`timescale 1ns / 1ps
`define INDEX (width+2)*(i/2+1)-1:(width+2)*i/2

module half_adder(
//inputs
	a,
	b,
//outputs
	o,
	cout
);

input wire a;
input wire b;
output wire o;
output wire cout;

`ifdef GSCL45NM
HAX1 HALFADD(.A(a),.B(b),.YS(o),.YC(cout));
`else
assign o = a^b;
assign cout = a&b;
`endif

endmodule

module compressor_3_2(
//inputs
	a,
	b,
	cin,
//outputs
	o,
	cout
);
input wire a;
input wire b;
input wire cin;
output wire o;
output wire cout;

`ifdef GSCL45NM
FAX1 FULLADD(.A(a),.B(b),.C(cin),.YS(o),.YC(cout));
`else
wire s = a^b;
wire g = a&b;

assign o = s^cin;
assign cout = s ? cin : g;
`endif

endmodule

module compressor_4_2(
//inputs
	a,
	b,
	c,
	d,
	cin,
//outputs
	o,
	co,
	cout
);

input wire a;
input wire b;
input wire c;
input wire d;
input wire cin;
output wire o;
output wire co;
output wire cout;
`ifdef FPGA_VERSION
wire carry;

compressor_3_2 FULLADD1(a,b,c,carry,cout);
compressor_3_2 FULLADD2(carry,d,cin,o,co);
`elsif GSCL45NM
wire carry;

FAX1 FULLADD1(.A(a),.B(b),.C(c),.YS(carry),.YC(cout));
FAX1 FULLADD2(.A(carry),.B(d),.C(cin),.YS(o),.YC(co));
`else
wire tmp1, tmp2, tmp3, tmp4, tmp5, tmp6;

assign tmp1 = ~(a&b);
assign tmp2 = ~(c&d);
assign tmp3 = ~((a|b)&tmp1);
assign tmp4 = ~((c|d)&tmp2);
assign tmp5 = ~((tmp1|tmp2)&(tmp3|tmp4));
assign tmp6 = tmp3^tmp4;
assign cout = ~(tmp1&tmp2);
assign co = tmp5|(tmp6&cin);
assign o = tmp6^cin;
`endif

endmodule

/********************************************************************************/

module _32_wallace_tree(
//inputs
	partial_products,
	carry,
//outputs
	compress_a,
	compress_b
);

localparam width = 32;

input wire [(width+2)*(width/2+1)-1:0] partial_products;
input wire [width/2-1:0] carry;
output wire [2*width-1:0] compress_a;
output wire [2*width-1:0] compress_b;

/* Input nets */
wire    s_0_0,    s_0_1,    s_1_0,    s_2_0,    s_2_1,    s_2_2;
wire    s_3_0,    s_3_1,    s_4_0,    s_4_1,    s_4_2,    s_4_3;
wire    s_5_0,    s_5_1,    s_5_2,    s_6_0,    s_6_1,    s_6_2;
wire    s_6_3,    s_6_4,    s_7_0,    s_7_1,    s_7_2,    s_7_3;
wire    s_8_0,    s_8_1,    s_8_2,    s_8_3,    s_8_4,    s_8_5;
wire    s_9_0,    s_9_1,    s_9_2,    s_9_3,    s_9_4,   s_10_0;
wire   s_10_1,   s_10_2,   s_10_3,   s_10_4,   s_10_5,   s_10_6;
wire   s_11_0,   s_11_1,   s_11_2,   s_11_3,   s_11_4,   s_11_5;
wire   s_12_0,   s_12_1,   s_12_2,   s_12_3,   s_12_4,   s_12_5;
wire   s_12_6,   s_12_7,   s_13_0,   s_13_1,   s_13_2,   s_13_3;
wire   s_13_4,   s_13_5,   s_13_6,   s_14_0,   s_14_1,   s_14_2;
wire   s_14_3,   s_14_4,   s_14_5,   s_14_6,   s_14_7,   s_14_8;
wire   s_15_0,   s_15_1,   s_15_2,   s_15_3,   s_15_4,   s_15_5;
wire   s_15_6,   s_15_7,   s_16_0,   s_16_1,   s_16_2,   s_16_3;
wire   s_16_4,   s_16_5,   s_16_6,   s_16_7,   s_16_8,   s_16_9;
wire   s_17_0,   s_17_1,   s_17_2,   s_17_3,   s_17_4,   s_17_5;
wire   s_17_6,   s_17_7,   s_17_8,   s_18_0,   s_18_1,   s_18_2;
wire   s_18_3,   s_18_4,   s_18_5,   s_18_6,   s_18_7,   s_18_8;
wire   s_18_9,  s_18_10,   s_19_0,   s_19_1,   s_19_2,   s_19_3;
wire   s_19_4,   s_19_5,   s_19_6,   s_19_7,   s_19_8,   s_19_9;
wire   s_20_0,   s_20_1,   s_20_2,   s_20_3,   s_20_4,   s_20_5;
wire   s_20_6,   s_20_7,   s_20_8,   s_20_9,  s_20_10,  s_20_11;
wire   s_21_0,   s_21_1,   s_21_2,   s_21_3,   s_21_4,   s_21_5;
wire   s_21_6,   s_21_7,   s_21_8,   s_21_9,  s_21_10,   s_22_0;
wire   s_22_1,   s_22_2,   s_22_3,   s_22_4,   s_22_5,   s_22_6;
wire   s_22_7,   s_22_8,   s_22_9,  s_22_10,  s_22_11,  s_22_12;
wire   s_23_0,   s_23_1,   s_23_2,   s_23_3,   s_23_4,   s_23_5;
wire   s_23_6,   s_23_7,   s_23_8,   s_23_9,  s_23_10,  s_23_11;
wire   s_24_0,   s_24_1,   s_24_2,   s_24_3,   s_24_4,   s_24_5;
wire   s_24_6,   s_24_7,   s_24_8,   s_24_9,  s_24_10,  s_24_11;
wire  s_24_12,  s_24_13,   s_25_0,   s_25_1,   s_25_2,   s_25_3;
wire   s_25_4,   s_25_5,   s_25_6,   s_25_7,   s_25_8,   s_25_9;
wire  s_25_10,  s_25_11,  s_25_12,   s_26_0,   s_26_1,   s_26_2;
wire   s_26_3,   s_26_4,   s_26_5,   s_26_6,   s_26_7,   s_26_8;
wire   s_26_9,  s_26_10,  s_26_11,  s_26_12,  s_26_13,  s_26_14;
wire   s_27_0,   s_27_1,   s_27_2,   s_27_3,   s_27_4,   s_27_5;
wire   s_27_6,   s_27_7,   s_27_8,   s_27_9,  s_27_10,  s_27_11;
wire  s_27_12,  s_27_13,   s_28_0,   s_28_1,   s_28_2,   s_28_3;
wire   s_28_4,   s_28_5,   s_28_6,   s_28_7,   s_28_8,   s_28_9;
wire  s_28_10,  s_28_11,  s_28_12,  s_28_13,  s_28_14,  s_28_15;
wire   s_29_0,   s_29_1,   s_29_2,   s_29_3,   s_29_4,   s_29_5;
wire   s_29_6,   s_29_7,   s_29_8,   s_29_9,  s_29_10,  s_29_11;
wire  s_29_12,  s_29_13,  s_29_14,   s_30_0,   s_30_1,   s_30_2;
wire   s_30_3,   s_30_4,   s_30_5,   s_30_6,   s_30_7,   s_30_8;
wire   s_30_9,  s_30_10,  s_30_11,  s_30_12,  s_30_13,  s_30_14;
wire  s_30_15,  s_30_16,   s_31_0,   s_31_1,   s_31_2,   s_31_3;
wire   s_31_4,   s_31_5,   s_31_6,   s_31_7,   s_31_8,   s_31_9;
wire  s_31_10,  s_31_11,  s_31_12,  s_31_13,  s_31_14,  s_31_15;
wire   s_32_0,   s_32_1,   s_32_2,   s_32_3,   s_32_4,   s_32_5;
wire   s_32_6,   s_32_7,   s_32_8,   s_32_9,  s_32_10,  s_32_11;
wire  s_32_12,  s_32_13,  s_32_14,  s_32_15,  s_32_16,   s_33_0;
wire   s_33_1,   s_33_2,   s_33_3,   s_33_4,   s_33_5,   s_33_6;
wire   s_33_7,   s_33_8,   s_33_9,  s_33_10,  s_33_11,  s_33_12;
wire  s_33_13,  s_33_14,  s_33_15,  s_33_16,   s_34_0,   s_34_1;
wire   s_34_2,   s_34_3,   s_34_4,   s_34_5,   s_34_6,   s_34_7;
wire   s_34_8,   s_34_9,  s_34_10,  s_34_11,  s_34_12,  s_34_13;
wire  s_34_14,  s_34_15,   s_35_0,   s_35_1,   s_35_2,   s_35_3;
wire   s_35_4,   s_35_5,   s_35_6,   s_35_7,   s_35_8,   s_35_9;
wire  s_35_10,  s_35_11,  s_35_12,  s_35_13,  s_35_14,  s_35_15;
wire   s_36_0,   s_36_1,   s_36_2,   s_36_3,   s_36_4,   s_36_5;
wire   s_36_6,   s_36_7,   s_36_8,   s_36_9,  s_36_10,  s_36_11;
wire  s_36_12,  s_36_13,  s_36_14,   s_37_0,   s_37_1,   s_37_2;
wire   s_37_3,   s_37_4,   s_37_5,   s_37_6,   s_37_7,   s_37_8;
wire   s_37_9,  s_37_10,  s_37_11,  s_37_12,  s_37_13,  s_37_14;
wire   s_38_0,   s_38_1,   s_38_2,   s_38_3,   s_38_4,   s_38_5;
wire   s_38_6,   s_38_7,   s_38_8,   s_38_9,  s_38_10,  s_38_11;
wire  s_38_12,  s_38_13,   s_39_0,   s_39_1,   s_39_2,   s_39_3;
wire   s_39_4,   s_39_5,   s_39_6,   s_39_7,   s_39_8,   s_39_9;
wire  s_39_10,  s_39_11,  s_39_12,  s_39_13,   s_40_0,   s_40_1;
wire   s_40_2,   s_40_3,   s_40_4,   s_40_5,   s_40_6,   s_40_7;
wire   s_40_8,   s_40_9,  s_40_10,  s_40_11,  s_40_12,   s_41_0;
wire   s_41_1,   s_41_2,   s_41_3,   s_41_4,   s_41_5,   s_41_6;
wire   s_41_7,   s_41_8,   s_41_9,  s_41_10,  s_41_11,  s_41_12;
wire   s_42_0,   s_42_1,   s_42_2,   s_42_3,   s_42_4,   s_42_5;
wire   s_42_6,   s_42_7,   s_42_8,   s_42_9,  s_42_10,  s_42_11;
wire   s_43_0,   s_43_1,   s_43_2,   s_43_3,   s_43_4,   s_43_5;
wire   s_43_6,   s_43_7,   s_43_8,   s_43_9,  s_43_10,  s_43_11;
wire   s_44_0,   s_44_1,   s_44_2,   s_44_3,   s_44_4,   s_44_5;
wire   s_44_6,   s_44_7,   s_44_8,   s_44_9,  s_44_10,   s_45_0;
wire   s_45_1,   s_45_2,   s_45_3,   s_45_4,   s_45_5,   s_45_6;
wire   s_45_7,   s_45_8,   s_45_9,  s_45_10,   s_46_0,   s_46_1;
wire   s_46_2,   s_46_3,   s_46_4,   s_46_5,   s_46_6,   s_46_7;
wire   s_46_8,   s_46_9,   s_47_0,   s_47_1,   s_47_2,   s_47_3;
wire   s_47_4,   s_47_5,   s_47_6,   s_47_7,   s_47_8,   s_47_9;
wire   s_48_0,   s_48_1,   s_48_2,   s_48_3,   s_48_4,   s_48_5;
wire   s_48_6,   s_48_7,   s_48_8,   s_49_0,   s_49_1,   s_49_2;
wire   s_49_3,   s_49_4,   s_49_5,   s_49_6,   s_49_7,   s_49_8;
wire   s_50_0,   s_50_1,   s_50_2,   s_50_3,   s_50_4,   s_50_5;
wire   s_50_6,   s_50_7,   s_51_0,   s_51_1,   s_51_2,   s_51_3;
wire   s_51_4,   s_51_5,   s_51_6,   s_51_7,   s_52_0,   s_52_1;
wire   s_52_2,   s_52_3,   s_52_4,   s_52_5,   s_52_6,   s_53_0;
wire   s_53_1,   s_53_2,   s_53_3,   s_53_4,   s_53_5,   s_53_6;
wire   s_54_0,   s_54_1,   s_54_2,   s_54_3,   s_54_4,   s_54_5;
wire   s_55_0,   s_55_1,   s_55_2,   s_55_3,   s_55_4,   s_55_5;
wire   s_56_0,   s_56_1,   s_56_2,   s_56_3,   s_56_4,   s_57_0;
wire   s_57_1,   s_57_2,   s_57_3,   s_57_4,   s_58_0,   s_58_1;
wire   s_58_2,   s_58_3,   s_59_0,   s_59_1,   s_59_2,   s_59_3;
wire   s_60_0,   s_60_1,   s_60_2,   s_61_0,   s_61_1,   s_61_2;
wire   s_62_0,   s_62_1,   s_63_0,   s_63_1;

assign {
 s_30_16,  s_28_15,  s_26_14,  s_24_13,  s_22_12,  s_20_11, 
 s_18_10,   s_16_9,   s_14_8,   s_12_7,   s_10_6,    s_8_5, 
   s_6_4,    s_4_3,    s_2_2,    s_0_1  
} = carry;

assign {
  s_33_0,   s_32_0,   s_31_0,   s_30_0,   s_29_0,   s_28_0, 
  s_27_0,   s_26_0,   s_25_0,   s_24_0,   s_23_0,   s_22_0, 
  s_21_0,   s_20_0,   s_19_0,   s_18_0,   s_17_0,   s_16_0, 
  s_15_0,   s_14_0,   s_13_0,   s_12_0,   s_11_0,   s_10_0, 
   s_9_0,    s_8_0,    s_7_0,    s_6_0,    s_5_0,    s_4_0, 
   s_3_0,    s_2_0,    s_1_0,    s_0_0  
} = partial_products[(width+2)*(0+1)-1:(width+2)*0];

assign {
  s_35_0,   s_34_0,   s_33_1,   s_32_1,   s_31_1,   s_30_1, 
  s_29_1,   s_28_1,   s_27_1,   s_26_1,   s_25_1,   s_24_1, 
  s_23_1,   s_22_1,   s_21_1,   s_20_1,   s_19_1,   s_18_1, 
  s_17_1,   s_16_1,   s_15_1,   s_14_1,   s_13_1,   s_12_1, 
  s_11_1,   s_10_1,    s_9_1,    s_8_1,    s_7_1,    s_6_1, 
   s_5_1,    s_4_1,    s_3_1,    s_2_1  
} = partial_products[(width+2)*(1+1)-1:(width+2)*1];

assign {
  s_37_0,   s_36_0,   s_35_1,   s_34_1,   s_33_2,   s_32_2, 
  s_31_2,   s_30_2,   s_29_2,   s_28_2,   s_27_2,   s_26_2, 
  s_25_2,   s_24_2,   s_23_2,   s_22_2,   s_21_2,   s_20_2, 
  s_19_2,   s_18_2,   s_17_2,   s_16_2,   s_15_2,   s_14_2, 
  s_13_2,   s_12_2,   s_11_2,   s_10_2,    s_9_2,    s_8_2, 
   s_7_2,    s_6_2,    s_5_2,    s_4_2  
} = partial_products[(width+2)*(2+1)-1:(width+2)*2];

assign {
  s_39_0,   s_38_0,   s_37_1,   s_36_1,   s_35_2,   s_34_2, 
  s_33_3,   s_32_3,   s_31_3,   s_30_3,   s_29_3,   s_28_3, 
  s_27_3,   s_26_3,   s_25_3,   s_24_3,   s_23_3,   s_22_3, 
  s_21_3,   s_20_3,   s_19_3,   s_18_3,   s_17_3,   s_16_3, 
  s_15_3,   s_14_3,   s_13_3,   s_12_3,   s_11_3,   s_10_3, 
   s_9_3,    s_8_3,    s_7_3,    s_6_3  
} = partial_products[(width+2)*(3+1)-1:(width+2)*3];

assign {
  s_41_0,   s_40_0,   s_39_1,   s_38_1,   s_37_2,   s_36_2, 
  s_35_3,   s_34_3,   s_33_4,   s_32_4,   s_31_4,   s_30_4, 
  s_29_4,   s_28_4,   s_27_4,   s_26_4,   s_25_4,   s_24_4, 
  s_23_4,   s_22_4,   s_21_4,   s_20_4,   s_19_4,   s_18_4, 
  s_17_4,   s_16_4,   s_15_4,   s_14_4,   s_13_4,   s_12_4, 
  s_11_4,   s_10_4,    s_9_4,    s_8_4  
} = partial_products[(width+2)*(4+1)-1:(width+2)*4];

assign {
  s_43_0,   s_42_0,   s_41_1,   s_40_1,   s_39_2,   s_38_2, 
  s_37_3,   s_36_3,   s_35_4,   s_34_4,   s_33_5,   s_32_5, 
  s_31_5,   s_30_5,   s_29_5,   s_28_5,   s_27_5,   s_26_5, 
  s_25_5,   s_24_5,   s_23_5,   s_22_5,   s_21_5,   s_20_5, 
  s_19_5,   s_18_5,   s_17_5,   s_16_5,   s_15_5,   s_14_5, 
  s_13_5,   s_12_5,   s_11_5,   s_10_5  
} = partial_products[(width+2)*(5+1)-1:(width+2)*5];

assign {
  s_45_0,   s_44_0,   s_43_1,   s_42_1,   s_41_2,   s_40_2, 
  s_39_3,   s_38_3,   s_37_4,   s_36_4,   s_35_5,   s_34_5, 
  s_33_6,   s_32_6,   s_31_6,   s_30_6,   s_29_6,   s_28_6, 
  s_27_6,   s_26_6,   s_25_6,   s_24_6,   s_23_6,   s_22_6, 
  s_21_6,   s_20_6,   s_19_6,   s_18_6,   s_17_6,   s_16_6, 
  s_15_6,   s_14_6,   s_13_6,   s_12_6  
} = partial_products[(width+2)*(6+1)-1:(width+2)*6];

assign {
  s_47_0,   s_46_0,   s_45_1,   s_44_1,   s_43_2,   s_42_2, 
  s_41_3,   s_40_3,   s_39_4,   s_38_4,   s_37_5,   s_36_5, 
  s_35_6,   s_34_6,   s_33_7,   s_32_7,   s_31_7,   s_30_7, 
  s_29_7,   s_28_7,   s_27_7,   s_26_7,   s_25_7,   s_24_7, 
  s_23_7,   s_22_7,   s_21_7,   s_20_7,   s_19_7,   s_18_7, 
  s_17_7,   s_16_7,   s_15_7,   s_14_7  
} = partial_products[(width+2)*(7+1)-1:(width+2)*7];

assign {
  s_49_0,   s_48_0,   s_47_1,   s_46_1,   s_45_2,   s_44_2, 
  s_43_3,   s_42_3,   s_41_4,   s_40_4,   s_39_5,   s_38_5, 
  s_37_6,   s_36_6,   s_35_7,   s_34_7,   s_33_8,   s_32_8, 
  s_31_8,   s_30_8,   s_29_8,   s_28_8,   s_27_8,   s_26_8, 
  s_25_8,   s_24_8,   s_23_8,   s_22_8,   s_21_8,   s_20_8, 
  s_19_8,   s_18_8,   s_17_8,   s_16_8  
} = partial_products[(width+2)*(8+1)-1:(width+2)*8];

assign {
  s_51_0,   s_50_0,   s_49_1,   s_48_1,   s_47_2,   s_46_2, 
  s_45_3,   s_44_3,   s_43_4,   s_42_4,   s_41_5,   s_40_5, 
  s_39_6,   s_38_6,   s_37_7,   s_36_7,   s_35_8,   s_34_8, 
  s_33_9,   s_32_9,   s_31_9,   s_30_9,   s_29_9,   s_28_9, 
  s_27_9,   s_26_9,   s_25_9,   s_24_9,   s_23_9,   s_22_9, 
  s_21_9,   s_20_9,   s_19_9,   s_18_9  
} = partial_products[(width+2)*(9+1)-1:(width+2)*9];

assign {
  s_53_0,   s_52_0,   s_51_1,   s_50_1,   s_49_2,   s_48_2, 
  s_47_3,   s_46_3,   s_45_4,   s_44_4,   s_43_5,   s_42_5, 
  s_41_6,   s_40_6,   s_39_7,   s_38_7,   s_37_8,   s_36_8, 
  s_35_9,   s_34_9,  s_33_10,  s_32_10,  s_31_10,  s_30_10, 
 s_29_10,  s_28_10,  s_27_10,  s_26_10,  s_25_10,  s_24_10, 
 s_23_10,  s_22_10,  s_21_10,  s_20_10  
} = partial_products[(width+2)*(10+1)-1:(width+2)*10];

assign {
  s_55_0,   s_54_0,   s_53_1,   s_52_1,   s_51_2,   s_50_2, 
  s_49_3,   s_48_3,   s_47_4,   s_46_4,   s_45_5,   s_44_5, 
  s_43_6,   s_42_6,   s_41_7,   s_40_7,   s_39_8,   s_38_8, 
  s_37_9,   s_36_9,  s_35_10,  s_34_10,  s_33_11,  s_32_11, 
 s_31_11,  s_30_11,  s_29_11,  s_28_11,  s_27_11,  s_26_11, 
 s_25_11,  s_24_11,  s_23_11,  s_22_11  
} = partial_products[(width+2)*(11+1)-1:(width+2)*11];

assign {
  s_57_0,   s_56_0,   s_55_1,   s_54_1,   s_53_2,   s_52_2, 
  s_51_3,   s_50_3,   s_49_4,   s_48_4,   s_47_5,   s_46_5, 
  s_45_6,   s_44_6,   s_43_7,   s_42_7,   s_41_8,   s_40_8, 
  s_39_9,   s_38_9,  s_37_10,  s_36_10,  s_35_11,  s_34_11, 
 s_33_12,  s_32_12,  s_31_12,  s_30_12,  s_29_12,  s_28_12, 
 s_27_12,  s_26_12,  s_25_12,  s_24_12  
} = partial_products[(width+2)*(12+1)-1:(width+2)*12];

assign {
  s_59_0,   s_58_0,   s_57_1,   s_56_1,   s_55_2,   s_54_2, 
  s_53_3,   s_52_3,   s_51_4,   s_50_4,   s_49_5,   s_48_5, 
  s_47_6,   s_46_6,   s_45_7,   s_44_7,   s_43_8,   s_42_8, 
  s_41_9,   s_40_9,  s_39_10,  s_38_10,  s_37_11,  s_36_11, 
 s_35_12,  s_34_12,  s_33_13,  s_32_13,  s_31_13,  s_30_13, 
 s_29_13,  s_28_13,  s_27_13,  s_26_13  
} = partial_products[(width+2)*(13+1)-1:(width+2)*13];

assign {
  s_61_0,   s_60_0,   s_59_1,   s_58_1,   s_57_2,   s_56_2, 
  s_55_3,   s_54_3,   s_53_4,   s_52_4,   s_51_5,   s_50_5, 
  s_49_6,   s_48_6,   s_47_7,   s_46_7,   s_45_8,   s_44_8, 
  s_43_9,   s_42_9,  s_41_10,  s_40_10,  s_39_11,  s_38_11, 
 s_37_12,  s_36_12,  s_35_13,  s_34_13,  s_33_14,  s_32_14, 
 s_31_14,  s_30_14,  s_29_14,  s_28_14  
} = partial_products[(width+2)*(14+1)-1:(width+2)*14];

assign {
  s_63_0,   s_62_0,   s_61_1,   s_60_1,   s_59_2,   s_58_2, 
  s_57_3,   s_56_3,   s_55_4,   s_54_4,   s_53_5,   s_52_5, 
  s_51_6,   s_50_6,   s_49_7,   s_48_7,   s_47_8,   s_46_8, 
  s_45_9,   s_44_9,  s_43_10,  s_42_10,  s_41_11,  s_40_11, 
 s_39_12,  s_38_12,  s_37_13,  s_36_13,  s_35_14,  s_34_14, 
 s_33_15,  s_32_15,  s_31_15,  s_30_15  
} = partial_products[(width+2)*(15+1)-1:(width+2)*15];

assign {
  s_63_1,   s_62_1,   s_61_2,   s_60_2,   s_59_3,   s_58_3, 
  s_57_4,   s_56_4,   s_55_5,   s_54_5,   s_53_6,   s_52_6, 
  s_51_7,   s_50_7,   s_49_8,   s_48_8,   s_47_9,   s_46_9, 
 s_45_10,  s_44_10,  s_43_11,  s_42_11,  s_41_12,  s_40_12, 
 s_39_13,  s_38_13,  s_37_14,  s_36_14,  s_35_15,  s_34_15, 
 s_33_16,  s_32_16  
} = partial_products[(width+2)*(width/2+1)-1:(width+2)*width/2+2];

/* u0_1 Output nets */
wire t_0,      t_1;
/* u1_2 Output nets */
wire t_2,      t_3;
/* u0_3 Output nets */
wire t_4,      t_5;
/* u2_4 Output nets */
wire t_6,      t_7,      t_8;
/* u1_5 Output nets */
wire t_9,     t_10;
/* u2_6 Output nets */
wire t_11,     t_12,     t_13;
/* u2_7 Output nets */
wire t_14,     t_15,     t_16;
/* u2_8 Output nets */
wire t_17,     t_18,     t_19;
/* u0_9 Output nets */
wire t_20,     t_21;
/* u2_10 Output nets */
wire t_22,     t_23,     t_24;
/* u0_11 Output nets */
wire t_25,     t_26;
/* u2_12 Output nets */
wire t_27,     t_28,     t_29;
/* u1_13 Output nets */
wire t_30,     t_31;
/* u2_14 Output nets */
wire t_32,     t_33,     t_34;
/* u1_15 Output nets */
wire t_35,     t_36;
/* u2_16 Output nets */
wire t_37,     t_38,     t_39;
/* u2_17 Output nets */
wire t_40,     t_41,     t_42;
/* u2_18 Output nets */
wire t_43,     t_44,     t_45;
/* u1_19 Output nets */
wire t_46,     t_47;
/* u2_20 Output nets */
wire t_48,     t_49,     t_50;
/* u2_21 Output nets */
wire t_51,     t_52,     t_53;
/* u2_22 Output nets */
wire t_54,     t_55,     t_56;
/* u2_23 Output nets */
wire t_57,     t_58,     t_59;
/* u2_24 Output nets */
wire t_60,     t_61,     t_62;
/* u2_25 Output nets */
wire t_63,     t_64,     t_65;
/* u0_26 Output nets */
wire t_66,     t_67;
/* u2_27 Output nets */
wire t_68,     t_69,     t_70;
/* u2_28 Output nets */
wire t_71,     t_72,     t_73;
/* u0_29 Output nets */
wire t_74,     t_75;
/* u2_30 Output nets */
wire t_76,     t_77,     t_78;
/* u2_31 Output nets */
wire t_79,     t_80,     t_81;
/* u1_32 Output nets */
wire t_82,     t_83;
/* u2_33 Output nets */
wire t_84,     t_85,     t_86;
/* u2_34 Output nets */
wire t_87,     t_88,     t_89;
/* u1_35 Output nets */
wire t_90,     t_91;
/* u2_36 Output nets */
wire t_92,     t_93,     t_94;
/* u2_37 Output nets */
wire t_95,     t_96,     t_97;
/* u2_38 Output nets */
wire t_98,     t_99,    t_100;
/* u2_39 Output nets */
wire t_101,    t_102,    t_103;
/* u2_40 Output nets */
wire t_104,    t_105,    t_106;
/* u1_41 Output nets */
wire t_107,    t_108;
/* u2_42 Output nets */
wire t_109,    t_110,    t_111;
/* u2_43 Output nets */
wire t_112,    t_113,    t_114;
/* u2_44 Output nets */
wire t_115,    t_116,    t_117;
/* u2_45 Output nets */
wire t_118,    t_119,    t_120;
/* u2_46 Output nets */
wire t_121,    t_122,    t_123;
/* u2_47 Output nets */
wire t_124,    t_125,    t_126;
/* u2_48 Output nets */
wire t_127,    t_128,    t_129;
/* u2_49 Output nets */
wire t_130,    t_131,    t_132;
/* u2_50 Output nets */
wire t_133,    t_134,    t_135;
/* u0_51 Output nets */
wire t_136,    t_137;
/* u2_52 Output nets */
wire t_138,    t_139,    t_140;
/* u2_53 Output nets */
wire t_141,    t_142,    t_143;
/* u2_54 Output nets */
wire t_144,    t_145,    t_146;
/* u0_55 Output nets */
wire t_147,    t_148;
/* u2_56 Output nets */
wire t_149,    t_150,    t_151;
/* u2_57 Output nets */
wire t_152,    t_153,    t_154;
/* u2_58 Output nets */
wire t_155,    t_156,    t_157;
/* u1_59 Output nets */
wire t_158,    t_159;
/* u2_60 Output nets */
wire t_160,    t_161,    t_162;
/* u2_61 Output nets */
wire t_163,    t_164,    t_165;
/* u2_62 Output nets */
wire t_166,    t_167,    t_168;
/* u1_63 Output nets */
wire t_169,    t_170;
/* u2_64 Output nets */
wire t_171,    t_172,    t_173;
/* u2_65 Output nets */
wire t_174,    t_175,    t_176;
/* u2_66 Output nets */
wire t_177,    t_178,    t_179;
/* u2_67 Output nets */
wire t_180,    t_181,    t_182;
/* u2_68 Output nets */
wire t_183,    t_184,    t_185;
/* u2_69 Output nets */
wire t_186,    t_187,    t_188;
/* u2_70 Output nets */
wire t_189,    t_190,    t_191;
/* u1_71 Output nets */
wire t_192,    t_193;
/* u2_72 Output nets */
wire t_194,    t_195,    t_196;
/* u2_73 Output nets */
wire t_197,    t_198,    t_199;
/* u2_74 Output nets */
wire t_200,    t_201,    t_202;
/* u2_75 Output nets */
wire t_203,    t_204,    t_205;
/* u2_76 Output nets */
wire t_206,    t_207,    t_208;
/* u2_77 Output nets */
wire t_209,    t_210,    t_211;
/* u2_78 Output nets */
wire t_212,    t_213,    t_214;
/* u2_79 Output nets */
wire t_215,    t_216,    t_217;
/* u2_80 Output nets */
wire t_218,    t_219,    t_220;
/* u2_81 Output nets */
wire t_221,    t_222,    t_223;
/* u2_82 Output nets */
wire t_224,    t_225,    t_226;
/* u2_83 Output nets */
wire t_227,    t_228,    t_229;
/* u2_84 Output nets */
wire t_230,    t_231,    t_232;
/* u2_85 Output nets */
wire t_233,    t_234,    t_235;
/* u2_86 Output nets */
wire t_236,    t_237,    t_238;
/* u2_87 Output nets */
wire t_239,    t_240,    t_241;
/* u2_88 Output nets */
wire t_242,    t_243,    t_244;
/* u2_89 Output nets */
wire t_245,    t_246,    t_247;
/* u2_90 Output nets */
wire t_248,    t_249,    t_250;
/* u2_91 Output nets */
wire t_251,    t_252,    t_253;
/* u2_92 Output nets */
wire t_254,    t_255,    t_256;
/* u2_93 Output nets */
wire t_257,    t_258,    t_259;
/* u2_94 Output nets */
wire t_260,    t_261,    t_262;
/* u2_95 Output nets */
wire t_263,    t_264,    t_265;
/* u2_96 Output nets */
wire t_266,    t_267,    t_268;
/* u2_97 Output nets */
wire t_269,    t_270,    t_271;
/* u2_98 Output nets */
wire t_272,    t_273,    t_274;
/* u1_99 Output nets */
wire t_275,    t_276;
/* u2_100 Output nets */
wire t_277,    t_278,    t_279;
/* u2_101 Output nets */
wire t_280,    t_281,    t_282;
/* u2_102 Output nets */
wire t_283,    t_284,    t_285;
/* u1_103 Output nets */
wire t_286,    t_287;
/* u2_104 Output nets */
wire t_288,    t_289,    t_290;
/* u2_105 Output nets */
wire t_291,    t_292,    t_293;
/* u2_106 Output nets */
wire t_294,    t_295,    t_296;
/* u1_107 Output nets */
wire t_297,    t_298;
/* u2_108 Output nets */
wire t_299,    t_300,    t_301;
/* u2_109 Output nets */
wire t_302,    t_303,    t_304;
/* u2_110 Output nets */
wire t_305,    t_306,    t_307;
/* u1_111 Output nets */
wire t_308,    t_309;
/* u2_112 Output nets */
wire t_310,    t_311,    t_312;
/* u2_113 Output nets */
wire t_313,    t_314,    t_315;
/* u2_114 Output nets */
wire t_316,    t_317,    t_318;
/* u0_115 Output nets */
wire t_319,    t_320;
/* u2_116 Output nets */
wire t_321,    t_322,    t_323;
/* u2_117 Output nets */
wire t_324,    t_325,    t_326;
/* u2_118 Output nets */
wire t_327,    t_328,    t_329;
/* u0_119 Output nets */
wire t_330,    t_331;
/* u2_120 Output nets */
wire t_332,    t_333,    t_334;
/* u2_121 Output nets */
wire t_335,    t_336,    t_337;
/* u2_122 Output nets */
wire t_338,    t_339,    t_340;
/* u2_123 Output nets */
wire t_341,    t_342,    t_343;
/* u2_124 Output nets */
wire t_344,    t_345,    t_346;
/* u2_125 Output nets */
wire t_347,    t_348,    t_349;
/* u2_126 Output nets */
wire t_350,    t_351,    t_352;
/* u2_127 Output nets */
wire t_353,    t_354,    t_355;
/* u1_128 Output nets */
wire t_356,    t_357;
/* u2_129 Output nets */
wire t_358,    t_359,    t_360;
/* u2_130 Output nets */
wire t_361,    t_362,    t_363;
/* u1_131 Output nets */
wire t_364,    t_365;
/* u2_132 Output nets */
wire t_366,    t_367,    t_368;
/* u2_133 Output nets */
wire t_369,    t_370,    t_371;
/* u1_134 Output nets */
wire t_372,    t_373;
/* u2_135 Output nets */
wire t_374,    t_375,    t_376;
/* u2_136 Output nets */
wire t_377,    t_378,    t_379;
/* u1_137 Output nets */
wire t_380,    t_381;
/* u2_138 Output nets */
wire t_382,    t_383,    t_384;
/* u2_139 Output nets */
wire t_385,    t_386,    t_387;
/* u0_140 Output nets */
wire t_388,    t_389;
/* u2_141 Output nets */
wire t_390,    t_391,    t_392;
/* u2_142 Output nets */
wire t_393,    t_394,    t_395;
/* u0_143 Output nets */
wire t_396,    t_397;
/* u2_144 Output nets */
wire t_398,    t_399,    t_400;
/* u2_145 Output nets */
wire t_401,    t_402,    t_403;
/* u2_146 Output nets */
wire t_404,    t_405,    t_406;
/* u2_147 Output nets */
wire t_407,    t_408,    t_409;
/* u2_148 Output nets */
wire t_410,    t_411,    t_412;
/* u1_149 Output nets */
wire t_413,    t_414;
/* u2_150 Output nets */
wire t_415,    t_416,    t_417;
/* u1_151 Output nets */
wire t_418,    t_419;
/* u2_152 Output nets */
wire t_420,    t_421,    t_422;
/* u1_153 Output nets */
wire t_423,    t_424;
/* u2_154 Output nets */
wire t_425,    t_426,    t_427;
/* u1_155 Output nets */
wire t_428,    t_429;
/* u2_156 Output nets */
wire t_430,    t_431,    t_432;
/* u0_157 Output nets */
wire t_433,    t_434;
/* u2_158 Output nets */
wire t_435,    t_436,    t_437;
/* u0_159 Output nets */
wire t_438,    t_439;
/* u2_160 Output nets */
wire t_440,    t_441,    t_442;
/* u2_161 Output nets */
wire t_443,    t_444,    t_445;
/* u1_162 Output nets */
wire t_446,    t_447;
/* u1_163 Output nets */
wire t_448,    t_449;
/* u0_164 Output nets */
wire t_450,    t_451;
/* u0_165 Output nets */
wire t_452;

/* compress stage 1 */
half_adder u0_1(.a(s_0_1), .b(s_0_0), .o(t_0), .cout(t_1));
compressor_3_2 u1_2(.a(s_2_2), .b(s_2_1), .cin(s_2_0), .o(t_2), .cout(t_3));
half_adder u0_3(.a(s_3_1), .b(s_3_0), .o(t_4), .cout(t_5));
compressor_4_2 u2_4(.a(s_4_3), .b(s_4_2), .c(s_4_1), .d(s_4_0), .cin(t_5), .o(t_6), .co(t_7), .cout(t_8));
compressor_3_2 u1_5(.a(s_5_1), .b(s_5_0), .cin(t_8), .o(t_9), .cout(t_10));
compressor_4_2 u2_6(.a(s_6_4), .b(s_6_3), .c(s_6_2), .d(s_6_1), .cin(s_6_0), .o(t_11), .co(t_12), .cout(t_13));
compressor_4_2 u2_7(.a(s_7_3), .b(s_7_2), .c(s_7_1), .d(s_7_0), .cin(t_13), .o(t_14), .co(t_15), .cout(t_16));
compressor_4_2 u2_8(.a(s_8_3), .b(s_8_2), .c(s_8_1), .d(s_8_0), .cin(t_16), .o(t_17), .co(t_18), .cout(t_19));
half_adder u0_9(.a(s_8_5), .b(s_8_4), .o(t_20), .cout(t_21));
compressor_4_2 u2_10(.a(s_9_2), .b(s_9_1), .c(s_9_0), .d(t_19), .cin(t_21), .o(t_22), .co(t_23), .cout(t_24));
half_adder u0_11(.a(s_9_4), .b(s_9_3), .o(t_25), .cout(t_26));
compressor_4_2 u2_12(.a(s_10_2), .b(s_10_1), .c(s_10_0), .d(t_24), .cin(t_26), .o(t_27), .co(t_28), .cout(t_29));
compressor_3_2 u1_13(.a(s_10_5), .b(s_10_4), .cin(s_10_3), .o(t_30), .cout(t_31));
compressor_4_2 u2_14(.a(s_11_2), .b(s_11_1), .c(s_11_0), .d(t_29), .cin(t_31), .o(t_32), .co(t_33), .cout(t_34));
compressor_3_2 u1_15(.a(s_11_5), .b(s_11_4), .cin(s_11_3), .o(t_35), .cout(t_36));
compressor_4_2 u2_16(.a(s_12_2), .b(s_12_1), .c(s_12_0), .d(t_34), .cin(t_36), .o(t_37), .co(t_38), .cout(t_39));
compressor_4_2 u2_17(.a(s_12_7), .b(s_12_6), .c(s_12_5), .d(s_12_4), .cin(s_12_3), .o(t_40), .co(t_41), .cout(t_42));
compressor_4_2 u2_18(.a(s_13_2), .b(s_13_1), .c(s_13_0), .d(t_39), .cin(t_42), .o(t_43), .co(t_44), .cout(t_45));
compressor_3_2 u1_19(.a(s_13_5), .b(s_13_4), .cin(s_13_3), .o(t_46), .cout(t_47));
compressor_4_2 u2_20(.a(s_14_2), .b(s_14_1), .c(s_14_0), .d(t_45), .cin(t_47), .o(t_48), .co(t_49), .cout(t_50));
compressor_4_2 u2_21(.a(s_14_7), .b(s_14_6), .c(s_14_5), .d(s_14_4), .cin(s_14_3), .o(t_51), .co(t_52), .cout(t_53));
compressor_4_2 u2_22(.a(s_15_2), .b(s_15_1), .c(s_15_0), .d(t_50), .cin(t_53), .o(t_54), .co(t_55), .cout(t_56));
compressor_4_2 u2_23(.a(s_15_7), .b(s_15_6), .c(s_15_5), .d(s_15_4), .cin(s_15_3), .o(t_57), .co(t_58), .cout(t_59));
compressor_4_2 u2_24(.a(s_16_2), .b(s_16_1), .c(s_16_0), .d(t_56), .cin(t_59), .o(t_60), .co(t_61), .cout(t_62));
compressor_4_2 u2_25(.a(s_16_7), .b(s_16_6), .c(s_16_5), .d(s_16_4), .cin(s_16_3), .o(t_63), .co(t_64), .cout(t_65));
half_adder u0_26(.a(s_16_9), .b(s_16_8), .o(t_66), .cout(t_67));
compressor_4_2 u2_27(.a(s_17_2), .b(s_17_1), .c(s_17_0), .d(t_62), .cin(t_65), .o(t_68), .co(t_69), .cout(t_70));
compressor_4_2 u2_28(.a(s_17_6), .b(s_17_5), .c(s_17_4), .d(s_17_3), .cin(t_67), .o(t_71), .co(t_72), .cout(t_73));
half_adder u0_29(.a(s_17_8), .b(s_17_7), .o(t_74), .cout(t_75));
compressor_4_2 u2_30(.a(s_18_2), .b(s_18_1), .c(s_18_0), .d(t_70), .cin(t_73), .o(t_76), .co(t_77), .cout(t_78));
compressor_4_2 u2_31(.a(s_18_6), .b(s_18_5), .c(s_18_4), .d(s_18_3), .cin(t_75), .o(t_79), .co(t_80), .cout(t_81));
compressor_3_2 u1_32(.a(s_18_9), .b(s_18_8), .cin(s_18_7), .o(t_82), .cout(t_83));
compressor_4_2 u2_33(.a(s_19_2), .b(s_19_1), .c(s_19_0), .d(t_78), .cin(t_81), .o(t_84), .co(t_85), .cout(t_86));
compressor_4_2 u2_34(.a(s_19_6), .b(s_19_5), .c(s_19_4), .d(s_19_3), .cin(t_83), .o(t_87), .co(t_88), .cout(t_89));
compressor_3_2 u1_35(.a(s_19_9), .b(s_19_8), .cin(s_19_7), .o(t_90), .cout(t_91));
compressor_4_2 u2_36(.a(s_20_2), .b(s_20_1), .c(s_20_0), .d(t_86), .cin(t_89), .o(t_92), .co(t_93), .cout(t_94));
compressor_4_2 u2_37(.a(s_20_6), .b(s_20_5), .c(s_20_4), .d(s_20_3), .cin(t_91), .o(t_95), .co(t_96), .cout(t_97));
compressor_4_2 u2_38(.a(s_20_11), .b(s_20_10), .c(s_20_9), .d(s_20_8), .cin(s_20_7), .o(t_98), .co(t_99), .cout(t_100));
compressor_4_2 u2_39(.a(s_21_2), .b(s_21_1), .c(s_21_0), .d(t_94), .cin(t_97), .o(t_101), .co(t_102), .cout(t_103));
compressor_4_2 u2_40(.a(s_21_6), .b(s_21_5), .c(s_21_4), .d(s_21_3), .cin(t_100), .o(t_104), .co(t_105), .cout(t_106));
compressor_3_2 u1_41(.a(s_21_9), .b(s_21_8), .cin(s_21_7), .o(t_107), .cout(t_108));
compressor_4_2 u2_42(.a(s_22_2), .b(s_22_1), .c(s_22_0), .d(t_103), .cin(t_106), .o(t_109), .co(t_110), .cout(t_111));
compressor_4_2 u2_43(.a(s_22_6), .b(s_22_5), .c(s_22_4), .d(s_22_3), .cin(t_108), .o(t_112), .co(t_113), .cout(t_114));
compressor_4_2 u2_44(.a(s_22_11), .b(s_22_10), .c(s_22_9), .d(s_22_8), .cin(s_22_7), .o(t_115), .co(t_116), .cout(t_117));
compressor_4_2 u2_45(.a(s_23_2), .b(s_23_1), .c(s_23_0), .d(t_111), .cin(t_114), .o(t_118), .co(t_119), .cout(t_120));
compressor_4_2 u2_46(.a(s_23_6), .b(s_23_5), .c(s_23_4), .d(s_23_3), .cin(t_117), .o(t_121), .co(t_122), .cout(t_123));
compressor_4_2 u2_47(.a(s_23_11), .b(s_23_10), .c(s_23_9), .d(s_23_8), .cin(s_23_7), .o(t_124), .co(t_125), .cout(t_126));
compressor_4_2 u2_48(.a(s_24_2), .b(s_24_1), .c(s_24_0), .d(t_120), .cin(t_123), .o(t_127), .co(t_128), .cout(t_129));
compressor_4_2 u2_49(.a(s_24_6), .b(s_24_5), .c(s_24_4), .d(s_24_3), .cin(t_126), .o(t_130), .co(t_131), .cout(t_132));
compressor_4_2 u2_50(.a(s_24_11), .b(s_24_10), .c(s_24_9), .d(s_24_8), .cin(s_24_7), .o(t_133), .co(t_134), .cout(t_135));
half_adder u0_51(.a(s_24_13), .b(s_24_12), .o(t_136), .cout(t_137));
compressor_4_2 u2_52(.a(s_25_2), .b(s_25_1), .c(s_25_0), .d(t_129), .cin(t_132), .o(t_138), .co(t_139), .cout(t_140));
compressor_4_2 u2_53(.a(s_25_5), .b(s_25_4), .c(s_25_3), .d(t_135), .cin(t_137), .o(t_141), .co(t_142), .cout(t_143));
compressor_4_2 u2_54(.a(s_25_10), .b(s_25_9), .c(s_25_8), .d(s_25_7), .cin(s_25_6), .o(t_144), .co(t_145), .cout(t_146));
half_adder u0_55(.a(s_25_12), .b(s_25_11), .o(t_147), .cout(t_148));
compressor_4_2 u2_56(.a(s_26_2), .b(s_26_1), .c(s_26_0), .d(t_140), .cin(t_143), .o(t_149), .co(t_150), .cout(t_151));
compressor_4_2 u2_57(.a(s_26_5), .b(s_26_4), .c(s_26_3), .d(t_146), .cin(t_148), .o(t_152), .co(t_153), .cout(t_154));
compressor_4_2 u2_58(.a(s_26_10), .b(s_26_9), .c(s_26_8), .d(s_26_7), .cin(s_26_6), .o(t_155), .co(t_156), .cout(t_157));
compressor_3_2 u1_59(.a(s_26_13), .b(s_26_12), .cin(s_26_11), .o(t_158), .cout(t_159));
compressor_4_2 u2_60(.a(s_27_2), .b(s_27_1), .c(s_27_0), .d(t_151), .cin(t_154), .o(t_160), .co(t_161), .cout(t_162));
compressor_4_2 u2_61(.a(s_27_5), .b(s_27_4), .c(s_27_3), .d(t_157), .cin(t_159), .o(t_163), .co(t_164), .cout(t_165));
compressor_4_2 u2_62(.a(s_27_10), .b(s_27_9), .c(s_27_8), .d(s_27_7), .cin(s_27_6), .o(t_166), .co(t_167), .cout(t_168));
compressor_3_2 u1_63(.a(s_27_13), .b(s_27_12), .cin(s_27_11), .o(t_169), .cout(t_170));
compressor_4_2 u2_64(.a(s_28_2), .b(s_28_1), .c(s_28_0), .d(t_162), .cin(t_165), .o(t_171), .co(t_172), .cout(t_173));
compressor_4_2 u2_65(.a(s_28_5), .b(s_28_4), .c(s_28_3), .d(t_168), .cin(t_170), .o(t_174), .co(t_175), .cout(t_176));
compressor_4_2 u2_66(.a(s_28_10), .b(s_28_9), .c(s_28_8), .d(s_28_7), .cin(s_28_6), .o(t_177), .co(t_178), .cout(t_179));
compressor_4_2 u2_67(.a(s_28_15), .b(s_28_14), .c(s_28_13), .d(s_28_12), .cin(s_28_11), .o(t_180), .co(t_181), .cout(t_182));
compressor_4_2 u2_68(.a(s_29_2), .b(s_29_1), .c(s_29_0), .d(t_173), .cin(t_176), .o(t_183), .co(t_184), .cout(t_185));
compressor_4_2 u2_69(.a(s_29_5), .b(s_29_4), .c(s_29_3), .d(t_179), .cin(t_182), .o(t_186), .co(t_187), .cout(t_188));
compressor_4_2 u2_70(.a(s_29_10), .b(s_29_9), .c(s_29_8), .d(s_29_7), .cin(s_29_6), .o(t_189), .co(t_190), .cout(t_191));
compressor_3_2 u1_71(.a(s_29_13), .b(s_29_12), .cin(s_29_11), .o(t_192), .cout(t_193));
compressor_4_2 u2_72(.a(s_30_2), .b(s_30_1), .c(s_30_0), .d(t_185), .cin(t_188), .o(t_194), .co(t_195), .cout(t_196));
compressor_4_2 u2_73(.a(s_30_5), .b(s_30_4), .c(s_30_3), .d(t_191), .cin(t_193), .o(t_197), .co(t_198), .cout(t_199));
compressor_4_2 u2_74(.a(s_30_10), .b(s_30_9), .c(s_30_8), .d(s_30_7), .cin(s_30_6), .o(t_200), .co(t_201), .cout(t_202));
compressor_4_2 u2_75(.a(s_30_15), .b(s_30_14), .c(s_30_13), .d(s_30_12), .cin(s_30_11), .o(t_203), .co(t_204), .cout(t_205));
compressor_4_2 u2_76(.a(s_31_2), .b(s_31_1), .c(s_31_0), .d(t_196), .cin(t_199), .o(t_206), .co(t_207), .cout(t_208));
compressor_4_2 u2_77(.a(s_31_5), .b(s_31_4), .c(s_31_3), .d(t_202), .cin(t_205), .o(t_209), .co(t_210), .cout(t_211));
compressor_4_2 u2_78(.a(s_31_10), .b(s_31_9), .c(s_31_8), .d(s_31_7), .cin(s_31_6), .o(t_212), .co(t_213), .cout(t_214));
compressor_4_2 u2_79(.a(s_31_15), .b(s_31_14), .c(s_31_13), .d(s_31_12), .cin(s_31_11), .o(t_215), .co(t_216), .cout(t_217));
compressor_4_2 u2_80(.a(s_32_2), .b(s_32_1), .c(s_32_0), .d(t_208), .cin(t_211), .o(t_218), .co(t_219), .cout(t_220));
compressor_4_2 u2_81(.a(s_32_5), .b(s_32_4), .c(s_32_3), .d(t_214), .cin(t_217), .o(t_221), .co(t_222), .cout(t_223));
compressor_4_2 u2_82(.a(s_32_10), .b(s_32_9), .c(s_32_8), .d(s_32_7), .cin(s_32_6), .o(t_224), .co(t_225), .cout(t_226));
compressor_4_2 u2_83(.a(s_32_15), .b(s_32_14), .c(s_32_13), .d(s_32_12), .cin(s_32_11), .o(t_227), .co(t_228), .cout(t_229));
compressor_4_2 u2_84(.a(s_33_2), .b(s_33_1), .c(s_33_0), .d(t_220), .cin(t_223), .o(t_230), .co(t_231), .cout(t_232));
compressor_4_2 u2_85(.a(s_33_5), .b(s_33_4), .c(s_33_3), .d(t_226), .cin(t_229), .o(t_233), .co(t_234), .cout(t_235));
compressor_4_2 u2_86(.a(s_33_10), .b(s_33_9), .c(s_33_8), .d(s_33_7), .cin(s_33_6), .o(t_236), .co(t_237), .cout(t_238));
compressor_4_2 u2_87(.a(s_33_15), .b(s_33_14), .c(s_33_13), .d(s_33_12), .cin(s_33_11), .o(t_239), .co(t_240), .cout(t_241));
compressor_4_2 u2_88(.a(s_34_2), .b(s_34_1), .c(s_34_0), .d(t_232), .cin(t_235), .o(t_242), .co(t_243), .cout(t_244));
compressor_4_2 u2_89(.a(s_34_5), .b(s_34_4), .c(s_34_3), .d(t_238), .cin(t_241), .o(t_245), .co(t_246), .cout(t_247));
compressor_4_2 u2_90(.a(s_34_10), .b(s_34_9), .c(s_34_8), .d(s_34_7), .cin(s_34_6), .o(t_248), .co(t_249), .cout(t_250));
compressor_4_2 u2_91(.a(s_34_15), .b(s_34_14), .c(s_34_13), .d(s_34_12), .cin(s_34_11), .o(t_251), .co(t_252), .cout(t_253));
compressor_4_2 u2_92(.a(s_35_2), .b(s_35_1), .c(s_35_0), .d(t_244), .cin(t_247), .o(t_254), .co(t_255), .cout(t_256));
compressor_4_2 u2_93(.a(s_35_5), .b(s_35_4), .c(s_35_3), .d(t_250), .cin(t_253), .o(t_257), .co(t_258), .cout(t_259));
compressor_4_2 u2_94(.a(s_35_10), .b(s_35_9), .c(s_35_8), .d(s_35_7), .cin(s_35_6), .o(t_260), .co(t_261), .cout(t_262));
compressor_4_2 u2_95(.a(s_35_15), .b(s_35_14), .c(s_35_13), .d(s_35_12), .cin(s_35_11), .o(t_263), .co(t_264), .cout(t_265));
compressor_4_2 u2_96(.a(s_36_2), .b(s_36_1), .c(s_36_0), .d(t_256), .cin(t_259), .o(t_266), .co(t_267), .cout(t_268));
compressor_4_2 u2_97(.a(s_36_5), .b(s_36_4), .c(s_36_3), .d(t_262), .cin(t_265), .o(t_269), .co(t_270), .cout(t_271));
compressor_4_2 u2_98(.a(s_36_10), .b(s_36_9), .c(s_36_8), .d(s_36_7), .cin(s_36_6), .o(t_272), .co(t_273), .cout(t_274));
compressor_3_2 u1_99(.a(s_36_13), .b(s_36_12), .cin(s_36_11), .o(t_275), .cout(t_276));
compressor_4_2 u2_100(.a(s_37_2), .b(s_37_1), .c(s_37_0), .d(t_268), .cin(t_271), .o(t_277), .co(t_278), .cout(t_279));
compressor_4_2 u2_101(.a(s_37_5), .b(s_37_4), .c(s_37_3), .d(t_274), .cin(t_276), .o(t_280), .co(t_281), .cout(t_282));
compressor_4_2 u2_102(.a(s_37_10), .b(s_37_9), .c(s_37_8), .d(s_37_7), .cin(s_37_6), .o(t_283), .co(t_284), .cout(t_285));
compressor_3_2 u1_103(.a(s_37_13), .b(s_37_12), .cin(s_37_11), .o(t_286), .cout(t_287));
compressor_4_2 u2_104(.a(s_38_2), .b(s_38_1), .c(s_38_0), .d(t_279), .cin(t_282), .o(t_288), .co(t_289), .cout(t_290));
compressor_4_2 u2_105(.a(s_38_5), .b(s_38_4), .c(s_38_3), .d(t_285), .cin(t_287), .o(t_291), .co(t_292), .cout(t_293));
compressor_4_2 u2_106(.a(s_38_10), .b(s_38_9), .c(s_38_8), .d(s_38_7), .cin(s_38_6), .o(t_294), .co(t_295), .cout(t_296));
compressor_3_2 u1_107(.a(s_38_13), .b(s_38_12), .cin(s_38_11), .o(t_297), .cout(t_298));
compressor_4_2 u2_108(.a(s_39_2), .b(s_39_1), .c(s_39_0), .d(t_290), .cin(t_293), .o(t_299), .co(t_300), .cout(t_301));
compressor_4_2 u2_109(.a(s_39_5), .b(s_39_4), .c(s_39_3), .d(t_296), .cin(t_298), .o(t_302), .co(t_303), .cout(t_304));
compressor_4_2 u2_110(.a(s_39_10), .b(s_39_9), .c(s_39_8), .d(s_39_7), .cin(s_39_6), .o(t_305), .co(t_306), .cout(t_307));
compressor_3_2 u1_111(.a(s_39_13), .b(s_39_12), .cin(s_39_11), .o(t_308), .cout(t_309));
compressor_4_2 u2_112(.a(s_40_2), .b(s_40_1), .c(s_40_0), .d(t_301), .cin(t_304), .o(t_310), .co(t_311), .cout(t_312));
compressor_4_2 u2_113(.a(s_40_5), .b(s_40_4), .c(s_40_3), .d(t_307), .cin(t_309), .o(t_313), .co(t_314), .cout(t_315));
compressor_4_2 u2_114(.a(s_40_10), .b(s_40_9), .c(s_40_8), .d(s_40_7), .cin(s_40_6), .o(t_316), .co(t_317), .cout(t_318));
half_adder u0_115(.a(s_40_12), .b(s_40_11), .o(t_319), .cout(t_320));
compressor_4_2 u2_116(.a(s_41_2), .b(s_41_1), .c(s_41_0), .d(t_312), .cin(t_315), .o(t_321), .co(t_322), .cout(t_323));
compressor_4_2 u2_117(.a(s_41_5), .b(s_41_4), .c(s_41_3), .d(t_318), .cin(t_320), .o(t_324), .co(t_325), .cout(t_326));
compressor_4_2 u2_118(.a(s_41_10), .b(s_41_9), .c(s_41_8), .d(s_41_7), .cin(s_41_6), .o(t_327), .co(t_328), .cout(t_329));
half_adder u0_119(.a(s_41_12), .b(s_41_11), .o(t_330), .cout(t_331));
compressor_4_2 u2_120(.a(s_42_2), .b(s_42_1), .c(s_42_0), .d(t_323), .cin(t_326), .o(t_332), .co(t_333), .cout(t_334));
compressor_4_2 u2_121(.a(s_42_5), .b(s_42_4), .c(s_42_3), .d(t_329), .cin(t_331), .o(t_335), .co(t_336), .cout(t_337));
compressor_4_2 u2_122(.a(s_42_10), .b(s_42_9), .c(s_42_8), .d(s_42_7), .cin(s_42_6), .o(t_338), .co(t_339), .cout(t_340));
compressor_4_2 u2_123(.a(s_43_2), .b(s_43_1), .c(s_43_0), .d(t_334), .cin(t_337), .o(t_341), .co(t_342), .cout(t_343));
compressor_4_2 u2_124(.a(s_43_6), .b(s_43_5), .c(s_43_4), .d(s_43_3), .cin(t_340), .o(t_344), .co(t_345), .cout(t_346));
compressor_4_2 u2_125(.a(s_43_11), .b(s_43_10), .c(s_43_9), .d(s_43_8), .cin(s_43_7), .o(t_347), .co(t_348), .cout(t_349));
compressor_4_2 u2_126(.a(s_44_2), .b(s_44_1), .c(s_44_0), .d(t_343), .cin(t_346), .o(t_350), .co(t_351), .cout(t_352));
compressor_4_2 u2_127(.a(s_44_6), .b(s_44_5), .c(s_44_4), .d(s_44_3), .cin(t_349), .o(t_353), .co(t_354), .cout(t_355));
compressor_3_2 u1_128(.a(s_44_9), .b(s_44_8), .cin(s_44_7), .o(t_356), .cout(t_357));
compressor_4_2 u2_129(.a(s_45_2), .b(s_45_1), .c(s_45_0), .d(t_352), .cin(t_355), .o(t_358), .co(t_359), .cout(t_360));
compressor_4_2 u2_130(.a(s_45_6), .b(s_45_5), .c(s_45_4), .d(s_45_3), .cin(t_357), .o(t_361), .co(t_362), .cout(t_363));
compressor_3_2 u1_131(.a(s_45_9), .b(s_45_8), .cin(s_45_7), .o(t_364), .cout(t_365));
compressor_4_2 u2_132(.a(s_46_2), .b(s_46_1), .c(s_46_0), .d(t_360), .cin(t_363), .o(t_366), .co(t_367), .cout(t_368));
compressor_4_2 u2_133(.a(s_46_6), .b(s_46_5), .c(s_46_4), .d(s_46_3), .cin(t_365), .o(t_369), .co(t_370), .cout(t_371));
compressor_3_2 u1_134(.a(s_46_9), .b(s_46_8), .cin(s_46_7), .o(t_372), .cout(t_373));
compressor_4_2 u2_135(.a(s_47_2), .b(s_47_1), .c(s_47_0), .d(t_368), .cin(t_371), .o(t_374), .co(t_375), .cout(t_376));
compressor_4_2 u2_136(.a(s_47_6), .b(s_47_5), .c(s_47_4), .d(s_47_3), .cin(t_373), .o(t_377), .co(t_378), .cout(t_379));
compressor_3_2 u1_137(.a(s_47_9), .b(s_47_8), .cin(s_47_7), .o(t_380), .cout(t_381));
compressor_4_2 u2_138(.a(s_48_2), .b(s_48_1), .c(s_48_0), .d(t_376), .cin(t_379), .o(t_382), .co(t_383), .cout(t_384));
compressor_4_2 u2_139(.a(s_48_6), .b(s_48_5), .c(s_48_4), .d(s_48_3), .cin(t_381), .o(t_385), .co(t_386), .cout(t_387));
half_adder u0_140(.a(s_48_8), .b(s_48_7), .o(t_388), .cout(t_389));
compressor_4_2 u2_141(.a(s_49_2), .b(s_49_1), .c(s_49_0), .d(t_384), .cin(t_387), .o(t_390), .co(t_391), .cout(t_392));
compressor_4_2 u2_142(.a(s_49_6), .b(s_49_5), .c(s_49_4), .d(s_49_3), .cin(t_389), .o(t_393), .co(t_394), .cout(t_395));
half_adder u0_143(.a(s_49_8), .b(s_49_7), .o(t_396), .cout(t_397));
compressor_4_2 u2_144(.a(s_50_2), .b(s_50_1), .c(s_50_0), .d(t_392), .cin(t_395), .o(t_398), .co(t_399), .cout(t_400));
compressor_4_2 u2_145(.a(s_50_6), .b(s_50_5), .c(s_50_4), .d(s_50_3), .cin(t_397), .o(t_401), .co(t_402), .cout(t_403));
compressor_4_2 u2_146(.a(s_51_2), .b(s_51_1), .c(s_51_0), .d(t_400), .cin(t_403), .o(t_404), .co(t_405), .cout(t_406));
compressor_4_2 u2_147(.a(s_51_7), .b(s_51_6), .c(s_51_5), .d(s_51_4), .cin(s_51_3), .o(t_407), .co(t_408), .cout(t_409));
compressor_4_2 u2_148(.a(s_52_2), .b(s_52_1), .c(s_52_0), .d(t_406), .cin(t_409), .o(t_410), .co(t_411), .cout(t_412));
compressor_3_2 u1_149(.a(s_52_5), .b(s_52_4), .cin(s_52_3), .o(t_413), .cout(t_414));
compressor_4_2 u2_150(.a(s_53_2), .b(s_53_1), .c(s_53_0), .d(t_412), .cin(t_414), .o(t_415), .co(t_416), .cout(t_417));
compressor_3_2 u1_151(.a(s_53_5), .b(s_53_4), .cin(s_53_3), .o(t_418), .cout(t_419));
compressor_4_2 u2_152(.a(s_54_2), .b(s_54_1), .c(s_54_0), .d(t_417), .cin(t_419), .o(t_420), .co(t_421), .cout(t_422));
compressor_3_2 u1_153(.a(s_54_5), .b(s_54_4), .cin(s_54_3), .o(t_423), .cout(t_424));
compressor_4_2 u2_154(.a(s_55_2), .b(s_55_1), .c(s_55_0), .d(t_422), .cin(t_424), .o(t_425), .co(t_426), .cout(t_427));
compressor_3_2 u1_155(.a(s_55_5), .b(s_55_4), .cin(s_55_3), .o(t_428), .cout(t_429));
compressor_4_2 u2_156(.a(s_56_2), .b(s_56_1), .c(s_56_0), .d(t_427), .cin(t_429), .o(t_430), .co(t_431), .cout(t_432));
half_adder u0_157(.a(s_56_4), .b(s_56_3), .o(t_433), .cout(t_434));
compressor_4_2 u2_158(.a(s_57_2), .b(s_57_1), .c(s_57_0), .d(t_432), .cin(t_434), .o(t_435), .co(t_436), .cout(t_437));
half_adder u0_159(.a(s_57_4), .b(s_57_3), .o(t_438), .cout(t_439));
compressor_4_2 u2_160(.a(s_58_2), .b(s_58_1), .c(s_58_0), .d(t_437), .cin(t_439), .o(t_440), .co(t_441), .cout(t_442));
compressor_4_2 u2_161(.a(s_59_3), .b(s_59_2), .c(s_59_1), .d(s_59_0), .cin(t_442), .o(t_443), .co(t_444), .cout(t_445));
compressor_3_2 u1_162(.a(s_60_1), .b(s_60_0), .cin(t_445), .o(t_446), .cout(t_447));
compressor_3_2 u1_163(.a(s_61_2), .b(s_61_1), .cin(s_61_0), .o(t_448), .cout(t_449));
half_adder u0_164(.a(s_62_1), .b(s_62_0), .o(t_450), .cout(t_451));
half_adder u0_165(.a(s_63_1), .b(s_63_0), .o(t_452), .cout());

/* u0_166 Output nets */
wire t_453,    t_454;
/* u0_167 Output nets */
wire t_455,    t_456;
/* u1_168 Output nets */
wire t_457,    t_458;
/* u0_169 Output nets */
wire t_459,    t_460;
/* u0_170 Output nets */
wire t_461,    t_462;
/* u1_171 Output nets */
wire t_463,    t_464;
/* u1_172 Output nets */
wire t_465,    t_466;
/* u2_173 Output nets */
wire t_467,    t_468,    t_469;
/* u1_174 Output nets */
wire t_470,    t_471;
/* u1_175 Output nets */
wire t_472,    t_473;
/* u2_176 Output nets */
wire t_474,    t_475,    t_476;
/* u2_177 Output nets */
wire t_477,    t_478,    t_479;
/* u2_178 Output nets */
wire t_480,    t_481,    t_482;
/* u2_179 Output nets */
wire t_483,    t_484,    t_485;
/* u2_180 Output nets */
wire t_486,    t_487,    t_488;
/* u2_181 Output nets */
wire t_489,    t_490,    t_491;
/* u0_182 Output nets */
wire t_492,    t_493;
/* u2_183 Output nets */
wire t_494,    t_495,    t_496;
/* u0_184 Output nets */
wire t_497,    t_498;
/* u2_185 Output nets */
wire t_499,    t_500,    t_501;
/* u0_186 Output nets */
wire t_502,    t_503;
/* u2_187 Output nets */
wire t_504,    t_505,    t_506;
/* u1_188 Output nets */
wire t_507,    t_508;
/* u2_189 Output nets */
wire t_509,    t_510,    t_511;
/* u1_190 Output nets */
wire t_512,    t_513;
/* u2_191 Output nets */
wire t_514,    t_515,    t_516;
/* u1_192 Output nets */
wire t_517,    t_518;
/* u2_193 Output nets */
wire t_519,    t_520,    t_521;
/* u1_194 Output nets */
wire t_522,    t_523;
/* u2_195 Output nets */
wire t_524,    t_525,    t_526;
/* u1_196 Output nets */
wire t_527,    t_528;
/* u2_197 Output nets */
wire t_529,    t_530,    t_531;
/* u2_198 Output nets */
wire t_532,    t_533,    t_534;
/* u2_199 Output nets */
wire t_535,    t_536,    t_537;
/* u1_200 Output nets */
wire t_538,    t_539;
/* u2_201 Output nets */
wire t_540,    t_541,    t_542;
/* u1_202 Output nets */
wire t_543,    t_544;
/* u2_203 Output nets */
wire t_545,    t_546,    t_547;
/* u2_204 Output nets */
wire t_548,    t_549,    t_550;
/* u2_205 Output nets */
wire t_551,    t_552,    t_553;
/* u2_206 Output nets */
wire t_554,    t_555,    t_556;
/* u2_207 Output nets */
wire t_557,    t_558,    t_559;
/* u2_208 Output nets */
wire t_560,    t_561,    t_562;
/* u2_209 Output nets */
wire t_563,    t_564,    t_565;
/* u2_210 Output nets */
wire t_566,    t_567,    t_568;
/* u2_211 Output nets */
wire t_569,    t_570,    t_571;
/* u2_212 Output nets */
wire t_572,    t_573,    t_574;
/* u2_213 Output nets */
wire t_575,    t_576,    t_577;
/* u2_214 Output nets */
wire t_578,    t_579,    t_580;
/* u2_215 Output nets */
wire t_581,    t_582,    t_583;
/* u2_216 Output nets */
wire t_584,    t_585,    t_586;
/* u2_217 Output nets */
wire t_587,    t_588,    t_589;
/* u2_218 Output nets */
wire t_590,    t_591,    t_592;
/* u2_219 Output nets */
wire t_593,    t_594,    t_595;
/* u2_220 Output nets */
wire t_596,    t_597,    t_598;
/* u2_221 Output nets */
wire t_599,    t_600,    t_601;
/* u1_222 Output nets */
wire t_602,    t_603;
/* u2_223 Output nets */
wire t_604,    t_605,    t_606;
/* u1_224 Output nets */
wire t_607,    t_608;
/* u2_225 Output nets */
wire t_609,    t_610,    t_611;
/* u1_226 Output nets */
wire t_612,    t_613;
/* u2_227 Output nets */
wire t_614,    t_615,    t_616;
/* u1_228 Output nets */
wire t_617,    t_618;
/* u2_229 Output nets */
wire t_619,    t_620,    t_621;
/* u1_230 Output nets */
wire t_622,    t_623;
/* u2_231 Output nets */
wire t_624,    t_625,    t_626;
/* u1_232 Output nets */
wire t_627,    t_628;
/* u2_233 Output nets */
wire t_629,    t_630,    t_631;
/* u1_234 Output nets */
wire t_632,    t_633;
/* u2_235 Output nets */
wire t_634,    t_635,    t_636;
/* u1_236 Output nets */
wire t_637,    t_638;
/* u2_237 Output nets */
wire t_639,    t_640,    t_641;
/* u0_238 Output nets */
wire t_642,    t_643;
/* u2_239 Output nets */
wire t_644,    t_645,    t_646;
/* u0_240 Output nets */
wire t_647,    t_648;
/* u2_241 Output nets */
wire t_649,    t_650,    t_651;
/* u0_242 Output nets */
wire t_652,    t_653;
/* u2_243 Output nets */
wire t_654,    t_655,    t_656;
/* u0_244 Output nets */
wire t_657,    t_658;
/* u2_245 Output nets */
wire t_659,    t_660,    t_661;
/* u0_246 Output nets */
wire t_662,    t_663;
/* u2_247 Output nets */
wire t_664,    t_665,    t_666;
/* u2_248 Output nets */
wire t_667,    t_668,    t_669;
/* u2_249 Output nets */
wire t_670,    t_671,    t_672;
/* u1_250 Output nets */
wire t_673,    t_674;
/* u1_251 Output nets */
wire t_675,    t_676;
/* u1_252 Output nets */
wire t_677,    t_678;
/* u1_253 Output nets */
wire t_679,    t_680;
/* u1_254 Output nets */
wire t_681,    t_682;
/* u0_255 Output nets */
wire t_683,    t_684;
/* u1_256 Output nets */
wire t_685,    t_686;
/* u0_257 Output nets */
wire t_687,    t_688;
/* u0_258 Output nets */
wire t_689,    t_690;
/* u0_259 Output nets */
wire t_691;

/* compress stage 2 */
half_adder u0_166(.a(t_1), .b(s_1_0), .o(t_453), .cout(t_454));
half_adder u0_167(.a(t_3), .b(t_4), .o(t_455), .cout(t_456));
compressor_3_2 u1_168(.a(t_7), .b(t_9), .cin(s_5_2), .o(t_457), .cout(t_458));
half_adder u0_169(.a(t_10), .b(t_11), .o(t_459), .cout(t_460));
half_adder u0_170(.a(t_12), .b(t_14), .o(t_461), .cout(t_462));
compressor_3_2 u1_171(.a(t_15), .b(t_20), .cin(t_17), .o(t_463), .cout(t_464));
compressor_3_2 u1_172(.a(t_18), .b(t_25), .cin(t_22), .o(t_465), .cout(t_466));
compressor_4_2 u2_173(.a(t_23), .b(t_30), .c(t_27), .d(s_10_6), .cin(t_466), .o(t_467), .co(t_468), .cout(t_469));
compressor_3_2 u1_174(.a(t_35), .b(t_32), .cin(t_469), .o(t_470), .cout(t_471));
compressor_3_2 u1_175(.a(t_33), .b(t_40), .cin(t_37), .o(t_472), .cout(t_473));
compressor_4_2 u2_176(.a(t_38), .b(t_46), .c(t_43), .d(s_13_6), .cin(t_473), .o(t_474), .co(t_475), .cout(t_476));
compressor_4_2 u2_177(.a(t_44), .b(t_51), .c(t_48), .d(s_14_8), .cin(t_476), .o(t_477), .co(t_478), .cout(t_479));
compressor_4_2 u2_178(.a(t_52), .b(t_49), .c(t_57), .d(t_54), .cin(t_479), .o(t_480), .co(t_481), .cout(t_482));
compressor_4_2 u2_179(.a(t_55), .b(t_66), .c(t_63), .d(t_60), .cin(t_482), .o(t_483), .co(t_484), .cout(t_485));
compressor_4_2 u2_180(.a(t_61), .b(t_74), .c(t_71), .d(t_68), .cin(t_485), .o(t_486), .co(t_487), .cout(t_488));
compressor_4_2 u2_181(.a(t_82), .b(t_79), .c(t_76), .d(s_18_10), .cin(t_488), .o(t_489), .co(t_490), .cout(t_491));
half_adder u0_182(.a(t_72), .b(t_69), .o(t_492), .cout(t_493));
compressor_4_2 u2_183(.a(t_90), .b(t_87), .c(t_84), .d(t_491), .cin(t_493), .o(t_494), .co(t_495), .cout(t_496));
half_adder u0_184(.a(t_80), .b(t_77), .o(t_497), .cout(t_498));
compressor_4_2 u2_185(.a(t_98), .b(t_95), .c(t_92), .d(t_496), .cin(t_498), .o(t_499), .co(t_500), .cout(t_501));
half_adder u0_186(.a(t_88), .b(t_85), .o(t_502), .cout(t_503));
compressor_4_2 u2_187(.a(t_104), .b(t_101), .c(s_21_10), .d(t_501), .cin(t_503), .o(t_504), .co(t_505), .cout(t_506));
compressor_3_2 u1_188(.a(t_96), .b(t_93), .cin(t_107), .o(t_507), .cout(t_508));
compressor_4_2 u2_189(.a(t_112), .b(t_109), .c(s_22_12), .d(t_506), .cin(t_508), .o(t_509), .co(t_510), .cout(t_511));
compressor_3_2 u1_190(.a(t_105), .b(t_102), .cin(t_115), .o(t_512), .cout(t_513));
compressor_4_2 u2_191(.a(t_124), .b(t_121), .c(t_118), .d(t_511), .cin(t_513), .o(t_514), .co(t_515), .cout(t_516));
compressor_3_2 u1_192(.a(t_116), .b(t_113), .cin(t_110), .o(t_517), .cout(t_518));
compressor_4_2 u2_193(.a(t_133), .b(t_130), .c(t_127), .d(t_516), .cin(t_518), .o(t_519), .co(t_520), .cout(t_521));
compressor_3_2 u1_194(.a(t_122), .b(t_119), .cin(t_136), .o(t_522), .cout(t_523));
compressor_4_2 u2_195(.a(t_144), .b(t_141), .c(t_138), .d(t_521), .cin(t_523), .o(t_524), .co(t_525), .cout(t_526));
compressor_3_2 u1_196(.a(t_131), .b(t_128), .cin(t_147), .o(t_527), .cout(t_528));
compressor_4_2 u2_197(.a(t_152), .b(t_149), .c(s_26_14), .d(t_526), .cin(t_528), .o(t_529), .co(t_530), .cout(t_531));
compressor_4_2 u2_198(.a(t_145), .b(t_142), .c(t_139), .d(t_158), .cin(t_155), .o(t_532), .co(t_533), .cout(t_534));
compressor_4_2 u2_199(.a(t_166), .b(t_163), .c(t_160), .d(t_531), .cin(t_534), .o(t_535), .co(t_536), .cout(t_537));
compressor_3_2 u1_200(.a(t_153), .b(t_150), .cin(t_169), .o(t_538), .cout(t_539));
compressor_4_2 u2_201(.a(t_177), .b(t_174), .c(t_171), .d(t_537), .cin(t_539), .o(t_540), .co(t_541), .cout(t_542));
compressor_3_2 u1_202(.a(t_164), .b(t_161), .cin(t_180), .o(t_543), .cout(t_544));
compressor_4_2 u2_203(.a(t_186), .b(t_183), .c(s_29_14), .d(t_542), .cin(t_544), .o(t_545), .co(t_546), .cout(t_547));
compressor_4_2 u2_204(.a(t_178), .b(t_175), .c(t_172), .d(t_192), .cin(t_189), .o(t_548), .co(t_549), .cout(t_550));
compressor_4_2 u2_205(.a(t_197), .b(t_194), .c(s_30_16), .d(t_547), .cin(t_550), .o(t_551), .co(t_552), .cout(t_553));
compressor_4_2 u2_206(.a(t_190), .b(t_187), .c(t_184), .d(t_203), .cin(t_200), .o(t_554), .co(t_555), .cout(t_556));
compressor_4_2 u2_207(.a(t_212), .b(t_209), .c(t_206), .d(t_553), .cin(t_556), .o(t_557), .co(t_558), .cout(t_559));
compressor_4_2 u2_208(.a(t_204), .b(t_201), .c(t_198), .d(t_195), .cin(t_215), .o(t_560), .co(t_561), .cout(t_562));
compressor_4_2 u2_209(.a(t_221), .b(t_218), .c(s_32_16), .d(t_559), .cin(t_562), .o(t_563), .co(t_564), .cout(t_565));
compressor_4_2 u2_210(.a(t_213), .b(t_210), .c(t_207), .d(t_227), .cin(t_224), .o(t_566), .co(t_567), .cout(t_568));
compressor_4_2 u2_211(.a(t_233), .b(t_230), .c(s_33_16), .d(t_565), .cin(t_568), .o(t_569), .co(t_570), .cout(t_571));
compressor_4_2 u2_212(.a(t_225), .b(t_222), .c(t_219), .d(t_239), .cin(t_236), .o(t_572), .co(t_573), .cout(t_574));
compressor_4_2 u2_213(.a(t_248), .b(t_245), .c(t_242), .d(t_571), .cin(t_574), .o(t_575), .co(t_576), .cout(t_577));
compressor_4_2 u2_214(.a(t_240), .b(t_237), .c(t_234), .d(t_231), .cin(t_251), .o(t_578), .co(t_579), .cout(t_580));
compressor_4_2 u2_215(.a(t_260), .b(t_257), .c(t_254), .d(t_577), .cin(t_580), .o(t_581), .co(t_582), .cout(t_583));
compressor_4_2 u2_216(.a(t_252), .b(t_249), .c(t_246), .d(t_243), .cin(t_263), .o(t_584), .co(t_585), .cout(t_586));
compressor_4_2 u2_217(.a(t_269), .b(t_266), .c(s_36_14), .d(t_583), .cin(t_586), .o(t_587), .co(t_588), .cout(t_589));
compressor_4_2 u2_218(.a(t_261), .b(t_258), .c(t_255), .d(t_275), .cin(t_272), .o(t_590), .co(t_591), .cout(t_592));
compressor_4_2 u2_219(.a(t_280), .b(t_277), .c(s_37_14), .d(t_589), .cin(t_592), .o(t_593), .co(t_594), .cout(t_595));
compressor_4_2 u2_220(.a(t_273), .b(t_270), .c(t_267), .d(t_286), .cin(t_283), .o(t_596), .co(t_597), .cout(t_598));
compressor_4_2 u2_221(.a(t_294), .b(t_291), .c(t_288), .d(t_595), .cin(t_598), .o(t_599), .co(t_600), .cout(t_601));
compressor_3_2 u1_222(.a(t_281), .b(t_278), .cin(t_297), .o(t_602), .cout(t_603));
compressor_4_2 u2_223(.a(t_305), .b(t_302), .c(t_299), .d(t_601), .cin(t_603), .o(t_604), .co(t_605), .cout(t_606));
compressor_3_2 u1_224(.a(t_292), .b(t_289), .cin(t_308), .o(t_607), .cout(t_608));
compressor_4_2 u2_225(.a(t_316), .b(t_313), .c(t_310), .d(t_606), .cin(t_608), .o(t_609), .co(t_610), .cout(t_611));
compressor_3_2 u1_226(.a(t_303), .b(t_300), .cin(t_319), .o(t_612), .cout(t_613));
compressor_4_2 u2_227(.a(t_327), .b(t_324), .c(t_321), .d(t_611), .cin(t_613), .o(t_614), .co(t_615), .cout(t_616));
compressor_3_2 u1_228(.a(t_314), .b(t_311), .cin(t_330), .o(t_617), .cout(t_618));
compressor_4_2 u2_229(.a(t_335), .b(t_332), .c(s_42_11), .d(t_616), .cin(t_618), .o(t_619), .co(t_620), .cout(t_621));
compressor_3_2 u1_230(.a(t_325), .b(t_322), .cin(t_338), .o(t_622), .cout(t_623));
compressor_4_2 u2_231(.a(t_347), .b(t_344), .c(t_341), .d(t_621), .cin(t_623), .o(t_624), .co(t_625), .cout(t_626));
compressor_3_2 u1_232(.a(t_339), .b(t_336), .cin(t_333), .o(t_627), .cout(t_628));
compressor_4_2 u2_233(.a(t_353), .b(t_350), .c(s_44_10), .d(t_626), .cin(t_628), .o(t_629), .co(t_630), .cout(t_631));
compressor_3_2 u1_234(.a(t_345), .b(t_342), .cin(t_356), .o(t_632), .cout(t_633));
compressor_4_2 u2_235(.a(t_361), .b(t_358), .c(s_45_10), .d(t_631), .cin(t_633), .o(t_634), .co(t_635), .cout(t_636));
compressor_3_2 u1_236(.a(t_354), .b(t_351), .cin(t_364), .o(t_637), .cout(t_638));
compressor_4_2 u2_237(.a(t_372), .b(t_369), .c(t_366), .d(t_636), .cin(t_638), .o(t_639), .co(t_640), .cout(t_641));
half_adder u0_238(.a(t_362), .b(t_359), .o(t_642), .cout(t_643));
compressor_4_2 u2_239(.a(t_380), .b(t_377), .c(t_374), .d(t_641), .cin(t_643), .o(t_644), .co(t_645), .cout(t_646));
half_adder u0_240(.a(t_370), .b(t_367), .o(t_647), .cout(t_648));
compressor_4_2 u2_241(.a(t_388), .b(t_385), .c(t_382), .d(t_646), .cin(t_648), .o(t_649), .co(t_650), .cout(t_651));
half_adder u0_242(.a(t_378), .b(t_375), .o(t_652), .cout(t_653));
compressor_4_2 u2_243(.a(t_396), .b(t_393), .c(t_390), .d(t_651), .cin(t_653), .o(t_654), .co(t_655), .cout(t_656));
half_adder u0_244(.a(t_386), .b(t_383), .o(t_657), .cout(t_658));
compressor_4_2 u2_245(.a(t_401), .b(t_398), .c(s_50_7), .d(t_656), .cin(t_658), .o(t_659), .co(t_660), .cout(t_661));
half_adder u0_246(.a(t_394), .b(t_391), .o(t_662), .cout(t_663));
compressor_4_2 u2_247(.a(t_399), .b(t_407), .c(t_404), .d(t_661), .cin(t_663), .o(t_664), .co(t_665), .cout(t_666));
compressor_4_2 u2_248(.a(t_405), .b(t_413), .c(t_410), .d(s_52_6), .cin(t_666), .o(t_667), .co(t_668), .cout(t_669));
compressor_4_2 u2_249(.a(t_411), .b(t_418), .c(t_415), .d(s_53_6), .cin(t_669), .o(t_670), .co(t_671), .cout(t_672));
compressor_3_2 u1_250(.a(t_423), .b(t_420), .cin(t_672), .o(t_673), .cout(t_674));
compressor_3_2 u1_251(.a(t_421), .b(t_428), .cin(t_425), .o(t_675), .cout(t_676));
compressor_3_2 u1_252(.a(t_426), .b(t_433), .cin(t_430), .o(t_677), .cout(t_678));
compressor_3_2 u1_253(.a(t_431), .b(t_438), .cin(t_435), .o(t_679), .cout(t_680));
compressor_3_2 u1_254(.a(t_436), .b(t_440), .cin(s_58_3), .o(t_681), .cout(t_682));
half_adder u0_255(.a(t_441), .b(t_443), .o(t_683), .cout(t_684));
compressor_3_2 u1_256(.a(t_444), .b(t_446), .cin(s_60_2), .o(t_685), .cout(t_686));
half_adder u0_257(.a(t_447), .b(t_448), .o(t_687), .cout(t_688));
half_adder u0_258(.a(t_449), .b(t_450), .o(t_689), .cout(t_690));
half_adder u0_259(.a(t_451), .b(t_452), .o(t_691), .cout());

/* u0_260 Output nets */
wire t_692,    t_693;
/* u0_261 Output nets */
wire t_694,    t_695;
/* u0_262 Output nets */
wire t_696,    t_697;
/* u0_263 Output nets */
wire t_698,    t_699;
/* u0_264 Output nets */
wire t_700,    t_701;
/* u0_265 Output nets */
wire t_702,    t_703;
/* u1_266 Output nets */
wire t_704,    t_705;
/* u0_267 Output nets */
wire t_706,    t_707;
/* u0_268 Output nets */
wire t_708,    t_709;
/* u0_269 Output nets */
wire t_710,    t_711;
/* u0_270 Output nets */
wire t_712,    t_713;
/* u1_271 Output nets */
wire t_714,    t_715;
/* u1_272 Output nets */
wire t_716,    t_717;
/* u1_273 Output nets */
wire t_718,    t_719;
/* u1_274 Output nets */
wire t_720,    t_721;
/* u1_275 Output nets */
wire t_722,    t_723;
/* u2_276 Output nets */
wire t_724,    t_725,    t_726;
/* u1_277 Output nets */
wire t_727,    t_728;
/* u1_278 Output nets */
wire t_729,    t_730;
/* u2_279 Output nets */
wire t_731,    t_732,    t_733;
/* u2_280 Output nets */
wire t_734,    t_735,    t_736;
/* u1_281 Output nets */
wire t_737,    t_738;
/* u2_282 Output nets */
wire t_739,    t_740,    t_741;
/* u2_283 Output nets */
wire t_742,    t_743,    t_744;
/* u2_284 Output nets */
wire t_745,    t_746,    t_747;
/* u2_285 Output nets */
wire t_748,    t_749,    t_750;
/* u2_286 Output nets */
wire t_751,    t_752,    t_753;
/* u2_287 Output nets */
wire t_754,    t_755,    t_756;
/* u2_288 Output nets */
wire t_757,    t_758,    t_759;
/* u2_289 Output nets */
wire t_760,    t_761,    t_762;
/* u2_290 Output nets */
wire t_763,    t_764,    t_765;
/* u2_291 Output nets */
wire t_766,    t_767,    t_768;
/* u2_292 Output nets */
wire t_769,    t_770,    t_771;
/* u2_293 Output nets */
wire t_772,    t_773,    t_774;
/* u2_294 Output nets */
wire t_775,    t_776,    t_777;
/* u2_295 Output nets */
wire t_778,    t_779,    t_780;
/* u2_296 Output nets */
wire t_781,    t_782,    t_783;
/* u2_297 Output nets */
wire t_784,    t_785,    t_786;
/* u1_298 Output nets */
wire t_787,    t_788;
/* u1_299 Output nets */
wire t_789,    t_790;
/* u1_300 Output nets */
wire t_791,    t_792;
/* u1_301 Output nets */
wire t_793,    t_794;
/* u1_302 Output nets */
wire t_795,    t_796;
/* u1_303 Output nets */
wire t_797,    t_798;
/* u1_304 Output nets */
wire t_799,    t_800;
/* u1_305 Output nets */
wire t_801,    t_802;
/* u1_306 Output nets */
wire t_803,    t_804;
/* u1_307 Output nets */
wire t_805,    t_806;
/* u0_308 Output nets */
wire t_807,    t_808;
/* u1_309 Output nets */
wire t_809,    t_810;
/* u0_310 Output nets */
wire t_811,    t_812;
/* u0_311 Output nets */
wire t_813,    t_814;
/* u0_312 Output nets */
wire t_815,    t_816;
/* u0_313 Output nets */
wire t_817,    t_818;
/* u0_314 Output nets */
wire t_819,    t_820;
/* u0_315 Output nets */
wire t_821,    t_822;
/* u0_316 Output nets */
wire t_823,    t_824;
/* u0_317 Output nets */
wire t_825,    t_826;
/* u0_318 Output nets */
wire t_827;

/* compress stage 3 */
half_adder u0_260(.a(t_454), .b(t_2), .o(t_692), .cout(t_693));
half_adder u0_261(.a(t_456), .b(t_6), .o(t_694), .cout(t_695));
half_adder u0_262(.a(t_458), .b(t_459), .o(t_696), .cout(t_697));
half_adder u0_263(.a(t_460), .b(t_461), .o(t_698), .cout(t_699));
half_adder u0_264(.a(t_462), .b(t_463), .o(t_700), .cout(t_701));
half_adder u0_265(.a(t_464), .b(t_465), .o(t_702), .cout(t_703));
compressor_3_2 u1_266(.a(t_468), .b(t_470), .cin(t_28), .o(t_704), .cout(t_705));
half_adder u0_267(.a(t_471), .b(t_472), .o(t_706), .cout(t_707));
half_adder u0_268(.a(t_474), .b(t_41), .o(t_708), .cout(t_709));
half_adder u0_269(.a(t_475), .b(t_477), .o(t_710), .cout(t_711));
half_adder u0_270(.a(t_478), .b(t_480), .o(t_712), .cout(t_713));
compressor_3_2 u1_271(.a(t_481), .b(t_483), .cin(t_58), .o(t_714), .cout(t_715));
compressor_3_2 u1_272(.a(t_484), .b(t_486), .cin(t_64), .o(t_716), .cout(t_717));
compressor_3_2 u1_273(.a(t_487), .b(t_492), .cin(t_489), .o(t_718), .cout(t_719));
compressor_3_2 u1_274(.a(t_490), .b(t_497), .cin(t_494), .o(t_720), .cout(t_721));
compressor_3_2 u1_275(.a(t_495), .b(t_502), .cin(t_499), .o(t_722), .cout(t_723));
compressor_4_2 u2_276(.a(t_500), .b(t_507), .c(t_504), .d(t_99), .cin(t_723), .o(t_724), .co(t_725), .cout(t_726));
compressor_3_2 u1_277(.a(t_512), .b(t_509), .cin(t_726), .o(t_727), .cout(t_728));
compressor_3_2 u1_278(.a(t_510), .b(t_517), .cin(t_514), .o(t_729), .cout(t_730));
compressor_4_2 u2_279(.a(t_515), .b(t_522), .c(t_519), .d(t_125), .cin(t_730), .o(t_731), .co(t_732), .cout(t_733));
compressor_4_2 u2_280(.a(t_520), .b(t_527), .c(t_524), .d(t_134), .cin(t_733), .o(t_734), .co(t_735), .cout(t_736));
compressor_3_2 u1_281(.a(t_532), .b(t_529), .cin(t_736), .o(t_737), .cout(t_738));
compressor_4_2 u2_282(.a(t_533), .b(t_530), .c(t_538), .d(t_535), .cin(t_156), .o(t_739), .co(t_740), .cout(t_741));
compressor_4_2 u2_283(.a(t_536), .b(t_543), .c(t_540), .d(t_167), .cin(t_741), .o(t_742), .co(t_743), .cout(t_744));
compressor_4_2 u2_284(.a(t_541), .b(t_548), .c(t_545), .d(t_181), .cin(t_744), .o(t_745), .co(t_746), .cout(t_747));
compressor_4_2 u2_285(.a(t_549), .b(t_546), .c(t_554), .d(t_551), .cin(t_747), .o(t_748), .co(t_749), .cout(t_750));
compressor_4_2 u2_286(.a(t_555), .b(t_552), .c(t_560), .d(t_557), .cin(t_750), .o(t_751), .co(t_752), .cout(t_753));
compressor_4_2 u2_287(.a(t_558), .b(t_566), .c(t_563), .d(t_216), .cin(t_753), .o(t_754), .co(t_755), .cout(t_756));
compressor_4_2 u2_288(.a(t_564), .b(t_572), .c(t_569), .d(t_228), .cin(t_756), .o(t_757), .co(t_758), .cout(t_759));
compressor_4_2 u2_289(.a(t_573), .b(t_570), .c(t_578), .d(t_575), .cin(t_759), .o(t_760), .co(t_761), .cout(t_762));
compressor_4_2 u2_290(.a(t_579), .b(t_576), .c(t_584), .d(t_581), .cin(t_762), .o(t_763), .co(t_764), .cout(t_765));
compressor_4_2 u2_291(.a(t_582), .b(t_590), .c(t_587), .d(t_264), .cin(t_765), .o(t_766), .co(t_767), .cout(t_768));
compressor_4_2 u2_292(.a(t_591), .b(t_588), .c(t_596), .d(t_593), .cin(t_768), .o(t_769), .co(t_770), .cout(t_771));
compressor_4_2 u2_293(.a(t_594), .b(t_602), .c(t_599), .d(t_284), .cin(t_771), .o(t_772), .co(t_773), .cout(t_774));
compressor_4_2 u2_294(.a(t_600), .b(t_607), .c(t_604), .d(t_295), .cin(t_774), .o(t_775), .co(t_776), .cout(t_777));
compressor_4_2 u2_295(.a(t_605), .b(t_612), .c(t_609), .d(t_306), .cin(t_777), .o(t_778), .co(t_779), .cout(t_780));
compressor_4_2 u2_296(.a(t_610), .b(t_617), .c(t_614), .d(t_317), .cin(t_780), .o(t_781), .co(t_782), .cout(t_783));
compressor_4_2 u2_297(.a(t_615), .b(t_622), .c(t_619), .d(t_328), .cin(t_783), .o(t_784), .co(t_785), .cout(t_786));
compressor_3_2 u1_298(.a(t_627), .b(t_624), .cin(t_786), .o(t_787), .cout(t_788));
compressor_3_2 u1_299(.a(t_632), .b(t_629), .cin(t_348), .o(t_789), .cout(t_790));
compressor_3_2 u1_300(.a(t_630), .b(t_637), .cin(t_634), .o(t_791), .cout(t_792));
compressor_3_2 u1_301(.a(t_635), .b(t_642), .cin(t_639), .o(t_793), .cout(t_794));
compressor_3_2 u1_302(.a(t_640), .b(t_647), .cin(t_644), .o(t_795), .cout(t_796));
compressor_3_2 u1_303(.a(t_645), .b(t_652), .cin(t_649), .o(t_797), .cout(t_798));
compressor_3_2 u1_304(.a(t_650), .b(t_657), .cin(t_654), .o(t_799), .cout(t_800));
compressor_3_2 u1_305(.a(t_655), .b(t_662), .cin(t_659), .o(t_801), .cout(t_802));
compressor_3_2 u1_306(.a(t_660), .b(t_664), .cin(t_402), .o(t_803), .cout(t_804));
compressor_3_2 u1_307(.a(t_665), .b(t_667), .cin(t_408), .o(t_805), .cout(t_806));
half_adder u0_308(.a(t_668), .b(t_670), .o(t_807), .cout(t_808));
compressor_3_2 u1_309(.a(t_671), .b(t_673), .cin(t_416), .o(t_809), .cout(t_810));
half_adder u0_310(.a(t_674), .b(t_675), .o(t_811), .cout(t_812));
half_adder u0_311(.a(t_676), .b(t_677), .o(t_813), .cout(t_814));
half_adder u0_312(.a(t_678), .b(t_679), .o(t_815), .cout(t_816));
half_adder u0_313(.a(t_680), .b(t_681), .o(t_817), .cout(t_818));
half_adder u0_314(.a(t_682), .b(t_683), .o(t_819), .cout(t_820));
half_adder u0_315(.a(t_684), .b(t_685), .o(t_821), .cout(t_822));
half_adder u0_316(.a(t_686), .b(t_687), .o(t_823), .cout(t_824));
half_adder u0_317(.a(t_688), .b(t_689), .o(t_825), .cout(t_826));
half_adder u0_318(.a(t_690), .b(t_691), .o(t_827), .cout());

/* u0_319 Output nets */
wire t_828,    t_829;
/* u0_320 Output nets */
wire t_830,    t_831;
/* u0_321 Output nets */
wire t_832,    t_833;
/* u0_322 Output nets */
wire t_834,    t_835;
/* u0_323 Output nets */
wire t_836,    t_837;
/* u0_324 Output nets */
wire t_838,    t_839;
/* u0_325 Output nets */
wire t_840,    t_841;
/* u0_326 Output nets */
wire t_842,    t_843;
/* u0_327 Output nets */
wire t_844,    t_845;
/* u0_328 Output nets */
wire t_846,    t_847;
/* u0_329 Output nets */
wire t_848,    t_849;
/* u0_330 Output nets */
wire t_850,    t_851;
/* u0_331 Output nets */
wire t_852,    t_853;
/* u0_332 Output nets */
wire t_854,    t_855;
/* u0_333 Output nets */
wire t_856,    t_857;
/* u1_334 Output nets */
wire t_858,    t_859;
/* u0_335 Output nets */
wire t_860,    t_861;
/* u0_336 Output nets */
wire t_862,    t_863;
/* u1_337 Output nets */
wire t_864,    t_865;
/* u0_338 Output nets */
wire t_866,    t_867;
/* u0_339 Output nets */
wire t_868,    t_869;
/* u0_340 Output nets */
wire t_870,    t_871;
/* u0_341 Output nets */
wire t_872,    t_873;
/* u0_342 Output nets */
wire t_874,    t_875;
/* u1_343 Output nets */
wire t_876,    t_877;
/* u1_344 Output nets */
wire t_878,    t_879;
/* u0_345 Output nets */
wire t_880,    t_881;
/* u0_346 Output nets */
wire t_882,    t_883;
/* u1_347 Output nets */
wire t_884,    t_885;
/* u0_348 Output nets */
wire t_886,    t_887;
/* u1_349 Output nets */
wire t_888,    t_889;
/* u0_350 Output nets */
wire t_890,    t_891;
/* u0_351 Output nets */
wire t_892,    t_893;
/* u0_352 Output nets */
wire t_894,    t_895;
/* u0_353 Output nets */
wire t_896,    t_897;
/* u1_354 Output nets */
wire t_898,    t_899;
/* u1_355 Output nets */
wire t_900,    t_901;
/* u0_356 Output nets */
wire t_902,    t_903;
/* u0_357 Output nets */
wire t_904,    t_905;
/* u0_358 Output nets */
wire t_906,    t_907;
/* u0_359 Output nets */
wire t_908,    t_909;
/* u0_360 Output nets */
wire t_910,    t_911;
/* u0_361 Output nets */
wire t_912,    t_913;
/* u0_362 Output nets */
wire t_914,    t_915;
/* u0_363 Output nets */
wire t_916,    t_917;
/* u0_364 Output nets */
wire t_918,    t_919;
/* u0_365 Output nets */
wire t_920,    t_921;
/* u0_366 Output nets */
wire t_922,    t_923;
/* u0_367 Output nets */
wire t_924,    t_925;
/* u0_368 Output nets */
wire t_926,    t_927;
/* u0_369 Output nets */
wire t_928,    t_929;
/* u0_370 Output nets */
wire t_930,    t_931;
/* u0_371 Output nets */
wire t_932,    t_933;
/* u0_372 Output nets */
wire t_934,    t_935;
/* u0_373 Output nets */
wire t_936,    t_937;
/* u0_374 Output nets */
wire t_938;

/* compress stage 4 */
half_adder u0_319(.a(t_693), .b(t_455), .o(t_828), .cout(t_829));
half_adder u0_320(.a(t_695), .b(t_457), .o(t_830), .cout(t_831));
half_adder u0_321(.a(t_697), .b(t_698), .o(t_832), .cout(t_833));
half_adder u0_322(.a(t_699), .b(t_700), .o(t_834), .cout(t_835));
half_adder u0_323(.a(t_701), .b(t_702), .o(t_836), .cout(t_837));
half_adder u0_324(.a(t_703), .b(t_467), .o(t_838), .cout(t_839));
half_adder u0_325(.a(t_705), .b(t_706), .o(t_840), .cout(t_841));
half_adder u0_326(.a(t_707), .b(t_708), .o(t_842), .cout(t_843));
half_adder u0_327(.a(t_709), .b(t_710), .o(t_844), .cout(t_845));
half_adder u0_328(.a(t_711), .b(t_712), .o(t_846), .cout(t_847));
half_adder u0_329(.a(t_713), .b(t_714), .o(t_848), .cout(t_849));
half_adder u0_330(.a(t_715), .b(t_716), .o(t_850), .cout(t_851));
half_adder u0_331(.a(t_717), .b(t_718), .o(t_852), .cout(t_853));
half_adder u0_332(.a(t_719), .b(t_720), .o(t_854), .cout(t_855));
half_adder u0_333(.a(t_721), .b(t_722), .o(t_856), .cout(t_857));
compressor_3_2 u1_334(.a(t_725), .b(t_727), .cin(t_505), .o(t_858), .cout(t_859));
half_adder u0_335(.a(t_728), .b(t_729), .o(t_860), .cout(t_861));
half_adder u0_336(.a(t_732), .b(t_734), .o(t_862), .cout(t_863));
compressor_3_2 u1_337(.a(t_735), .b(t_737), .cin(t_525), .o(t_864), .cout(t_865));
half_adder u0_338(.a(t_738), .b(t_739), .o(t_866), .cout(t_867));
half_adder u0_339(.a(t_740), .b(t_742), .o(t_868), .cout(t_869));
half_adder u0_340(.a(t_743), .b(t_745), .o(t_870), .cout(t_871));
half_adder u0_341(.a(t_746), .b(t_748), .o(t_872), .cout(t_873));
half_adder u0_342(.a(t_749), .b(t_751), .o(t_874), .cout(t_875));
compressor_3_2 u1_343(.a(t_752), .b(t_754), .cin(t_561), .o(t_876), .cout(t_877));
compressor_3_2 u1_344(.a(t_755), .b(t_757), .cin(t_567), .o(t_878), .cout(t_879));
half_adder u0_345(.a(t_758), .b(t_760), .o(t_880), .cout(t_881));
half_adder u0_346(.a(t_761), .b(t_763), .o(t_882), .cout(t_883));
compressor_3_2 u1_347(.a(t_764), .b(t_766), .cin(t_585), .o(t_884), .cout(t_885));
half_adder u0_348(.a(t_767), .b(t_769), .o(t_886), .cout(t_887));
compressor_3_2 u1_349(.a(t_770), .b(t_772), .cin(t_597), .o(t_888), .cout(t_889));
half_adder u0_350(.a(t_773), .b(t_775), .o(t_890), .cout(t_891));
half_adder u0_351(.a(t_776), .b(t_778), .o(t_892), .cout(t_893));
half_adder u0_352(.a(t_779), .b(t_781), .o(t_894), .cout(t_895));
half_adder u0_353(.a(t_782), .b(t_784), .o(t_896), .cout(t_897));
compressor_3_2 u1_354(.a(t_785), .b(t_787), .cin(t_620), .o(t_898), .cout(t_899));
compressor_3_2 u1_355(.a(t_788), .b(t_789), .cin(t_625), .o(t_900), .cout(t_901));
half_adder u0_356(.a(t_790), .b(t_791), .o(t_902), .cout(t_903));
half_adder u0_357(.a(t_792), .b(t_793), .o(t_904), .cout(t_905));
half_adder u0_358(.a(t_794), .b(t_795), .o(t_906), .cout(t_907));
half_adder u0_359(.a(t_796), .b(t_797), .o(t_908), .cout(t_909));
half_adder u0_360(.a(t_798), .b(t_799), .o(t_910), .cout(t_911));
half_adder u0_361(.a(t_800), .b(t_801), .o(t_912), .cout(t_913));
half_adder u0_362(.a(t_802), .b(t_803), .o(t_914), .cout(t_915));
half_adder u0_363(.a(t_804), .b(t_805), .o(t_916), .cout(t_917));
half_adder u0_364(.a(t_806), .b(t_807), .o(t_918), .cout(t_919));
half_adder u0_365(.a(t_808), .b(t_809), .o(t_920), .cout(t_921));
half_adder u0_366(.a(t_810), .b(t_811), .o(t_922), .cout(t_923));
half_adder u0_367(.a(t_812), .b(t_813), .o(t_924), .cout(t_925));
half_adder u0_368(.a(t_814), .b(t_815), .o(t_926), .cout(t_927));
half_adder u0_369(.a(t_816), .b(t_817), .o(t_928), .cout(t_929));
half_adder u0_370(.a(t_818), .b(t_819), .o(t_930), .cout(t_931));
half_adder u0_371(.a(t_820), .b(t_821), .o(t_932), .cout(t_933));
half_adder u0_372(.a(t_822), .b(t_823), .o(t_934), .cout(t_935));
half_adder u0_373(.a(t_824), .b(t_825), .o(t_936), .cout(t_937));
half_adder u0_374(.a(t_826), .b(t_827), .o(t_938), .cout());

/* Output nets Compression result */
assign compress_a = {
   t_938,   t_936,   t_934,   t_932,
   t_930,   t_928,   t_926,   t_924,
   t_922,   t_920,   t_918,   t_916,
   t_914,   t_912,   t_910,   t_908,
   t_906,   t_904,   t_902,   t_900,
   t_898,   t_896,   t_894,   t_892,
   t_890,   t_888,   t_886,   t_884,
   t_882,   t_880,   t_878,   t_876,
   t_874,   t_872,   t_870,   t_868,
   t_866,   t_864,   t_862,   t_731,
   t_860,   t_858,   t_724,   t_856,
   t_854,   t_852,   t_850,   t_848,
   t_846,   t_844,   t_842,   t_840,
   t_704,   t_838,   t_836,   t_834,
   t_832,   t_696,   t_830,   t_694,
   t_828,   t_692,   t_453,     t_0
};
assign compress_b = {
   t_937,   t_935,   t_933,   t_931,
   t_929,   t_927,   t_925,   t_923,
   t_921,   t_919,   t_917,   t_915,
   t_913,   t_911,   t_909,   t_907,
   t_905,   t_903,   t_901,   t_899,
   t_897,   t_895,   t_893,   t_891,
   t_889,   t_887,   t_885,   t_883,
   t_881,   t_879,   t_877,   t_875,
   t_873,   t_871,   t_869,   t_867,
   t_865,   t_863,    1'b0,   t_861,
   t_859,    1'b0,   t_857,   t_855,
   t_853,   t_851,   t_849,   t_847,
   t_845,   t_843,   t_841,    1'b0,
   t_839,   t_837,   t_835,   t_833,
    1'b0,   t_831,    1'b0,   t_829,
    1'b0,    1'b0,    1'b0,    1'b0
};

endmodule

/********************************************************************************/

module _64_wallace_tree(
//inputs
	partial_products,
	carry,
//outputs
	compress_a,
	compress_b
);

localparam width = 64;

input wire [(width+2)*(width/2+1)-1:0] partial_products;
input wire [width/2-1:0] carry;
output wire [2*width-1:0] compress_a;
output wire [2*width-1:0] compress_b;

/* Input nets */
wire    s_0_0,    s_0_1,    s_1_0,    s_2_0,    s_2_1,    s_2_2;
wire    s_3_0,    s_3_1,    s_4_0,    s_4_1,    s_4_2,    s_4_3;
wire    s_5_0,    s_5_1,    s_5_2,    s_6_0,    s_6_1,    s_6_2;
wire    s_6_3,    s_6_4,    s_7_0,    s_7_1,    s_7_2,    s_7_3;
wire    s_8_0,    s_8_1,    s_8_2,    s_8_3,    s_8_4,    s_8_5;
wire    s_9_0,    s_9_1,    s_9_2,    s_9_3,    s_9_4,   s_10_0;
wire   s_10_1,   s_10_2,   s_10_3,   s_10_4,   s_10_5,   s_10_6;
wire   s_11_0,   s_11_1,   s_11_2,   s_11_3,   s_11_4,   s_11_5;
wire   s_12_0,   s_12_1,   s_12_2,   s_12_3,   s_12_4,   s_12_5;
wire   s_12_6,   s_12_7,   s_13_0,   s_13_1,   s_13_2,   s_13_3;
wire   s_13_4,   s_13_5,   s_13_6,   s_14_0,   s_14_1,   s_14_2;
wire   s_14_3,   s_14_4,   s_14_5,   s_14_6,   s_14_7,   s_14_8;
wire   s_15_0,   s_15_1,   s_15_2,   s_15_3,   s_15_4,   s_15_5;
wire   s_15_6,   s_15_7,   s_16_0,   s_16_1,   s_16_2,   s_16_3;
wire   s_16_4,   s_16_5,   s_16_6,   s_16_7,   s_16_8,   s_16_9;
wire   s_17_0,   s_17_1,   s_17_2,   s_17_3,   s_17_4,   s_17_5;
wire   s_17_6,   s_17_7,   s_17_8,   s_18_0,   s_18_1,   s_18_2;
wire   s_18_3,   s_18_4,   s_18_5,   s_18_6,   s_18_7,   s_18_8;
wire   s_18_9,  s_18_10,   s_19_0,   s_19_1,   s_19_2,   s_19_3;
wire   s_19_4,   s_19_5,   s_19_6,   s_19_7,   s_19_8,   s_19_9;
wire   s_20_0,   s_20_1,   s_20_2,   s_20_3,   s_20_4,   s_20_5;
wire   s_20_6,   s_20_7,   s_20_8,   s_20_9,  s_20_10,  s_20_11;
wire   s_21_0,   s_21_1,   s_21_2,   s_21_3,   s_21_4,   s_21_5;
wire   s_21_6,   s_21_7,   s_21_8,   s_21_9,  s_21_10,   s_22_0;
wire   s_22_1,   s_22_2,   s_22_3,   s_22_4,   s_22_5,   s_22_6;
wire   s_22_7,   s_22_8,   s_22_9,  s_22_10,  s_22_11,  s_22_12;
wire   s_23_0,   s_23_1,   s_23_2,   s_23_3,   s_23_4,   s_23_5;
wire   s_23_6,   s_23_7,   s_23_8,   s_23_9,  s_23_10,  s_23_11;
wire   s_24_0,   s_24_1,   s_24_2,   s_24_3,   s_24_4,   s_24_5;
wire   s_24_6,   s_24_7,   s_24_8,   s_24_9,  s_24_10,  s_24_11;
wire  s_24_12,  s_24_13,   s_25_0,   s_25_1,   s_25_2,   s_25_3;
wire   s_25_4,   s_25_5,   s_25_6,   s_25_7,   s_25_8,   s_25_9;
wire  s_25_10,  s_25_11,  s_25_12,   s_26_0,   s_26_1,   s_26_2;
wire   s_26_3,   s_26_4,   s_26_5,   s_26_6,   s_26_7,   s_26_8;
wire   s_26_9,  s_26_10,  s_26_11,  s_26_12,  s_26_13,  s_26_14;
wire   s_27_0,   s_27_1,   s_27_2,   s_27_3,   s_27_4,   s_27_5;
wire   s_27_6,   s_27_7,   s_27_8,   s_27_9,  s_27_10,  s_27_11;
wire  s_27_12,  s_27_13,   s_28_0,   s_28_1,   s_28_2,   s_28_3;
wire   s_28_4,   s_28_5,   s_28_6,   s_28_7,   s_28_8,   s_28_9;
wire  s_28_10,  s_28_11,  s_28_12,  s_28_13,  s_28_14,  s_28_15;
wire   s_29_0,   s_29_1,   s_29_2,   s_29_3,   s_29_4,   s_29_5;
wire   s_29_6,   s_29_7,   s_29_8,   s_29_9,  s_29_10,  s_29_11;
wire  s_29_12,  s_29_13,  s_29_14,   s_30_0,   s_30_1,   s_30_2;
wire   s_30_3,   s_30_4,   s_30_5,   s_30_6,   s_30_7,   s_30_8;
wire   s_30_9,  s_30_10,  s_30_11,  s_30_12,  s_30_13,  s_30_14;
wire  s_30_15,  s_30_16,   s_31_0,   s_31_1,   s_31_2,   s_31_3;
wire   s_31_4,   s_31_5,   s_31_6,   s_31_7,   s_31_8,   s_31_9;
wire  s_31_10,  s_31_11,  s_31_12,  s_31_13,  s_31_14,  s_31_15;
wire   s_32_0,   s_32_1,   s_32_2,   s_32_3,   s_32_4,   s_32_5;
wire   s_32_6,   s_32_7,   s_32_8,   s_32_9,  s_32_10,  s_32_11;
wire  s_32_12,  s_32_13,  s_32_14,  s_32_15,  s_32_16,  s_32_17;
wire   s_33_0,   s_33_1,   s_33_2,   s_33_3,   s_33_4,   s_33_5;
wire   s_33_6,   s_33_7,   s_33_8,   s_33_9,  s_33_10,  s_33_11;
wire  s_33_12,  s_33_13,  s_33_14,  s_33_15,  s_33_16,   s_34_0;
wire   s_34_1,   s_34_2,   s_34_3,   s_34_4,   s_34_5,   s_34_6;
wire   s_34_7,   s_34_8,   s_34_9,  s_34_10,  s_34_11,  s_34_12;
wire  s_34_13,  s_34_14,  s_34_15,  s_34_16,  s_34_17,  s_34_18;
wire   s_35_0,   s_35_1,   s_35_2,   s_35_3,   s_35_4,   s_35_5;
wire   s_35_6,   s_35_7,   s_35_8,   s_35_9,  s_35_10,  s_35_11;
wire  s_35_12,  s_35_13,  s_35_14,  s_35_15,  s_35_16,  s_35_17;
wire   s_36_0,   s_36_1,   s_36_2,   s_36_3,   s_36_4,   s_36_5;
wire   s_36_6,   s_36_7,   s_36_8,   s_36_9,  s_36_10,  s_36_11;
wire  s_36_12,  s_36_13,  s_36_14,  s_36_15,  s_36_16,  s_36_17;
wire  s_36_18,  s_36_19,   s_37_0,   s_37_1,   s_37_2,   s_37_3;
wire   s_37_4,   s_37_5,   s_37_6,   s_37_7,   s_37_8,   s_37_9;
wire  s_37_10,  s_37_11,  s_37_12,  s_37_13,  s_37_14,  s_37_15;
wire  s_37_16,  s_37_17,  s_37_18,   s_38_0,   s_38_1,   s_38_2;
wire   s_38_3,   s_38_4,   s_38_5,   s_38_6,   s_38_7,   s_38_8;
wire   s_38_9,  s_38_10,  s_38_11,  s_38_12,  s_38_13,  s_38_14;
wire  s_38_15,  s_38_16,  s_38_17,  s_38_18,  s_38_19,  s_38_20;
wire   s_39_0,   s_39_1,   s_39_2,   s_39_3,   s_39_4,   s_39_5;
wire   s_39_6,   s_39_7,   s_39_8,   s_39_9,  s_39_10,  s_39_11;
wire  s_39_12,  s_39_13,  s_39_14,  s_39_15,  s_39_16,  s_39_17;
wire  s_39_18,  s_39_19,   s_40_0,   s_40_1,   s_40_2,   s_40_3;
wire   s_40_4,   s_40_5,   s_40_6,   s_40_7,   s_40_8,   s_40_9;
wire  s_40_10,  s_40_11,  s_40_12,  s_40_13,  s_40_14,  s_40_15;
wire  s_40_16,  s_40_17,  s_40_18,  s_40_19,  s_40_20,  s_40_21;
wire   s_41_0,   s_41_1,   s_41_2,   s_41_3,   s_41_4,   s_41_5;
wire   s_41_6,   s_41_7,   s_41_8,   s_41_9,  s_41_10,  s_41_11;
wire  s_41_12,  s_41_13,  s_41_14,  s_41_15,  s_41_16,  s_41_17;
wire  s_41_18,  s_41_19,  s_41_20,   s_42_0,   s_42_1,   s_42_2;
wire   s_42_3,   s_42_4,   s_42_5,   s_42_6,   s_42_7,   s_42_8;
wire   s_42_9,  s_42_10,  s_42_11,  s_42_12,  s_42_13,  s_42_14;
wire  s_42_15,  s_42_16,  s_42_17,  s_42_18,  s_42_19,  s_42_20;
wire  s_42_21,  s_42_22,   s_43_0,   s_43_1,   s_43_2,   s_43_3;
wire   s_43_4,   s_43_5,   s_43_6,   s_43_7,   s_43_8,   s_43_9;
wire  s_43_10,  s_43_11,  s_43_12,  s_43_13,  s_43_14,  s_43_15;
wire  s_43_16,  s_43_17,  s_43_18,  s_43_19,  s_43_20,  s_43_21;
wire   s_44_0,   s_44_1,   s_44_2,   s_44_3,   s_44_4,   s_44_5;
wire   s_44_6,   s_44_7,   s_44_8,   s_44_9,  s_44_10,  s_44_11;
wire  s_44_12,  s_44_13,  s_44_14,  s_44_15,  s_44_16,  s_44_17;
wire  s_44_18,  s_44_19,  s_44_20,  s_44_21,  s_44_22,  s_44_23;
wire   s_45_0,   s_45_1,   s_45_2,   s_45_3,   s_45_4,   s_45_5;
wire   s_45_6,   s_45_7,   s_45_8,   s_45_9,  s_45_10,  s_45_11;
wire  s_45_12,  s_45_13,  s_45_14,  s_45_15,  s_45_16,  s_45_17;
wire  s_45_18,  s_45_19,  s_45_20,  s_45_21,  s_45_22,   s_46_0;
wire   s_46_1,   s_46_2,   s_46_3,   s_46_4,   s_46_5,   s_46_6;
wire   s_46_7,   s_46_8,   s_46_9,  s_46_10,  s_46_11,  s_46_12;
wire  s_46_13,  s_46_14,  s_46_15,  s_46_16,  s_46_17,  s_46_18;
wire  s_46_19,  s_46_20,  s_46_21,  s_46_22,  s_46_23,  s_46_24;
wire   s_47_0,   s_47_1,   s_47_2,   s_47_3,   s_47_4,   s_47_5;
wire   s_47_6,   s_47_7,   s_47_8,   s_47_9,  s_47_10,  s_47_11;
wire  s_47_12,  s_47_13,  s_47_14,  s_47_15,  s_47_16,  s_47_17;
wire  s_47_18,  s_47_19,  s_47_20,  s_47_21,  s_47_22,  s_47_23;
wire   s_48_0,   s_48_1,   s_48_2,   s_48_3,   s_48_4,   s_48_5;
wire   s_48_6,   s_48_7,   s_48_8,   s_48_9,  s_48_10,  s_48_11;
wire  s_48_12,  s_48_13,  s_48_14,  s_48_15,  s_48_16,  s_48_17;
wire  s_48_18,  s_48_19,  s_48_20,  s_48_21,  s_48_22,  s_48_23;
wire  s_48_24,  s_48_25,   s_49_0,   s_49_1,   s_49_2,   s_49_3;
wire   s_49_4,   s_49_5,   s_49_6,   s_49_7,   s_49_8,   s_49_9;
wire  s_49_10,  s_49_11,  s_49_12,  s_49_13,  s_49_14,  s_49_15;
wire  s_49_16,  s_49_17,  s_49_18,  s_49_19,  s_49_20,  s_49_21;
wire  s_49_22,  s_49_23,  s_49_24,   s_50_0,   s_50_1,   s_50_2;
wire   s_50_3,   s_50_4,   s_50_5,   s_50_6,   s_50_7,   s_50_8;
wire   s_50_9,  s_50_10,  s_50_11,  s_50_12,  s_50_13,  s_50_14;
wire  s_50_15,  s_50_16,  s_50_17,  s_50_18,  s_50_19,  s_50_20;
wire  s_50_21,  s_50_22,  s_50_23,  s_50_24,  s_50_25,  s_50_26;
wire   s_51_0,   s_51_1,   s_51_2,   s_51_3,   s_51_4,   s_51_5;
wire   s_51_6,   s_51_7,   s_51_8,   s_51_9,  s_51_10,  s_51_11;
wire  s_51_12,  s_51_13,  s_51_14,  s_51_15,  s_51_16,  s_51_17;
wire  s_51_18,  s_51_19,  s_51_20,  s_51_21,  s_51_22,  s_51_23;
wire  s_51_24,  s_51_25,   s_52_0,   s_52_1,   s_52_2,   s_52_3;
wire   s_52_4,   s_52_5,   s_52_6,   s_52_7,   s_52_8,   s_52_9;
wire  s_52_10,  s_52_11,  s_52_12,  s_52_13,  s_52_14,  s_52_15;
wire  s_52_16,  s_52_17,  s_52_18,  s_52_19,  s_52_20,  s_52_21;
wire  s_52_22,  s_52_23,  s_52_24,  s_52_25,  s_52_26,  s_52_27;
wire   s_53_0,   s_53_1,   s_53_2,   s_53_3,   s_53_4,   s_53_5;
wire   s_53_6,   s_53_7,   s_53_8,   s_53_9,  s_53_10,  s_53_11;
wire  s_53_12,  s_53_13,  s_53_14,  s_53_15,  s_53_16,  s_53_17;
wire  s_53_18,  s_53_19,  s_53_20,  s_53_21,  s_53_22,  s_53_23;
wire  s_53_24,  s_53_25,  s_53_26,   s_54_0,   s_54_1,   s_54_2;
wire   s_54_3,   s_54_4,   s_54_5,   s_54_6,   s_54_7,   s_54_8;
wire   s_54_9,  s_54_10,  s_54_11,  s_54_12,  s_54_13,  s_54_14;
wire  s_54_15,  s_54_16,  s_54_17,  s_54_18,  s_54_19,  s_54_20;
wire  s_54_21,  s_54_22,  s_54_23,  s_54_24,  s_54_25,  s_54_26;
wire  s_54_27,  s_54_28,   s_55_0,   s_55_1,   s_55_2,   s_55_3;
wire   s_55_4,   s_55_5,   s_55_6,   s_55_7,   s_55_8,   s_55_9;
wire  s_55_10,  s_55_11,  s_55_12,  s_55_13,  s_55_14,  s_55_15;
wire  s_55_16,  s_55_17,  s_55_18,  s_55_19,  s_55_20,  s_55_21;
wire  s_55_22,  s_55_23,  s_55_24,  s_55_25,  s_55_26,  s_55_27;
wire   s_56_0,   s_56_1,   s_56_2,   s_56_3,   s_56_4,   s_56_5;
wire   s_56_6,   s_56_7,   s_56_8,   s_56_9,  s_56_10,  s_56_11;
wire  s_56_12,  s_56_13,  s_56_14,  s_56_15,  s_56_16,  s_56_17;
wire  s_56_18,  s_56_19,  s_56_20,  s_56_21,  s_56_22,  s_56_23;
wire  s_56_24,  s_56_25,  s_56_26,  s_56_27,  s_56_28,  s_56_29;
wire   s_57_0,   s_57_1,   s_57_2,   s_57_3,   s_57_4,   s_57_5;
wire   s_57_6,   s_57_7,   s_57_8,   s_57_9,  s_57_10,  s_57_11;
wire  s_57_12,  s_57_13,  s_57_14,  s_57_15,  s_57_16,  s_57_17;
wire  s_57_18,  s_57_19,  s_57_20,  s_57_21,  s_57_22,  s_57_23;
wire  s_57_24,  s_57_25,  s_57_26,  s_57_27,  s_57_28,   s_58_0;
wire   s_58_1,   s_58_2,   s_58_3,   s_58_4,   s_58_5,   s_58_6;
wire   s_58_7,   s_58_8,   s_58_9,  s_58_10,  s_58_11,  s_58_12;
wire  s_58_13,  s_58_14,  s_58_15,  s_58_16,  s_58_17,  s_58_18;
wire  s_58_19,  s_58_20,  s_58_21,  s_58_22,  s_58_23,  s_58_24;
wire  s_58_25,  s_58_26,  s_58_27,  s_58_28,  s_58_29,  s_58_30;
wire   s_59_0,   s_59_1,   s_59_2,   s_59_3,   s_59_4,   s_59_5;
wire   s_59_6,   s_59_7,   s_59_8,   s_59_9,  s_59_10,  s_59_11;
wire  s_59_12,  s_59_13,  s_59_14,  s_59_15,  s_59_16,  s_59_17;
wire  s_59_18,  s_59_19,  s_59_20,  s_59_21,  s_59_22,  s_59_23;
wire  s_59_24,  s_59_25,  s_59_26,  s_59_27,  s_59_28,  s_59_29;
wire   s_60_0,   s_60_1,   s_60_2,   s_60_3,   s_60_4,   s_60_5;
wire   s_60_6,   s_60_7,   s_60_8,   s_60_9,  s_60_10,  s_60_11;
wire  s_60_12,  s_60_13,  s_60_14,  s_60_15,  s_60_16,  s_60_17;
wire  s_60_18,  s_60_19,  s_60_20,  s_60_21,  s_60_22,  s_60_23;
wire  s_60_24,  s_60_25,  s_60_26,  s_60_27,  s_60_28,  s_60_29;
wire  s_60_30,  s_60_31,   s_61_0,   s_61_1,   s_61_2,   s_61_3;
wire   s_61_4,   s_61_5,   s_61_6,   s_61_7,   s_61_8,   s_61_9;
wire  s_61_10,  s_61_11,  s_61_12,  s_61_13,  s_61_14,  s_61_15;
wire  s_61_16,  s_61_17,  s_61_18,  s_61_19,  s_61_20,  s_61_21;
wire  s_61_22,  s_61_23,  s_61_24,  s_61_25,  s_61_26,  s_61_27;
wire  s_61_28,  s_61_29,  s_61_30,   s_62_0,   s_62_1,   s_62_2;
wire   s_62_3,   s_62_4,   s_62_5,   s_62_6,   s_62_7,   s_62_8;
wire   s_62_9,  s_62_10,  s_62_11,  s_62_12,  s_62_13,  s_62_14;
wire  s_62_15,  s_62_16,  s_62_17,  s_62_18,  s_62_19,  s_62_20;
wire  s_62_21,  s_62_22,  s_62_23,  s_62_24,  s_62_25,  s_62_26;
wire  s_62_27,  s_62_28,  s_62_29,  s_62_30,  s_62_31,  s_62_32;
wire   s_63_0,   s_63_1,   s_63_2,   s_63_3,   s_63_4,   s_63_5;
wire   s_63_6,   s_63_7,   s_63_8,   s_63_9,  s_63_10,  s_63_11;
wire  s_63_12,  s_63_13,  s_63_14,  s_63_15,  s_63_16,  s_63_17;
wire  s_63_18,  s_63_19,  s_63_20,  s_63_21,  s_63_22,  s_63_23;
wire  s_63_24,  s_63_25,  s_63_26,  s_63_27,  s_63_28,  s_63_29;
wire  s_63_30,  s_63_31,   s_64_0,   s_64_1,   s_64_2,   s_64_3;
wire   s_64_4,   s_64_5,   s_64_6,   s_64_7,   s_64_8,   s_64_9;
wire  s_64_10,  s_64_11,  s_64_12,  s_64_13,  s_64_14,  s_64_15;
wire  s_64_16,  s_64_17,  s_64_18,  s_64_19,  s_64_20,  s_64_21;
wire  s_64_22,  s_64_23,  s_64_24,  s_64_25,  s_64_26,  s_64_27;
wire  s_64_28,  s_64_29,  s_64_30,  s_64_31,  s_64_32,   s_65_0;
wire   s_65_1,   s_65_2,   s_65_3,   s_65_4,   s_65_5,   s_65_6;
wire   s_65_7,   s_65_8,   s_65_9,  s_65_10,  s_65_11,  s_65_12;
wire  s_65_13,  s_65_14,  s_65_15,  s_65_16,  s_65_17,  s_65_18;
wire  s_65_19,  s_65_20,  s_65_21,  s_65_22,  s_65_23,  s_65_24;
wire  s_65_25,  s_65_26,  s_65_27,  s_65_28,  s_65_29,  s_65_30;
wire  s_65_31,  s_65_32,   s_66_0,   s_66_1,   s_66_2,   s_66_3;
wire   s_66_4,   s_66_5,   s_66_6,   s_66_7,   s_66_8,   s_66_9;
wire  s_66_10,  s_66_11,  s_66_12,  s_66_13,  s_66_14,  s_66_15;
wire  s_66_16,  s_66_17,  s_66_18,  s_66_19,  s_66_20,  s_66_21;
wire  s_66_22,  s_66_23,  s_66_24,  s_66_25,  s_66_26,  s_66_27;
wire  s_66_28,  s_66_29,  s_66_30,  s_66_31,   s_67_0,   s_67_1;
wire   s_67_2,   s_67_3,   s_67_4,   s_67_5,   s_67_6,   s_67_7;
wire   s_67_8,   s_67_9,  s_67_10,  s_67_11,  s_67_12,  s_67_13;
wire  s_67_14,  s_67_15,  s_67_16,  s_67_17,  s_67_18,  s_67_19;
wire  s_67_20,  s_67_21,  s_67_22,  s_67_23,  s_67_24,  s_67_25;
wire  s_67_26,  s_67_27,  s_67_28,  s_67_29,  s_67_30,  s_67_31;
wire   s_68_0,   s_68_1,   s_68_2,   s_68_3,   s_68_4,   s_68_5;
wire   s_68_6,   s_68_7,   s_68_8,   s_68_9,  s_68_10,  s_68_11;
wire  s_68_12,  s_68_13,  s_68_14,  s_68_15,  s_68_16,  s_68_17;
wire  s_68_18,  s_68_19,  s_68_20,  s_68_21,  s_68_22,  s_68_23;
wire  s_68_24,  s_68_25,  s_68_26,  s_68_27,  s_68_28,  s_68_29;
wire  s_68_30,   s_69_0,   s_69_1,   s_69_2,   s_69_3,   s_69_4;
wire   s_69_5,   s_69_6,   s_69_7,   s_69_8,   s_69_9,  s_69_10;
wire  s_69_11,  s_69_12,  s_69_13,  s_69_14,  s_69_15,  s_69_16;
wire  s_69_17,  s_69_18,  s_69_19,  s_69_20,  s_69_21,  s_69_22;
wire  s_69_23,  s_69_24,  s_69_25,  s_69_26,  s_69_27,  s_69_28;
wire  s_69_29,  s_69_30,   s_70_0,   s_70_1,   s_70_2,   s_70_3;
wire   s_70_4,   s_70_5,   s_70_6,   s_70_7,   s_70_8,   s_70_9;
wire  s_70_10,  s_70_11,  s_70_12,  s_70_13,  s_70_14,  s_70_15;
wire  s_70_16,  s_70_17,  s_70_18,  s_70_19,  s_70_20,  s_70_21;
wire  s_70_22,  s_70_23,  s_70_24,  s_70_25,  s_70_26,  s_70_27;
wire  s_70_28,  s_70_29,   s_71_0,   s_71_1,   s_71_2,   s_71_3;
wire   s_71_4,   s_71_5,   s_71_6,   s_71_7,   s_71_8,   s_71_9;
wire  s_71_10,  s_71_11,  s_71_12,  s_71_13,  s_71_14,  s_71_15;
wire  s_71_16,  s_71_17,  s_71_18,  s_71_19,  s_71_20,  s_71_21;
wire  s_71_22,  s_71_23,  s_71_24,  s_71_25,  s_71_26,  s_71_27;
wire  s_71_28,  s_71_29,   s_72_0,   s_72_1,   s_72_2,   s_72_3;
wire   s_72_4,   s_72_5,   s_72_6,   s_72_7,   s_72_8,   s_72_9;
wire  s_72_10,  s_72_11,  s_72_12,  s_72_13,  s_72_14,  s_72_15;
wire  s_72_16,  s_72_17,  s_72_18,  s_72_19,  s_72_20,  s_72_21;
wire  s_72_22,  s_72_23,  s_72_24,  s_72_25,  s_72_26,  s_72_27;
wire  s_72_28,   s_73_0,   s_73_1,   s_73_2,   s_73_3,   s_73_4;
wire   s_73_5,   s_73_6,   s_73_7,   s_73_8,   s_73_9,  s_73_10;
wire  s_73_11,  s_73_12,  s_73_13,  s_73_14,  s_73_15,  s_73_16;
wire  s_73_17,  s_73_18,  s_73_19,  s_73_20,  s_73_21,  s_73_22;
wire  s_73_23,  s_73_24,  s_73_25,  s_73_26,  s_73_27,  s_73_28;
wire   s_74_0,   s_74_1,   s_74_2,   s_74_3,   s_74_4,   s_74_5;
wire   s_74_6,   s_74_7,   s_74_8,   s_74_9,  s_74_10,  s_74_11;
wire  s_74_12,  s_74_13,  s_74_14,  s_74_15,  s_74_16,  s_74_17;
wire  s_74_18,  s_74_19,  s_74_20,  s_74_21,  s_74_22,  s_74_23;
wire  s_74_24,  s_74_25,  s_74_26,  s_74_27,   s_75_0,   s_75_1;
wire   s_75_2,   s_75_3,   s_75_4,   s_75_5,   s_75_6,   s_75_7;
wire   s_75_8,   s_75_9,  s_75_10,  s_75_11,  s_75_12,  s_75_13;
wire  s_75_14,  s_75_15,  s_75_16,  s_75_17,  s_75_18,  s_75_19;
wire  s_75_20,  s_75_21,  s_75_22,  s_75_23,  s_75_24,  s_75_25;
wire  s_75_26,  s_75_27,   s_76_0,   s_76_1,   s_76_2,   s_76_3;
wire   s_76_4,   s_76_5,   s_76_6,   s_76_7,   s_76_8,   s_76_9;
wire  s_76_10,  s_76_11,  s_76_12,  s_76_13,  s_76_14,  s_76_15;
wire  s_76_16,  s_76_17,  s_76_18,  s_76_19,  s_76_20,  s_76_21;
wire  s_76_22,  s_76_23,  s_76_24,  s_76_25,  s_76_26,   s_77_0;
wire   s_77_1,   s_77_2,   s_77_3,   s_77_4,   s_77_5,   s_77_6;
wire   s_77_7,   s_77_8,   s_77_9,  s_77_10,  s_77_11,  s_77_12;
wire  s_77_13,  s_77_14,  s_77_15,  s_77_16,  s_77_17,  s_77_18;
wire  s_77_19,  s_77_20,  s_77_21,  s_77_22,  s_77_23,  s_77_24;
wire  s_77_25,  s_77_26,   s_78_0,   s_78_1,   s_78_2,   s_78_3;
wire   s_78_4,   s_78_5,   s_78_6,   s_78_7,   s_78_8,   s_78_9;
wire  s_78_10,  s_78_11,  s_78_12,  s_78_13,  s_78_14,  s_78_15;
wire  s_78_16,  s_78_17,  s_78_18,  s_78_19,  s_78_20,  s_78_21;
wire  s_78_22,  s_78_23,  s_78_24,  s_78_25,   s_79_0,   s_79_1;
wire   s_79_2,   s_79_3,   s_79_4,   s_79_5,   s_79_6,   s_79_7;
wire   s_79_8,   s_79_9,  s_79_10,  s_79_11,  s_79_12,  s_79_13;
wire  s_79_14,  s_79_15,  s_79_16,  s_79_17,  s_79_18,  s_79_19;
wire  s_79_20,  s_79_21,  s_79_22,  s_79_23,  s_79_24,  s_79_25;
wire   s_80_0,   s_80_1,   s_80_2,   s_80_3,   s_80_4,   s_80_5;
wire   s_80_6,   s_80_7,   s_80_8,   s_80_9,  s_80_10,  s_80_11;
wire  s_80_12,  s_80_13,  s_80_14,  s_80_15,  s_80_16,  s_80_17;
wire  s_80_18,  s_80_19,  s_80_20,  s_80_21,  s_80_22,  s_80_23;
wire  s_80_24,   s_81_0,   s_81_1,   s_81_2,   s_81_3,   s_81_4;
wire   s_81_5,   s_81_6,   s_81_7,   s_81_8,   s_81_9,  s_81_10;
wire  s_81_11,  s_81_12,  s_81_13,  s_81_14,  s_81_15,  s_81_16;
wire  s_81_17,  s_81_18,  s_81_19,  s_81_20,  s_81_21,  s_81_22;
wire  s_81_23,  s_81_24,   s_82_0,   s_82_1,   s_82_2,   s_82_3;
wire   s_82_4,   s_82_5,   s_82_6,   s_82_7,   s_82_8,   s_82_9;
wire  s_82_10,  s_82_11,  s_82_12,  s_82_13,  s_82_14,  s_82_15;
wire  s_82_16,  s_82_17,  s_82_18,  s_82_19,  s_82_20,  s_82_21;
wire  s_82_22,  s_82_23,   s_83_0,   s_83_1,   s_83_2,   s_83_3;
wire   s_83_4,   s_83_5,   s_83_6,   s_83_7,   s_83_8,   s_83_9;
wire  s_83_10,  s_83_11,  s_83_12,  s_83_13,  s_83_14,  s_83_15;
wire  s_83_16,  s_83_17,  s_83_18,  s_83_19,  s_83_20,  s_83_21;
wire  s_83_22,  s_83_23,   s_84_0,   s_84_1,   s_84_2,   s_84_3;
wire   s_84_4,   s_84_5,   s_84_6,   s_84_7,   s_84_8,   s_84_9;
wire  s_84_10,  s_84_11,  s_84_12,  s_84_13,  s_84_14,  s_84_15;
wire  s_84_16,  s_84_17,  s_84_18,  s_84_19,  s_84_20,  s_84_21;
wire  s_84_22,   s_85_0,   s_85_1,   s_85_2,   s_85_3,   s_85_4;
wire   s_85_5,   s_85_6,   s_85_7,   s_85_8,   s_85_9,  s_85_10;
wire  s_85_11,  s_85_12,  s_85_13,  s_85_14,  s_85_15,  s_85_16;
wire  s_85_17,  s_85_18,  s_85_19,  s_85_20,  s_85_21,  s_85_22;
wire   s_86_0,   s_86_1,   s_86_2,   s_86_3,   s_86_4,   s_86_5;
wire   s_86_6,   s_86_7,   s_86_8,   s_86_9,  s_86_10,  s_86_11;
wire  s_86_12,  s_86_13,  s_86_14,  s_86_15,  s_86_16,  s_86_17;
wire  s_86_18,  s_86_19,  s_86_20,  s_86_21,   s_87_0,   s_87_1;
wire   s_87_2,   s_87_3,   s_87_4,   s_87_5,   s_87_6,   s_87_7;
wire   s_87_8,   s_87_9,  s_87_10,  s_87_11,  s_87_12,  s_87_13;
wire  s_87_14,  s_87_15,  s_87_16,  s_87_17,  s_87_18,  s_87_19;
wire  s_87_20,  s_87_21,   s_88_0,   s_88_1,   s_88_2,   s_88_3;
wire   s_88_4,   s_88_5,   s_88_6,   s_88_7,   s_88_8,   s_88_9;
wire  s_88_10,  s_88_11,  s_88_12,  s_88_13,  s_88_14,  s_88_15;
wire  s_88_16,  s_88_17,  s_88_18,  s_88_19,  s_88_20,   s_89_0;
wire   s_89_1,   s_89_2,   s_89_3,   s_89_4,   s_89_5,   s_89_6;
wire   s_89_7,   s_89_8,   s_89_9,  s_89_10,  s_89_11,  s_89_12;
wire  s_89_13,  s_89_14,  s_89_15,  s_89_16,  s_89_17,  s_89_18;
wire  s_89_19,  s_89_20,   s_90_0,   s_90_1,   s_90_2,   s_90_3;
wire   s_90_4,   s_90_5,   s_90_6,   s_90_7,   s_90_8,   s_90_9;
wire  s_90_10,  s_90_11,  s_90_12,  s_90_13,  s_90_14,  s_90_15;
wire  s_90_16,  s_90_17,  s_90_18,  s_90_19,   s_91_0,   s_91_1;
wire   s_91_2,   s_91_3,   s_91_4,   s_91_5,   s_91_6,   s_91_7;
wire   s_91_8,   s_91_9,  s_91_10,  s_91_11,  s_91_12,  s_91_13;
wire  s_91_14,  s_91_15,  s_91_16,  s_91_17,  s_91_18,  s_91_19;
wire   s_92_0,   s_92_1,   s_92_2,   s_92_3,   s_92_4,   s_92_5;
wire   s_92_6,   s_92_7,   s_92_8,   s_92_9,  s_92_10,  s_92_11;
wire  s_92_12,  s_92_13,  s_92_14,  s_92_15,  s_92_16,  s_92_17;
wire  s_92_18,   s_93_0,   s_93_1,   s_93_2,   s_93_3,   s_93_4;
wire   s_93_5,   s_93_6,   s_93_7,   s_93_8,   s_93_9,  s_93_10;
wire  s_93_11,  s_93_12,  s_93_13,  s_93_14,  s_93_15,  s_93_16;
wire  s_93_17,  s_93_18,   s_94_0,   s_94_1,   s_94_2,   s_94_3;
wire   s_94_4,   s_94_5,   s_94_6,   s_94_7,   s_94_8,   s_94_9;
wire  s_94_10,  s_94_11,  s_94_12,  s_94_13,  s_94_14,  s_94_15;
wire  s_94_16,  s_94_17,   s_95_0,   s_95_1,   s_95_2,   s_95_3;
wire   s_95_4,   s_95_5,   s_95_6,   s_95_7,   s_95_8,   s_95_9;
wire  s_95_10,  s_95_11,  s_95_12,  s_95_13,  s_95_14,  s_95_15;
wire  s_95_16,  s_95_17,   s_96_0,   s_96_1,   s_96_2,   s_96_3;
wire   s_96_4,   s_96_5,   s_96_6,   s_96_7,   s_96_8,   s_96_9;
wire  s_96_10,  s_96_11,  s_96_12,  s_96_13,  s_96_14,  s_96_15;
wire  s_96_16,   s_97_0,   s_97_1,   s_97_2,   s_97_3,   s_97_4;
wire   s_97_5,   s_97_6,   s_97_7,   s_97_8,   s_97_9,  s_97_10;
wire  s_97_11,  s_97_12,  s_97_13,  s_97_14,  s_97_15,  s_97_16;
wire   s_98_0,   s_98_1,   s_98_2,   s_98_3,   s_98_4,   s_98_5;
wire   s_98_6,   s_98_7,   s_98_8,   s_98_9,  s_98_10,  s_98_11;
wire  s_98_12,  s_98_13,  s_98_14,  s_98_15,   s_99_0,   s_99_1;
wire   s_99_2,   s_99_3,   s_99_4,   s_99_5,   s_99_6,   s_99_7;
wire   s_99_8,   s_99_9,  s_99_10,  s_99_11,  s_99_12,  s_99_13;
wire  s_99_14,  s_99_15,  s_100_0,  s_100_1,  s_100_2,  s_100_3;
wire  s_100_4,  s_100_5,  s_100_6,  s_100_7,  s_100_8,  s_100_9;
wire s_100_10, s_100_11, s_100_12, s_100_13, s_100_14,  s_101_0;
wire  s_101_1,  s_101_2,  s_101_3,  s_101_4,  s_101_5,  s_101_6;
wire  s_101_7,  s_101_8,  s_101_9, s_101_10, s_101_11, s_101_12;
wire s_101_13, s_101_14,  s_102_0,  s_102_1,  s_102_2,  s_102_3;
wire  s_102_4,  s_102_5,  s_102_6,  s_102_7,  s_102_8,  s_102_9;
wire s_102_10, s_102_11, s_102_12, s_102_13,  s_103_0,  s_103_1;
wire  s_103_2,  s_103_3,  s_103_4,  s_103_5,  s_103_6,  s_103_7;
wire  s_103_8,  s_103_9, s_103_10, s_103_11, s_103_12, s_103_13;
wire  s_104_0,  s_104_1,  s_104_2,  s_104_3,  s_104_4,  s_104_5;
wire  s_104_6,  s_104_7,  s_104_8,  s_104_9, s_104_10, s_104_11;
wire s_104_12,  s_105_0,  s_105_1,  s_105_2,  s_105_3,  s_105_4;
wire  s_105_5,  s_105_6,  s_105_7,  s_105_8,  s_105_9, s_105_10;
wire s_105_11, s_105_12,  s_106_0,  s_106_1,  s_106_2,  s_106_3;
wire  s_106_4,  s_106_5,  s_106_6,  s_106_7,  s_106_8,  s_106_9;
wire s_106_10, s_106_11,  s_107_0,  s_107_1,  s_107_2,  s_107_3;
wire  s_107_4,  s_107_5,  s_107_6,  s_107_7,  s_107_8,  s_107_9;
wire s_107_10, s_107_11,  s_108_0,  s_108_1,  s_108_2,  s_108_3;
wire  s_108_4,  s_108_5,  s_108_6,  s_108_7,  s_108_8,  s_108_9;
wire s_108_10,  s_109_0,  s_109_1,  s_109_2,  s_109_3,  s_109_4;
wire  s_109_5,  s_109_6,  s_109_7,  s_109_8,  s_109_9, s_109_10;
wire  s_110_0,  s_110_1,  s_110_2,  s_110_3,  s_110_4,  s_110_5;
wire  s_110_6,  s_110_7,  s_110_8,  s_110_9,  s_111_0,  s_111_1;
wire  s_111_2,  s_111_3,  s_111_4,  s_111_5,  s_111_6,  s_111_7;
wire  s_111_8,  s_111_9,  s_112_0,  s_112_1,  s_112_2,  s_112_3;
wire  s_112_4,  s_112_5,  s_112_6,  s_112_7,  s_112_8,  s_113_0;
wire  s_113_1,  s_113_2,  s_113_3,  s_113_4,  s_113_5,  s_113_6;
wire  s_113_7,  s_113_8,  s_114_0,  s_114_1,  s_114_2,  s_114_3;
wire  s_114_4,  s_114_5,  s_114_6,  s_114_7,  s_115_0,  s_115_1;
wire  s_115_2,  s_115_3,  s_115_4,  s_115_5,  s_115_6,  s_115_7;
wire  s_116_0,  s_116_1,  s_116_2,  s_116_3,  s_116_4,  s_116_5;
wire  s_116_6,  s_117_0,  s_117_1,  s_117_2,  s_117_3,  s_117_4;
wire  s_117_5,  s_117_6,  s_118_0,  s_118_1,  s_118_2,  s_118_3;
wire  s_118_4,  s_118_5,  s_119_0,  s_119_1,  s_119_2,  s_119_3;
wire  s_119_4,  s_119_5,  s_120_0,  s_120_1,  s_120_2,  s_120_3;
wire  s_120_4,  s_121_0,  s_121_1,  s_121_2,  s_121_3,  s_121_4;
wire  s_122_0,  s_122_1,  s_122_2,  s_122_3,  s_123_0,  s_123_1;
wire  s_123_2,  s_123_3,  s_124_0,  s_124_1,  s_124_2,  s_125_0;
wire  s_125_1,  s_125_2,  s_126_0,  s_126_1,  s_127_0,  s_127_1;

assign {
 s_62_32,  s_60_31,  s_58_30,  s_56_29,  s_54_28,  s_52_27, 
 s_50_26,  s_48_25,  s_46_24,  s_44_23,  s_42_22,  s_40_21, 
 s_38_20,  s_36_19,  s_34_18,  s_32_17,  s_30_16,  s_28_15, 
 s_26_14,  s_24_13,  s_22_12,  s_20_11,  s_18_10,   s_16_9, 
  s_14_8,   s_12_7,   s_10_6,    s_8_5,    s_6_4,    s_4_3, 
   s_2_2,    s_0_1
} = carry;

assign {
  s_65_0,   s_64_0,   s_63_0,   s_62_0,   s_61_0,   s_60_0, 
  s_59_0,   s_58_0,   s_57_0,   s_56_0,   s_55_0,   s_54_0, 
  s_53_0,   s_52_0,   s_51_0,   s_50_0,   s_49_0,   s_48_0, 
  s_47_0,   s_46_0,   s_45_0,   s_44_0,   s_43_0,   s_42_0, 
  s_41_0,   s_40_0,   s_39_0,   s_38_0,   s_37_0,   s_36_0, 
  s_35_0,   s_34_0,   s_33_0,   s_32_0,   s_31_0,   s_30_0, 
  s_29_0,   s_28_0,   s_27_0,   s_26_0,   s_25_0,   s_24_0, 
  s_23_0,   s_22_0,   s_21_0,   s_20_0,   s_19_0,   s_18_0, 
  s_17_0,   s_16_0,   s_15_0,   s_14_0,   s_13_0,   s_12_0, 
  s_11_0,   s_10_0,    s_9_0,    s_8_0,    s_7_0,    s_6_0, 
   s_5_0,    s_4_0,    s_3_0,    s_2_0,    s_1_0,    s_0_0
} = partial_products[(width+2)*(0+1)-1:(width+2)*0];

assign {
  s_67_0,   s_66_0,   s_65_1,   s_64_1,   s_63_1,   s_62_1, 
  s_61_1,   s_60_1,   s_59_1,   s_58_1,   s_57_1,   s_56_1, 
  s_55_1,   s_54_1,   s_53_1,   s_52_1,   s_51_1,   s_50_1, 
  s_49_1,   s_48_1,   s_47_1,   s_46_1,   s_45_1,   s_44_1, 
  s_43_1,   s_42_1,   s_41_1,   s_40_1,   s_39_1,   s_38_1, 
  s_37_1,   s_36_1,   s_35_1,   s_34_1,   s_33_1,   s_32_1, 
  s_31_1,   s_30_1,   s_29_1,   s_28_1,   s_27_1,   s_26_1, 
  s_25_1,   s_24_1,   s_23_1,   s_22_1,   s_21_1,   s_20_1, 
  s_19_1,   s_18_1,   s_17_1,   s_16_1,   s_15_1,   s_14_1, 
  s_13_1,   s_12_1,   s_11_1,   s_10_1,    s_9_1,    s_8_1, 
   s_7_1,    s_6_1,    s_5_1,    s_4_1,    s_3_1,    s_2_1
} = partial_products[(width+2)*(1+1)-1:(width+2)*1];

assign {
  s_69_0,   s_68_0,   s_67_1,   s_66_1,   s_65_2,   s_64_2, 
  s_63_2,   s_62_2,   s_61_2,   s_60_2,   s_59_2,   s_58_2, 
  s_57_2,   s_56_2,   s_55_2,   s_54_2,   s_53_2,   s_52_2, 
  s_51_2,   s_50_2,   s_49_2,   s_48_2,   s_47_2,   s_46_2, 
  s_45_2,   s_44_2,   s_43_2,   s_42_2,   s_41_2,   s_40_2, 
  s_39_2,   s_38_2,   s_37_2,   s_36_2,   s_35_2,   s_34_2, 
  s_33_2,   s_32_2,   s_31_2,   s_30_2,   s_29_2,   s_28_2, 
  s_27_2,   s_26_2,   s_25_2,   s_24_2,   s_23_2,   s_22_2, 
  s_21_2,   s_20_2,   s_19_2,   s_18_2,   s_17_2,   s_16_2, 
  s_15_2,   s_14_2,   s_13_2,   s_12_2,   s_11_2,   s_10_2, 
   s_9_2,    s_8_2,    s_7_2,    s_6_2,    s_5_2,    s_4_2
} = partial_products[(width+2)*(2+1)-1:(width+2)*2];

assign {
  s_71_0,   s_70_0,   s_69_1,   s_68_1,   s_67_2,   s_66_2, 
  s_65_3,   s_64_3,   s_63_3,   s_62_3,   s_61_3,   s_60_3, 
  s_59_3,   s_58_3,   s_57_3,   s_56_3,   s_55_3,   s_54_3, 
  s_53_3,   s_52_3,   s_51_3,   s_50_3,   s_49_3,   s_48_3, 
  s_47_3,   s_46_3,   s_45_3,   s_44_3,   s_43_3,   s_42_3, 
  s_41_3,   s_40_3,   s_39_3,   s_38_3,   s_37_3,   s_36_3, 
  s_35_3,   s_34_3,   s_33_3,   s_32_3,   s_31_3,   s_30_3, 
  s_29_3,   s_28_3,   s_27_3,   s_26_3,   s_25_3,   s_24_3, 
  s_23_3,   s_22_3,   s_21_3,   s_20_3,   s_19_3,   s_18_3, 
  s_17_3,   s_16_3,   s_15_3,   s_14_3,   s_13_3,   s_12_3, 
  s_11_3,   s_10_3,    s_9_3,    s_8_3,    s_7_3,    s_6_3
} = partial_products[(width+2)*(3+1)-1:(width+2)*3];

assign {
  s_73_0,   s_72_0,   s_71_1,   s_70_1,   s_69_2,   s_68_2, 
  s_67_3,   s_66_3,   s_65_4,   s_64_4,   s_63_4,   s_62_4, 
  s_61_4,   s_60_4,   s_59_4,   s_58_4,   s_57_4,   s_56_4, 
  s_55_4,   s_54_4,   s_53_4,   s_52_4,   s_51_4,   s_50_4, 
  s_49_4,   s_48_4,   s_47_4,   s_46_4,   s_45_4,   s_44_4, 
  s_43_4,   s_42_4,   s_41_4,   s_40_4,   s_39_4,   s_38_4, 
  s_37_4,   s_36_4,   s_35_4,   s_34_4,   s_33_4,   s_32_4, 
  s_31_4,   s_30_4,   s_29_4,   s_28_4,   s_27_4,   s_26_4, 
  s_25_4,   s_24_4,   s_23_4,   s_22_4,   s_21_4,   s_20_4, 
  s_19_4,   s_18_4,   s_17_4,   s_16_4,   s_15_4,   s_14_4, 
  s_13_4,   s_12_4,   s_11_4,   s_10_4,    s_9_4,    s_8_4
} = partial_products[(width+2)*(4+1)-1:(width+2)*4];

assign {
  s_75_0,   s_74_0,   s_73_1,   s_72_1,   s_71_2,   s_70_2, 
  s_69_3,   s_68_3,   s_67_4,   s_66_4,   s_65_5,   s_64_5, 
  s_63_5,   s_62_5,   s_61_5,   s_60_5,   s_59_5,   s_58_5, 
  s_57_5,   s_56_5,   s_55_5,   s_54_5,   s_53_5,   s_52_5, 
  s_51_5,   s_50_5,   s_49_5,   s_48_5,   s_47_5,   s_46_5, 
  s_45_5,   s_44_5,   s_43_5,   s_42_5,   s_41_5,   s_40_5, 
  s_39_5,   s_38_5,   s_37_5,   s_36_5,   s_35_5,   s_34_5, 
  s_33_5,   s_32_5,   s_31_5,   s_30_5,   s_29_5,   s_28_5, 
  s_27_5,   s_26_5,   s_25_5,   s_24_5,   s_23_5,   s_22_5, 
  s_21_5,   s_20_5,   s_19_5,   s_18_5,   s_17_5,   s_16_5, 
  s_15_5,   s_14_5,   s_13_5,   s_12_5,   s_11_5,   s_10_5
} = partial_products[(width+2)*(5+1)-1:(width+2)*5];

assign {
  s_77_0,   s_76_0,   s_75_1,   s_74_1,   s_73_2,   s_72_2, 
  s_71_3,   s_70_3,   s_69_4,   s_68_4,   s_67_5,   s_66_5, 
  s_65_6,   s_64_6,   s_63_6,   s_62_6,   s_61_6,   s_60_6, 
  s_59_6,   s_58_6,   s_57_6,   s_56_6,   s_55_6,   s_54_6, 
  s_53_6,   s_52_6,   s_51_6,   s_50_6,   s_49_6,   s_48_6, 
  s_47_6,   s_46_6,   s_45_6,   s_44_6,   s_43_6,   s_42_6, 
  s_41_6,   s_40_6,   s_39_6,   s_38_6,   s_37_6,   s_36_6, 
  s_35_6,   s_34_6,   s_33_6,   s_32_6,   s_31_6,   s_30_6, 
  s_29_6,   s_28_6,   s_27_6,   s_26_6,   s_25_6,   s_24_6, 
  s_23_6,   s_22_6,   s_21_6,   s_20_6,   s_19_6,   s_18_6, 
  s_17_6,   s_16_6,   s_15_6,   s_14_6,   s_13_6,   s_12_6
} = partial_products[(width+2)*(6+1)-1:(width+2)*6];

assign {
  s_79_0,   s_78_0,   s_77_1,   s_76_1,   s_75_2,   s_74_2, 
  s_73_3,   s_72_3,   s_71_4,   s_70_4,   s_69_5,   s_68_5, 
  s_67_6,   s_66_6,   s_65_7,   s_64_7,   s_63_7,   s_62_7, 
  s_61_7,   s_60_7,   s_59_7,   s_58_7,   s_57_7,   s_56_7, 
  s_55_7,   s_54_7,   s_53_7,   s_52_7,   s_51_7,   s_50_7, 
  s_49_7,   s_48_7,   s_47_7,   s_46_7,   s_45_7,   s_44_7, 
  s_43_7,   s_42_7,   s_41_7,   s_40_7,   s_39_7,   s_38_7, 
  s_37_7,   s_36_7,   s_35_7,   s_34_7,   s_33_7,   s_32_7, 
  s_31_7,   s_30_7,   s_29_7,   s_28_7,   s_27_7,   s_26_7, 
  s_25_7,   s_24_7,   s_23_7,   s_22_7,   s_21_7,   s_20_7, 
  s_19_7,   s_18_7,   s_17_7,   s_16_7,   s_15_7,   s_14_7
} = partial_products[(width+2)*(7+1)-1:(width+2)*7];

assign {
  s_81_0,   s_80_0,   s_79_1,   s_78_1,   s_77_2,   s_76_2, 
  s_75_3,   s_74_3,   s_73_4,   s_72_4,   s_71_5,   s_70_5, 
  s_69_6,   s_68_6,   s_67_7,   s_66_7,   s_65_8,   s_64_8, 
  s_63_8,   s_62_8,   s_61_8,   s_60_8,   s_59_8,   s_58_8, 
  s_57_8,   s_56_8,   s_55_8,   s_54_8,   s_53_8,   s_52_8, 
  s_51_8,   s_50_8,   s_49_8,   s_48_8,   s_47_8,   s_46_8, 
  s_45_8,   s_44_8,   s_43_8,   s_42_8,   s_41_8,   s_40_8, 
  s_39_8,   s_38_8,   s_37_8,   s_36_8,   s_35_8,   s_34_8, 
  s_33_8,   s_32_8,   s_31_8,   s_30_8,   s_29_8,   s_28_8, 
  s_27_8,   s_26_8,   s_25_8,   s_24_8,   s_23_8,   s_22_8, 
  s_21_8,   s_20_8,   s_19_8,   s_18_8,   s_17_8,   s_16_8
} = partial_products[(width+2)*(8+1)-1:(width+2)*8];

assign {
  s_83_0,   s_82_0,   s_81_1,   s_80_1,   s_79_2,   s_78_2, 
  s_77_3,   s_76_3,   s_75_4,   s_74_4,   s_73_5,   s_72_5, 
  s_71_6,   s_70_6,   s_69_7,   s_68_7,   s_67_8,   s_66_8, 
  s_65_9,   s_64_9,   s_63_9,   s_62_9,   s_61_9,   s_60_9, 
  s_59_9,   s_58_9,   s_57_9,   s_56_9,   s_55_9,   s_54_9, 
  s_53_9,   s_52_9,   s_51_9,   s_50_9,   s_49_9,   s_48_9, 
  s_47_9,   s_46_9,   s_45_9,   s_44_9,   s_43_9,   s_42_9, 
  s_41_9,   s_40_9,   s_39_9,   s_38_9,   s_37_9,   s_36_9, 
  s_35_9,   s_34_9,   s_33_9,   s_32_9,   s_31_9,   s_30_9, 
  s_29_9,   s_28_9,   s_27_9,   s_26_9,   s_25_9,   s_24_9, 
  s_23_9,   s_22_9,   s_21_9,   s_20_9,   s_19_9,   s_18_9
} = partial_products[(width+2)*(9+1)-1:(width+2)*9];

assign {
  s_85_0,   s_84_0,   s_83_1,   s_82_1,   s_81_2,   s_80_2, 
  s_79_3,   s_78_3,   s_77_4,   s_76_4,   s_75_5,   s_74_5, 
  s_73_6,   s_72_6,   s_71_7,   s_70_7,   s_69_8,   s_68_8, 
  s_67_9,   s_66_9,  s_65_10,  s_64_10,  s_63_10,  s_62_10, 
 s_61_10,  s_60_10,  s_59_10,  s_58_10,  s_57_10,  s_56_10, 
 s_55_10,  s_54_10,  s_53_10,  s_52_10,  s_51_10,  s_50_10, 
 s_49_10,  s_48_10,  s_47_10,  s_46_10,  s_45_10,  s_44_10, 
 s_43_10,  s_42_10,  s_41_10,  s_40_10,  s_39_10,  s_38_10, 
 s_37_10,  s_36_10,  s_35_10,  s_34_10,  s_33_10,  s_32_10, 
 s_31_10,  s_30_10,  s_29_10,  s_28_10,  s_27_10,  s_26_10, 
 s_25_10,  s_24_10,  s_23_10,  s_22_10,  s_21_10,  s_20_10
} = partial_products[(width+2)*(10+1)-1:(width+2)*10];

assign {
  s_87_0,   s_86_0,   s_85_1,   s_84_1,   s_83_2,   s_82_2, 
  s_81_3,   s_80_3,   s_79_4,   s_78_4,   s_77_5,   s_76_5, 
  s_75_6,   s_74_6,   s_73_7,   s_72_7,   s_71_8,   s_70_8, 
  s_69_9,   s_68_9,  s_67_10,  s_66_10,  s_65_11,  s_64_11, 
 s_63_11,  s_62_11,  s_61_11,  s_60_11,  s_59_11,  s_58_11, 
 s_57_11,  s_56_11,  s_55_11,  s_54_11,  s_53_11,  s_52_11, 
 s_51_11,  s_50_11,  s_49_11,  s_48_11,  s_47_11,  s_46_11, 
 s_45_11,  s_44_11,  s_43_11,  s_42_11,  s_41_11,  s_40_11, 
 s_39_11,  s_38_11,  s_37_11,  s_36_11,  s_35_11,  s_34_11, 
 s_33_11,  s_32_11,  s_31_11,  s_30_11,  s_29_11,  s_28_11, 
 s_27_11,  s_26_11,  s_25_11,  s_24_11,  s_23_11,  s_22_11
} = partial_products[(width+2)*(11+1)-1:(width+2)*11];

assign {
  s_89_0,   s_88_0,   s_87_1,   s_86_1,   s_85_2,   s_84_2, 
  s_83_3,   s_82_3,   s_81_4,   s_80_4,   s_79_5,   s_78_5, 
  s_77_6,   s_76_6,   s_75_7,   s_74_7,   s_73_8,   s_72_8, 
  s_71_9,   s_70_9,  s_69_10,  s_68_10,  s_67_11,  s_66_11, 
 s_65_12,  s_64_12,  s_63_12,  s_62_12,  s_61_12,  s_60_12, 
 s_59_12,  s_58_12,  s_57_12,  s_56_12,  s_55_12,  s_54_12, 
 s_53_12,  s_52_12,  s_51_12,  s_50_12,  s_49_12,  s_48_12, 
 s_47_12,  s_46_12,  s_45_12,  s_44_12,  s_43_12,  s_42_12, 
 s_41_12,  s_40_12,  s_39_12,  s_38_12,  s_37_12,  s_36_12, 
 s_35_12,  s_34_12,  s_33_12,  s_32_12,  s_31_12,  s_30_12, 
 s_29_12,  s_28_12,  s_27_12,  s_26_12,  s_25_12,  s_24_12
} = partial_products[(width+2)*(12+1)-1:(width+2)*12];

assign {
  s_91_0,   s_90_0,   s_89_1,   s_88_1,   s_87_2,   s_86_2, 
  s_85_3,   s_84_3,   s_83_4,   s_82_4,   s_81_5,   s_80_5, 
  s_79_6,   s_78_6,   s_77_7,   s_76_7,   s_75_8,   s_74_8, 
  s_73_9,   s_72_9,  s_71_10,  s_70_10,  s_69_11,  s_68_11, 
 s_67_12,  s_66_12,  s_65_13,  s_64_13,  s_63_13,  s_62_13, 
 s_61_13,  s_60_13,  s_59_13,  s_58_13,  s_57_13,  s_56_13, 
 s_55_13,  s_54_13,  s_53_13,  s_52_13,  s_51_13,  s_50_13, 
 s_49_13,  s_48_13,  s_47_13,  s_46_13,  s_45_13,  s_44_13, 
 s_43_13,  s_42_13,  s_41_13,  s_40_13,  s_39_13,  s_38_13, 
 s_37_13,  s_36_13,  s_35_13,  s_34_13,  s_33_13,  s_32_13, 
 s_31_13,  s_30_13,  s_29_13,  s_28_13,  s_27_13,  s_26_13
} = partial_products[(width+2)*(13+1)-1:(width+2)*13];

assign {
  s_93_0,   s_92_0,   s_91_1,   s_90_1,   s_89_2,   s_88_2, 
  s_87_3,   s_86_3,   s_85_4,   s_84_4,   s_83_5,   s_82_5, 
  s_81_6,   s_80_6,   s_79_7,   s_78_7,   s_77_8,   s_76_8, 
  s_75_9,   s_74_9,  s_73_10,  s_72_10,  s_71_11,  s_70_11, 
 s_69_12,  s_68_12,  s_67_13,  s_66_13,  s_65_14,  s_64_14, 
 s_63_14,  s_62_14,  s_61_14,  s_60_14,  s_59_14,  s_58_14, 
 s_57_14,  s_56_14,  s_55_14,  s_54_14,  s_53_14,  s_52_14, 
 s_51_14,  s_50_14,  s_49_14,  s_48_14,  s_47_14,  s_46_14, 
 s_45_14,  s_44_14,  s_43_14,  s_42_14,  s_41_14,  s_40_14, 
 s_39_14,  s_38_14,  s_37_14,  s_36_14,  s_35_14,  s_34_14, 
 s_33_14,  s_32_14,  s_31_14,  s_30_14,  s_29_14,  s_28_14
} = partial_products[(width+2)*(14+1)-1:(width+2)*14];

assign {
  s_95_0,   s_94_0,   s_93_1,   s_92_1,   s_91_2,   s_90_2, 
  s_89_3,   s_88_3,   s_87_4,   s_86_4,   s_85_5,   s_84_5, 
  s_83_6,   s_82_6,   s_81_7,   s_80_7,   s_79_8,   s_78_8, 
  s_77_9,   s_76_9,  s_75_10,  s_74_10,  s_73_11,  s_72_11, 
 s_71_12,  s_70_12,  s_69_13,  s_68_13,  s_67_14,  s_66_14, 
 s_65_15,  s_64_15,  s_63_15,  s_62_15,  s_61_15,  s_60_15, 
 s_59_15,  s_58_15,  s_57_15,  s_56_15,  s_55_15,  s_54_15, 
 s_53_15,  s_52_15,  s_51_15,  s_50_15,  s_49_15,  s_48_15, 
 s_47_15,  s_46_15,  s_45_15,  s_44_15,  s_43_15,  s_42_15, 
 s_41_15,  s_40_15,  s_39_15,  s_38_15,  s_37_15,  s_36_15, 
 s_35_15,  s_34_15,  s_33_15,  s_32_15,  s_31_15,  s_30_15
} = partial_products[(width+2)*(15+1)-1:(width+2)*15];

assign {
  s_97_0,   s_96_0,   s_95_1,   s_94_1,   s_93_2,   s_92_2, 
  s_91_3,   s_90_3,   s_89_4,   s_88_4,   s_87_5,   s_86_5, 
  s_85_6,   s_84_6,   s_83_7,   s_82_7,   s_81_8,   s_80_8, 
  s_79_9,   s_78_9,  s_77_10,  s_76_10,  s_75_11,  s_74_11, 
 s_73_12,  s_72_12,  s_71_13,  s_70_13,  s_69_14,  s_68_14, 
 s_67_15,  s_66_15,  s_65_16,  s_64_16,  s_63_16,  s_62_16, 
 s_61_16,  s_60_16,  s_59_16,  s_58_16,  s_57_16,  s_56_16, 
 s_55_16,  s_54_16,  s_53_16,  s_52_16,  s_51_16,  s_50_16, 
 s_49_16,  s_48_16,  s_47_16,  s_46_16,  s_45_16,  s_44_16, 
 s_43_16,  s_42_16,  s_41_16,  s_40_16,  s_39_16,  s_38_16, 
 s_37_16,  s_36_16,  s_35_16,  s_34_16,  s_33_16,  s_32_16
} = partial_products[(width+2)*(16+1)-1:(width+2)*16];

assign {
  s_99_0,   s_98_0,   s_97_1,   s_96_1,   s_95_2,   s_94_2, 
  s_93_3,   s_92_3,   s_91_4,   s_90_4,   s_89_5,   s_88_5, 
  s_87_6,   s_86_6,   s_85_7,   s_84_7,   s_83_8,   s_82_8, 
  s_81_9,   s_80_9,  s_79_10,  s_78_10,  s_77_11,  s_76_11, 
 s_75_12,  s_74_12,  s_73_13,  s_72_13,  s_71_14,  s_70_14, 
 s_69_15,  s_68_15,  s_67_16,  s_66_16,  s_65_17,  s_64_17, 
 s_63_17,  s_62_17,  s_61_17,  s_60_17,  s_59_17,  s_58_17, 
 s_57_17,  s_56_17,  s_55_17,  s_54_17,  s_53_17,  s_52_17, 
 s_51_17,  s_50_17,  s_49_17,  s_48_17,  s_47_17,  s_46_17, 
 s_45_17,  s_44_17,  s_43_17,  s_42_17,  s_41_17,  s_40_17, 
 s_39_17,  s_38_17,  s_37_17,  s_36_17,  s_35_17,  s_34_17
} = partial_products[(width+2)*(17+1)-1:(width+2)*17];

assign {
 s_101_0,  s_100_0,   s_99_1,   s_98_1,   s_97_2,   s_96_2, 
  s_95_3,   s_94_3,   s_93_4,   s_92_4,   s_91_5,   s_90_5, 
  s_89_6,   s_88_6,   s_87_7,   s_86_7,   s_85_8,   s_84_8, 
  s_83_9,   s_82_9,  s_81_10,  s_80_10,  s_79_11,  s_78_11, 
 s_77_12,  s_76_12,  s_75_13,  s_74_13,  s_73_14,  s_72_14, 
 s_71_15,  s_70_15,  s_69_16,  s_68_16,  s_67_17,  s_66_17, 
 s_65_18,  s_64_18,  s_63_18,  s_62_18,  s_61_18,  s_60_18, 
 s_59_18,  s_58_18,  s_57_18,  s_56_18,  s_55_18,  s_54_18, 
 s_53_18,  s_52_18,  s_51_18,  s_50_18,  s_49_18,  s_48_18, 
 s_47_18,  s_46_18,  s_45_18,  s_44_18,  s_43_18,  s_42_18, 
 s_41_18,  s_40_18,  s_39_18,  s_38_18,  s_37_18,  s_36_18
} = partial_products[(width+2)*(18+1)-1:(width+2)*18];

assign {
 s_103_0,  s_102_0,  s_101_1,  s_100_1,   s_99_2,   s_98_2, 
  s_97_3,   s_96_3,   s_95_4,   s_94_4,   s_93_5,   s_92_5, 
  s_91_6,   s_90_6,   s_89_7,   s_88_7,   s_87_8,   s_86_8, 
  s_85_9,   s_84_9,  s_83_10,  s_82_10,  s_81_11,  s_80_11, 
 s_79_12,  s_78_12,  s_77_13,  s_76_13,  s_75_14,  s_74_14, 
 s_73_15,  s_72_15,  s_71_16,  s_70_16,  s_69_17,  s_68_17, 
 s_67_18,  s_66_18,  s_65_19,  s_64_19,  s_63_19,  s_62_19, 
 s_61_19,  s_60_19,  s_59_19,  s_58_19,  s_57_19,  s_56_19, 
 s_55_19,  s_54_19,  s_53_19,  s_52_19,  s_51_19,  s_50_19, 
 s_49_19,  s_48_19,  s_47_19,  s_46_19,  s_45_19,  s_44_19, 
 s_43_19,  s_42_19,  s_41_19,  s_40_19,  s_39_19,  s_38_19
} = partial_products[(width+2)*(19+1)-1:(width+2)*19];

assign {
 s_105_0,  s_104_0,  s_103_1,  s_102_1,  s_101_2,  s_100_2, 
  s_99_3,   s_98_3,   s_97_4,   s_96_4,   s_95_5,   s_94_5, 
  s_93_6,   s_92_6,   s_91_7,   s_90_7,   s_89_8,   s_88_8, 
  s_87_9,   s_86_9,  s_85_10,  s_84_10,  s_83_11,  s_82_11, 
 s_81_12,  s_80_12,  s_79_13,  s_78_13,  s_77_14,  s_76_14, 
 s_75_15,  s_74_15,  s_73_16,  s_72_16,  s_71_17,  s_70_17, 
 s_69_18,  s_68_18,  s_67_19,  s_66_19,  s_65_20,  s_64_20, 
 s_63_20,  s_62_20,  s_61_20,  s_60_20,  s_59_20,  s_58_20, 
 s_57_20,  s_56_20,  s_55_20,  s_54_20,  s_53_20,  s_52_20, 
 s_51_20,  s_50_20,  s_49_20,  s_48_20,  s_47_20,  s_46_20, 
 s_45_20,  s_44_20,  s_43_20,  s_42_20,  s_41_20,  s_40_20
} = partial_products[(width+2)*(20+1)-1:(width+2)*20];

assign {
 s_107_0,  s_106_0,  s_105_1,  s_104_1,  s_103_2,  s_102_2, 
 s_101_3,  s_100_3,   s_99_4,   s_98_4,   s_97_5,   s_96_5, 
  s_95_6,   s_94_6,   s_93_7,   s_92_7,   s_91_8,   s_90_8, 
  s_89_9,   s_88_9,  s_87_10,  s_86_10,  s_85_11,  s_84_11, 
 s_83_12,  s_82_12,  s_81_13,  s_80_13,  s_79_14,  s_78_14, 
 s_77_15,  s_76_15,  s_75_16,  s_74_16,  s_73_17,  s_72_17, 
 s_71_18,  s_70_18,  s_69_19,  s_68_19,  s_67_20,  s_66_20, 
 s_65_21,  s_64_21,  s_63_21,  s_62_21,  s_61_21,  s_60_21, 
 s_59_21,  s_58_21,  s_57_21,  s_56_21,  s_55_21,  s_54_21, 
 s_53_21,  s_52_21,  s_51_21,  s_50_21,  s_49_21,  s_48_21, 
 s_47_21,  s_46_21,  s_45_21,  s_44_21,  s_43_21,  s_42_21
} = partial_products[(width+2)*(21+1)-1:(width+2)*21];

assign {
 s_109_0,  s_108_0,  s_107_1,  s_106_1,  s_105_2,  s_104_2, 
 s_103_3,  s_102_3,  s_101_4,  s_100_4,   s_99_5,   s_98_5, 
  s_97_6,   s_96_6,   s_95_7,   s_94_7,   s_93_8,   s_92_8, 
  s_91_9,   s_90_9,  s_89_10,  s_88_10,  s_87_11,  s_86_11, 
 s_85_12,  s_84_12,  s_83_13,  s_82_13,  s_81_14,  s_80_14, 
 s_79_15,  s_78_15,  s_77_16,  s_76_16,  s_75_17,  s_74_17, 
 s_73_18,  s_72_18,  s_71_19,  s_70_19,  s_69_20,  s_68_20, 
 s_67_21,  s_66_21,  s_65_22,  s_64_22,  s_63_22,  s_62_22, 
 s_61_22,  s_60_22,  s_59_22,  s_58_22,  s_57_22,  s_56_22, 
 s_55_22,  s_54_22,  s_53_22,  s_52_22,  s_51_22,  s_50_22, 
 s_49_22,  s_48_22,  s_47_22,  s_46_22,  s_45_22,  s_44_22
} = partial_products[(width+2)*(22+1)-1:(width+2)*22];

assign {
 s_111_0,  s_110_0,  s_109_1,  s_108_1,  s_107_2,  s_106_2, 
 s_105_3,  s_104_3,  s_103_4,  s_102_4,  s_101_5,  s_100_5, 
  s_99_6,   s_98_6,   s_97_7,   s_96_7,   s_95_8,   s_94_8, 
  s_93_9,   s_92_9,  s_91_10,  s_90_10,  s_89_11,  s_88_11, 
 s_87_12,  s_86_12,  s_85_13,  s_84_13,  s_83_14,  s_82_14, 
 s_81_15,  s_80_15,  s_79_16,  s_78_16,  s_77_17,  s_76_17, 
 s_75_18,  s_74_18,  s_73_19,  s_72_19,  s_71_20,  s_70_20, 
 s_69_21,  s_68_21,  s_67_22,  s_66_22,  s_65_23,  s_64_23, 
 s_63_23,  s_62_23,  s_61_23,  s_60_23,  s_59_23,  s_58_23, 
 s_57_23,  s_56_23,  s_55_23,  s_54_23,  s_53_23,  s_52_23, 
 s_51_23,  s_50_23,  s_49_23,  s_48_23,  s_47_23,  s_46_23
} = partial_products[(width+2)*(23+1)-1:(width+2)*23];

assign {
 s_113_0,  s_112_0,  s_111_1,  s_110_1,  s_109_2,  s_108_2, 
 s_107_3,  s_106_3,  s_105_4,  s_104_4,  s_103_5,  s_102_5, 
 s_101_6,  s_100_6,   s_99_7,   s_98_7,   s_97_8,   s_96_8, 
  s_95_9,   s_94_9,  s_93_10,  s_92_10,  s_91_11,  s_90_11, 
 s_89_12,  s_88_12,  s_87_13,  s_86_13,  s_85_14,  s_84_14, 
 s_83_15,  s_82_15,  s_81_16,  s_80_16,  s_79_17,  s_78_17, 
 s_77_18,  s_76_18,  s_75_19,  s_74_19,  s_73_20,  s_72_20, 
 s_71_21,  s_70_21,  s_69_22,  s_68_22,  s_67_23,  s_66_23, 
 s_65_24,  s_64_24,  s_63_24,  s_62_24,  s_61_24,  s_60_24, 
 s_59_24,  s_58_24,  s_57_24,  s_56_24,  s_55_24,  s_54_24, 
 s_53_24,  s_52_24,  s_51_24,  s_50_24,  s_49_24,  s_48_24
} = partial_products[(width+2)*(24+1)-1:(width+2)*24];

assign {
 s_115_0,  s_114_0,  s_113_1,  s_112_1,  s_111_2,  s_110_2, 
 s_109_3,  s_108_3,  s_107_4,  s_106_4,  s_105_5,  s_104_5, 
 s_103_6,  s_102_6,  s_101_7,  s_100_7,   s_99_8,   s_98_8, 
  s_97_9,   s_96_9,  s_95_10,  s_94_10,  s_93_11,  s_92_11, 
 s_91_12,  s_90_12,  s_89_13,  s_88_13,  s_87_14,  s_86_14, 
 s_85_15,  s_84_15,  s_83_16,  s_82_16,  s_81_17,  s_80_17, 
 s_79_18,  s_78_18,  s_77_19,  s_76_19,  s_75_20,  s_74_20, 
 s_73_21,  s_72_21,  s_71_22,  s_70_22,  s_69_23,  s_68_23, 
 s_67_24,  s_66_24,  s_65_25,  s_64_25,  s_63_25,  s_62_25, 
 s_61_25,  s_60_25,  s_59_25,  s_58_25,  s_57_25,  s_56_25, 
 s_55_25,  s_54_25,  s_53_25,  s_52_25,  s_51_25,  s_50_25
} = partial_products[(width+2)*(25+1)-1:(width+2)*25];

assign {
 s_117_0,  s_116_0,  s_115_1,  s_114_1,  s_113_2,  s_112_2, 
 s_111_3,  s_110_3,  s_109_4,  s_108_4,  s_107_5,  s_106_5, 
 s_105_6,  s_104_6,  s_103_7,  s_102_7,  s_101_8,  s_100_8, 
  s_99_9,   s_98_9,  s_97_10,  s_96_10,  s_95_11,  s_94_11, 
 s_93_12,  s_92_12,  s_91_13,  s_90_13,  s_89_14,  s_88_14, 
 s_87_15,  s_86_15,  s_85_16,  s_84_16,  s_83_17,  s_82_17, 
 s_81_18,  s_80_18,  s_79_19,  s_78_19,  s_77_20,  s_76_20, 
 s_75_21,  s_74_21,  s_73_22,  s_72_22,  s_71_23,  s_70_23, 
 s_69_24,  s_68_24,  s_67_25,  s_66_25,  s_65_26,  s_64_26, 
 s_63_26,  s_62_26,  s_61_26,  s_60_26,  s_59_26,  s_58_26, 
 s_57_26,  s_56_26,  s_55_26,  s_54_26,  s_53_26,  s_52_26
} = partial_products[(width+2)*(26+1)-1:(width+2)*26];

assign {
 s_119_0,  s_118_0,  s_117_1,  s_116_1,  s_115_2,  s_114_2, 
 s_113_3,  s_112_3,  s_111_4,  s_110_4,  s_109_5,  s_108_5, 
 s_107_6,  s_106_6,  s_105_7,  s_104_7,  s_103_8,  s_102_8, 
 s_101_9,  s_100_9,  s_99_10,  s_98_10,  s_97_11,  s_96_11, 
 s_95_12,  s_94_12,  s_93_13,  s_92_13,  s_91_14,  s_90_14, 
 s_89_15,  s_88_15,  s_87_16,  s_86_16,  s_85_17,  s_84_17, 
 s_83_18,  s_82_18,  s_81_19,  s_80_19,  s_79_20,  s_78_20, 
 s_77_21,  s_76_21,  s_75_22,  s_74_22,  s_73_23,  s_72_23, 
 s_71_24,  s_70_24,  s_69_25,  s_68_25,  s_67_26,  s_66_26, 
 s_65_27,  s_64_27,  s_63_27,  s_62_27,  s_61_27,  s_60_27, 
 s_59_27,  s_58_27,  s_57_27,  s_56_27,  s_55_27,  s_54_27
} = partial_products[(width+2)*(27+1)-1:(width+2)*27];

assign {
 s_121_0,  s_120_0,  s_119_1,  s_118_1,  s_117_2,  s_116_2, 
 s_115_3,  s_114_3,  s_113_4,  s_112_4,  s_111_5,  s_110_5, 
 s_109_6,  s_108_6,  s_107_7,  s_106_7,  s_105_8,  s_104_8, 
 s_103_9,  s_102_9, s_101_10, s_100_10,  s_99_11,  s_98_11, 
 s_97_12,  s_96_12,  s_95_13,  s_94_13,  s_93_14,  s_92_14, 
 s_91_15,  s_90_15,  s_89_16,  s_88_16,  s_87_17,  s_86_17, 
 s_85_18,  s_84_18,  s_83_19,  s_82_19,  s_81_20,  s_80_20, 
 s_79_21,  s_78_21,  s_77_22,  s_76_22,  s_75_23,  s_74_23, 
 s_73_24,  s_72_24,  s_71_25,  s_70_25,  s_69_26,  s_68_26, 
 s_67_27,  s_66_27,  s_65_28,  s_64_28,  s_63_28,  s_62_28, 
 s_61_28,  s_60_28,  s_59_28,  s_58_28,  s_57_28,  s_56_28
} = partial_products[(width+2)*(28+1)-1:(width+2)*28];

assign {
 s_123_0,  s_122_0,  s_121_1,  s_120_1,  s_119_2,  s_118_2, 
 s_117_3,  s_116_3,  s_115_4,  s_114_4,  s_113_5,  s_112_5, 
 s_111_6,  s_110_6,  s_109_7,  s_108_7,  s_107_8,  s_106_8, 
 s_105_9,  s_104_9, s_103_10, s_102_10, s_101_11, s_100_11, 
 s_99_12,  s_98_12,  s_97_13,  s_96_13,  s_95_14,  s_94_14, 
 s_93_15,  s_92_15,  s_91_16,  s_90_16,  s_89_17,  s_88_17, 
 s_87_18,  s_86_18,  s_85_19,  s_84_19,  s_83_20,  s_82_20, 
 s_81_21,  s_80_21,  s_79_22,  s_78_22,  s_77_23,  s_76_23, 
 s_75_24,  s_74_24,  s_73_25,  s_72_25,  s_71_26,  s_70_26, 
 s_69_27,  s_68_27,  s_67_28,  s_66_28,  s_65_29,  s_64_29, 
 s_63_29,  s_62_29,  s_61_29,  s_60_29,  s_59_29,  s_58_29
} = partial_products[(width+2)*(29+1)-1:(width+2)*29];

assign {
 s_125_0,  s_124_0,  s_123_1,  s_122_1,  s_121_2,  s_120_2, 
 s_119_3,  s_118_3,  s_117_4,  s_116_4,  s_115_5,  s_114_5, 
 s_113_6,  s_112_6,  s_111_7,  s_110_7,  s_109_8,  s_108_8, 
 s_107_9,  s_106_9, s_105_10, s_104_10, s_103_11, s_102_11, 
s_101_12, s_100_12,  s_99_13,  s_98_13,  s_97_14,  s_96_14, 
 s_95_15,  s_94_15,  s_93_16,  s_92_16,  s_91_17,  s_90_17, 
 s_89_18,  s_88_18,  s_87_19,  s_86_19,  s_85_20,  s_84_20, 
 s_83_21,  s_82_21,  s_81_22,  s_80_22,  s_79_23,  s_78_23, 
 s_77_24,  s_76_24,  s_75_25,  s_74_25,  s_73_26,  s_72_26, 
 s_71_27,  s_70_27,  s_69_28,  s_68_28,  s_67_29,  s_66_29, 
 s_65_30,  s_64_30,  s_63_30,  s_62_30,  s_61_30,  s_60_30
} = partial_products[(width+2)*(30+1)-1:(width+2)*30];

assign {
 s_127_0,  s_126_0,  s_125_1,  s_124_1,  s_123_2,  s_122_2, 
 s_121_3,  s_120_3,  s_119_4,  s_118_4,  s_117_5,  s_116_5, 
 s_115_6,  s_114_6,  s_113_7,  s_112_7,  s_111_8,  s_110_8, 
 s_109_9,  s_108_9, s_107_10, s_106_10, s_105_11, s_104_11, 
s_103_12, s_102_12, s_101_13, s_100_13,  s_99_14,  s_98_14, 
 s_97_15,  s_96_15,  s_95_16,  s_94_16,  s_93_17,  s_92_17, 
 s_91_18,  s_90_18,  s_89_19,  s_88_19,  s_87_20,  s_86_20, 
 s_85_21,  s_84_21,  s_83_22,  s_82_22,  s_81_23,  s_80_23, 
 s_79_24,  s_78_24,  s_77_25,  s_76_25,  s_75_26,  s_74_26, 
 s_73_27,  s_72_27,  s_71_28,  s_70_28,  s_69_29,  s_68_29, 
 s_67_30,  s_66_30,  s_65_31,  s_64_31,  s_63_31,  s_62_31
} = partial_products[(width+2)*(31+1)-1:(width+2)*31];

assign {
 s_127_1,  s_126_1,  s_125_2,  s_124_2,  s_123_3,  s_122_3, 
 s_121_4,  s_120_4,  s_119_5,  s_118_5,  s_117_6,  s_116_6, 
 s_115_7,  s_114_7,  s_113_8,  s_112_8,  s_111_9,  s_110_9, 
s_109_10, s_108_10, s_107_11, s_106_11, s_105_12, s_104_12, 
s_103_13, s_102_13, s_101_14, s_100_14,  s_99_15,  s_98_15, 
 s_97_16,  s_96_16,  s_95_17,  s_94_17,  s_93_18,  s_92_18, 
 s_91_19,  s_90_19,  s_89_20,  s_88_20,  s_87_21,  s_86_21, 
 s_85_22,  s_84_22,  s_83_23,  s_82_23,  s_81_24,  s_80_24, 
 s_79_25,  s_78_25,  s_77_26,  s_76_26,  s_75_27,  s_74_27, 
 s_73_28,  s_72_28,  s_71_29,  s_70_29,  s_69_30,  s_68_30, 
 s_67_31,  s_66_31,  s_65_32,  s_64_32
} = partial_products[(width+2)*(width/2+1)-1:(width+2)*width/2+2];

/* u0_1 Output nets */
wire t_0,      t_1;
/* u1_2 Output nets */
wire t_2,      t_3;
/* u0_3 Output nets */
wire t_4,      t_5;
/* u2_4 Output nets */
wire t_6,      t_7,      t_8;
/* u1_5 Output nets */
wire t_9,     t_10;
/* u2_6 Output nets */
wire t_11,     t_12,     t_13;
/* u2_7 Output nets */
wire t_14,     t_15,     t_16;
/* u2_8 Output nets */
wire t_17,     t_18,     t_19;
/* u0_9 Output nets */
wire t_20,     t_21;
/* u2_10 Output nets */
wire t_22,     t_23,     t_24;
/* u0_11 Output nets */
wire t_25,     t_26;
/* u2_12 Output nets */
wire t_27,     t_28,     t_29;
/* u1_13 Output nets */
wire t_30,     t_31;
/* u2_14 Output nets */
wire t_32,     t_33,     t_34;
/* u1_15 Output nets */
wire t_35,     t_36;
/* u2_16 Output nets */
wire t_37,     t_38,     t_39;
/* u2_17 Output nets */
wire t_40,     t_41,     t_42;
/* u2_18 Output nets */
wire t_43,     t_44,     t_45;
/* u1_19 Output nets */
wire t_46,     t_47;
/* u2_20 Output nets */
wire t_48,     t_49,     t_50;
/* u2_21 Output nets */
wire t_51,     t_52,     t_53;
/* u2_22 Output nets */
wire t_54,     t_55,     t_56;
/* u2_23 Output nets */
wire t_57,     t_58,     t_59;
/* u2_24 Output nets */
wire t_60,     t_61,     t_62;
/* u2_25 Output nets */
wire t_63,     t_64,     t_65;
/* u0_26 Output nets */
wire t_66,     t_67;
/* u2_27 Output nets */
wire t_68,     t_69,     t_70;
/* u2_28 Output nets */
wire t_71,     t_72,     t_73;
/* u0_29 Output nets */
wire t_74,     t_75;
/* u2_30 Output nets */
wire t_76,     t_77,     t_78;
/* u2_31 Output nets */
wire t_79,     t_80,     t_81;
/* u1_32 Output nets */
wire t_82,     t_83;
/* u2_33 Output nets */
wire t_84,     t_85,     t_86;
/* u2_34 Output nets */
wire t_87,     t_88,     t_89;
/* u1_35 Output nets */
wire t_90,     t_91;
/* u2_36 Output nets */
wire t_92,     t_93,     t_94;
/* u2_37 Output nets */
wire t_95,     t_96,     t_97;
/* u2_38 Output nets */
wire t_98,     t_99,    t_100;
/* u2_39 Output nets */
wire t_101,    t_102,    t_103;
/* u2_40 Output nets */
wire t_104,    t_105,    t_106;
/* u1_41 Output nets */
wire t_107,    t_108;
/* u2_42 Output nets */
wire t_109,    t_110,    t_111;
/* u2_43 Output nets */
wire t_112,    t_113,    t_114;
/* u2_44 Output nets */
wire t_115,    t_116,    t_117;
/* u2_45 Output nets */
wire t_118,    t_119,    t_120;
/* u2_46 Output nets */
wire t_121,    t_122,    t_123;
/* u2_47 Output nets */
wire t_124,    t_125,    t_126;
/* u2_48 Output nets */
wire t_127,    t_128,    t_129;
/* u2_49 Output nets */
wire t_130,    t_131,    t_132;
/* u2_50 Output nets */
wire t_133,    t_134,    t_135;
/* u0_51 Output nets */
wire t_136,    t_137;
/* u2_52 Output nets */
wire t_138,    t_139,    t_140;
/* u2_53 Output nets */
wire t_141,    t_142,    t_143;
/* u2_54 Output nets */
wire t_144,    t_145,    t_146;
/* u0_55 Output nets */
wire t_147,    t_148;
/* u2_56 Output nets */
wire t_149,    t_150,    t_151;
/* u2_57 Output nets */
wire t_152,    t_153,    t_154;
/* u2_58 Output nets */
wire t_155,    t_156,    t_157;
/* u1_59 Output nets */
wire t_158,    t_159;
/* u2_60 Output nets */
wire t_160,    t_161,    t_162;
/* u2_61 Output nets */
wire t_163,    t_164,    t_165;
/* u2_62 Output nets */
wire t_166,    t_167,    t_168;
/* u1_63 Output nets */
wire t_169,    t_170;
/* u2_64 Output nets */
wire t_171,    t_172,    t_173;
/* u2_65 Output nets */
wire t_174,    t_175,    t_176;
/* u2_66 Output nets */
wire t_177,    t_178,    t_179;
/* u2_67 Output nets */
wire t_180,    t_181,    t_182;
/* u2_68 Output nets */
wire t_183,    t_184,    t_185;
/* u2_69 Output nets */
wire t_186,    t_187,    t_188;
/* u2_70 Output nets */
wire t_189,    t_190,    t_191;
/* u1_71 Output nets */
wire t_192,    t_193;
/* u2_72 Output nets */
wire t_194,    t_195,    t_196;
/* u2_73 Output nets */
wire t_197,    t_198,    t_199;
/* u2_74 Output nets */
wire t_200,    t_201,    t_202;
/* u2_75 Output nets */
wire t_203,    t_204,    t_205;
/* u2_76 Output nets */
wire t_206,    t_207,    t_208;
/* u2_77 Output nets */
wire t_209,    t_210,    t_211;
/* u2_78 Output nets */
wire t_212,    t_213,    t_214;
/* u2_79 Output nets */
wire t_215,    t_216,    t_217;
/* u2_80 Output nets */
wire t_218,    t_219,    t_220;
/* u2_81 Output nets */
wire t_221,    t_222,    t_223;
/* u2_82 Output nets */
wire t_224,    t_225,    t_226;
/* u2_83 Output nets */
wire t_227,    t_228,    t_229;
/* u0_84 Output nets */
wire t_230,    t_231;
/* u2_85 Output nets */
wire t_232,    t_233,    t_234;
/* u2_86 Output nets */
wire t_235,    t_236,    t_237;
/* u2_87 Output nets */
wire t_238,    t_239,    t_240;
/* u2_88 Output nets */
wire t_241,    t_242,    t_243;
/* u0_89 Output nets */
wire t_244,    t_245;
/* u2_90 Output nets */
wire t_246,    t_247,    t_248;
/* u2_91 Output nets */
wire t_249,    t_250,    t_251;
/* u2_92 Output nets */
wire t_252,    t_253,    t_254;
/* u2_93 Output nets */
wire t_255,    t_256,    t_257;
/* u1_94 Output nets */
wire t_258,    t_259;
/* u2_95 Output nets */
wire t_260,    t_261,    t_262;
/* u2_96 Output nets */
wire t_263,    t_264,    t_265;
/* u2_97 Output nets */
wire t_266,    t_267,    t_268;
/* u2_98 Output nets */
wire t_269,    t_270,    t_271;
/* u1_99 Output nets */
wire t_272,    t_273;
/* u2_100 Output nets */
wire t_274,    t_275,    t_276;
/* u2_101 Output nets */
wire t_277,    t_278,    t_279;
/* u2_102 Output nets */
wire t_280,    t_281,    t_282;
/* u2_103 Output nets */
wire t_283,    t_284,    t_285;
/* u2_104 Output nets */
wire t_286,    t_287,    t_288;
/* u2_105 Output nets */
wire t_289,    t_290,    t_291;
/* u2_106 Output nets */
wire t_292,    t_293,    t_294;
/* u2_107 Output nets */
wire t_295,    t_296,    t_297;
/* u2_108 Output nets */
wire t_298,    t_299,    t_300;
/* u1_109 Output nets */
wire t_301,    t_302;
/* u2_110 Output nets */
wire t_303,    t_304,    t_305;
/* u2_111 Output nets */
wire t_306,    t_307,    t_308;
/* u2_112 Output nets */
wire t_309,    t_310,    t_311;
/* u2_113 Output nets */
wire t_312,    t_313,    t_314;
/* u2_114 Output nets */
wire t_315,    t_316,    t_317;
/* u2_115 Output nets */
wire t_318,    t_319,    t_320;
/* u2_116 Output nets */
wire t_321,    t_322,    t_323;
/* u2_117 Output nets */
wire t_324,    t_325,    t_326;
/* u2_118 Output nets */
wire t_327,    t_328,    t_329;
/* u2_119 Output nets */
wire t_330,    t_331,    t_332;
/* u2_120 Output nets */
wire t_333,    t_334,    t_335;
/* u2_121 Output nets */
wire t_336,    t_337,    t_338;
/* u2_122 Output nets */
wire t_339,    t_340,    t_341;
/* u2_123 Output nets */
wire t_342,    t_343,    t_344;
/* u2_124 Output nets */
wire t_345,    t_346,    t_347;
/* u0_125 Output nets */
wire t_348,    t_349;
/* u2_126 Output nets */
wire t_350,    t_351,    t_352;
/* u2_127 Output nets */
wire t_353,    t_354,    t_355;
/* u2_128 Output nets */
wire t_356,    t_357,    t_358;
/* u2_129 Output nets */
wire t_359,    t_360,    t_361;
/* u2_130 Output nets */
wire t_362,    t_363,    t_364;
/* u0_131 Output nets */
wire t_365,    t_366;
/* u2_132 Output nets */
wire t_367,    t_368,    t_369;
/* u2_133 Output nets */
wire t_370,    t_371,    t_372;
/* u2_134 Output nets */
wire t_373,    t_374,    t_375;
/* u2_135 Output nets */
wire t_376,    t_377,    t_378;
/* u2_136 Output nets */
wire t_379,    t_380,    t_381;
/* u1_137 Output nets */
wire t_382,    t_383;
/* u2_138 Output nets */
wire t_384,    t_385,    t_386;
/* u2_139 Output nets */
wire t_387,    t_388,    t_389;
/* u2_140 Output nets */
wire t_390,    t_391,    t_392;
/* u2_141 Output nets */
wire t_393,    t_394,    t_395;
/* u2_142 Output nets */
wire t_396,    t_397,    t_398;
/* u1_143 Output nets */
wire t_399,    t_400;
/* u2_144 Output nets */
wire t_401,    t_402,    t_403;
/* u2_145 Output nets */
wire t_404,    t_405,    t_406;
/* u2_146 Output nets */
wire t_407,    t_408,    t_409;
/* u2_147 Output nets */
wire t_410,    t_411,    t_412;
/* u2_148 Output nets */
wire t_413,    t_414,    t_415;
/* u2_149 Output nets */
wire t_416,    t_417,    t_418;
/* u2_150 Output nets */
wire t_419,    t_420,    t_421;
/* u2_151 Output nets */
wire t_422,    t_423,    t_424;
/* u2_152 Output nets */
wire t_425,    t_426,    t_427;
/* u2_153 Output nets */
wire t_428,    t_429,    t_430;
/* u2_154 Output nets */
wire t_431,    t_432,    t_433;
/* u1_155 Output nets */
wire t_434,    t_435;
/* u2_156 Output nets */
wire t_436,    t_437,    t_438;
/* u2_157 Output nets */
wire t_439,    t_440,    t_441;
/* u2_158 Output nets */
wire t_442,    t_443,    t_444;
/* u2_159 Output nets */
wire t_445,    t_446,    t_447;
/* u2_160 Output nets */
wire t_448,    t_449,    t_450;
/* u2_161 Output nets */
wire t_451,    t_452,    t_453;
/* u2_162 Output nets */
wire t_454,    t_455,    t_456;
/* u2_163 Output nets */
wire t_457,    t_458,    t_459;
/* u2_164 Output nets */
wire t_460,    t_461,    t_462;
/* u2_165 Output nets */
wire t_463,    t_464,    t_465;
/* u2_166 Output nets */
wire t_466,    t_467,    t_468;
/* u2_167 Output nets */
wire t_469,    t_470,    t_471;
/* u2_168 Output nets */
wire t_472,    t_473,    t_474;
/* u2_169 Output nets */
wire t_475,    t_476,    t_477;
/* u2_170 Output nets */
wire t_478,    t_479,    t_480;
/* u2_171 Output nets */
wire t_481,    t_482,    t_483;
/* u2_172 Output nets */
wire t_484,    t_485,    t_486;
/* u2_173 Output nets */
wire t_487,    t_488,    t_489;
/* u0_174 Output nets */
wire t_490,    t_491;
/* u2_175 Output nets */
wire t_492,    t_493,    t_494;
/* u2_176 Output nets */
wire t_495,    t_496,    t_497;
/* u2_177 Output nets */
wire t_498,    t_499,    t_500;
/* u2_178 Output nets */
wire t_501,    t_502,    t_503;
/* u2_179 Output nets */
wire t_504,    t_505,    t_506;
/* u2_180 Output nets */
wire t_507,    t_508,    t_509;
/* u0_181 Output nets */
wire t_510,    t_511;
/* u2_182 Output nets */
wire t_512,    t_513,    t_514;
/* u2_183 Output nets */
wire t_515,    t_516,    t_517;
/* u2_184 Output nets */
wire t_518,    t_519,    t_520;
/* u2_185 Output nets */
wire t_521,    t_522,    t_523;
/* u2_186 Output nets */
wire t_524,    t_525,    t_526;
/* u2_187 Output nets */
wire t_527,    t_528,    t_529;
/* u1_188 Output nets */
wire t_530,    t_531;
/* u2_189 Output nets */
wire t_532,    t_533,    t_534;
/* u2_190 Output nets */
wire t_535,    t_536,    t_537;
/* u2_191 Output nets */
wire t_538,    t_539,    t_540;
/* u2_192 Output nets */
wire t_541,    t_542,    t_543;
/* u2_193 Output nets */
wire t_544,    t_545,    t_546;
/* u2_194 Output nets */
wire t_547,    t_548,    t_549;
/* u1_195 Output nets */
wire t_550,    t_551;
/* u2_196 Output nets */
wire t_552,    t_553,    t_554;
/* u2_197 Output nets */
wire t_555,    t_556,    t_557;
/* u2_198 Output nets */
wire t_558,    t_559,    t_560;
/* u2_199 Output nets */
wire t_561,    t_562,    t_563;
/* u2_200 Output nets */
wire t_564,    t_565,    t_566;
/* u2_201 Output nets */
wire t_567,    t_568,    t_569;
/* u2_202 Output nets */
wire t_570,    t_571,    t_572;
/* u2_203 Output nets */
wire t_573,    t_574,    t_575;
/* u2_204 Output nets */
wire t_576,    t_577,    t_578;
/* u2_205 Output nets */
wire t_579,    t_580,    t_581;
/* u2_206 Output nets */
wire t_582,    t_583,    t_584;
/* u2_207 Output nets */
wire t_585,    t_586,    t_587;
/* u2_208 Output nets */
wire t_588,    t_589,    t_590;
/* u1_209 Output nets */
wire t_591,    t_592;
/* u2_210 Output nets */
wire t_593,    t_594,    t_595;
/* u2_211 Output nets */
wire t_596,    t_597,    t_598;
/* u2_212 Output nets */
wire t_599,    t_600,    t_601;
/* u2_213 Output nets */
wire t_602,    t_603,    t_604;
/* u2_214 Output nets */
wire t_605,    t_606,    t_607;
/* u2_215 Output nets */
wire t_608,    t_609,    t_610;
/* u2_216 Output nets */
wire t_611,    t_612,    t_613;
/* u2_217 Output nets */
wire t_614,    t_615,    t_616;
/* u2_218 Output nets */
wire t_617,    t_618,    t_619;
/* u2_219 Output nets */
wire t_620,    t_621,    t_622;
/* u2_220 Output nets */
wire t_623,    t_624,    t_625;
/* u2_221 Output nets */
wire t_626,    t_627,    t_628;
/* u2_222 Output nets */
wire t_629,    t_630,    t_631;
/* u2_223 Output nets */
wire t_632,    t_633,    t_634;
/* u2_224 Output nets */
wire t_635,    t_636,    t_637;
/* u2_225 Output nets */
wire t_638,    t_639,    t_640;
/* u2_226 Output nets */
wire t_641,    t_642,    t_643;
/* u2_227 Output nets */
wire t_644,    t_645,    t_646;
/* u2_228 Output nets */
wire t_647,    t_648,    t_649;
/* u2_229 Output nets */
wire t_650,    t_651,    t_652;
/* u2_230 Output nets */
wire t_653,    t_654,    t_655;
/* u0_231 Output nets */
wire t_656,    t_657;
/* u2_232 Output nets */
wire t_658,    t_659,    t_660;
/* u2_233 Output nets */
wire t_661,    t_662,    t_663;
/* u2_234 Output nets */
wire t_664,    t_665,    t_666;
/* u2_235 Output nets */
wire t_667,    t_668,    t_669;
/* u2_236 Output nets */
wire t_670,    t_671,    t_672;
/* u2_237 Output nets */
wire t_673,    t_674,    t_675;
/* u2_238 Output nets */
wire t_676,    t_677,    t_678;
/* u0_239 Output nets */
wire t_679,    t_680;
/* u2_240 Output nets */
wire t_681,    t_682,    t_683;
/* u2_241 Output nets */
wire t_684,    t_685,    t_686;
/* u2_242 Output nets */
wire t_687,    t_688,    t_689;
/* u2_243 Output nets */
wire t_690,    t_691,    t_692;
/* u2_244 Output nets */
wire t_693,    t_694,    t_695;
/* u2_245 Output nets */
wire t_696,    t_697,    t_698;
/* u2_246 Output nets */
wire t_699,    t_700,    t_701;
/* u1_247 Output nets */
wire t_702,    t_703;
/* u2_248 Output nets */
wire t_704,    t_705,    t_706;
/* u2_249 Output nets */
wire t_707,    t_708,    t_709;
/* u2_250 Output nets */
wire t_710,    t_711,    t_712;
/* u2_251 Output nets */
wire t_713,    t_714,    t_715;
/* u2_252 Output nets */
wire t_716,    t_717,    t_718;
/* u2_253 Output nets */
wire t_719,    t_720,    t_721;
/* u2_254 Output nets */
wire t_722,    t_723,    t_724;
/* u1_255 Output nets */
wire t_725,    t_726;
/* u2_256 Output nets */
wire t_727,    t_728,    t_729;
/* u2_257 Output nets */
wire t_730,    t_731,    t_732;
/* u2_258 Output nets */
wire t_733,    t_734,    t_735;
/* u2_259 Output nets */
wire t_736,    t_737,    t_738;
/* u2_260 Output nets */
wire t_739,    t_740,    t_741;
/* u2_261 Output nets */
wire t_742,    t_743,    t_744;
/* u2_262 Output nets */
wire t_745,    t_746,    t_747;
/* u2_263 Output nets */
wire t_748,    t_749,    t_750;
/* u2_264 Output nets */
wire t_751,    t_752,    t_753;
/* u2_265 Output nets */
wire t_754,    t_755,    t_756;
/* u2_266 Output nets */
wire t_757,    t_758,    t_759;
/* u2_267 Output nets */
wire t_760,    t_761,    t_762;
/* u2_268 Output nets */
wire t_763,    t_764,    t_765;
/* u2_269 Output nets */
wire t_766,    t_767,    t_768;
/* u2_270 Output nets */
wire t_769,    t_770,    t_771;
/* u1_271 Output nets */
wire t_772,    t_773;
/* u2_272 Output nets */
wire t_774,    t_775,    t_776;
/* u2_273 Output nets */
wire t_777,    t_778,    t_779;
/* u2_274 Output nets */
wire t_780,    t_781,    t_782;
/* u2_275 Output nets */
wire t_783,    t_784,    t_785;
/* u2_276 Output nets */
wire t_786,    t_787,    t_788;
/* u2_277 Output nets */
wire t_789,    t_790,    t_791;
/* u2_278 Output nets */
wire t_792,    t_793,    t_794;
/* u2_279 Output nets */
wire t_795,    t_796,    t_797;
/* u2_280 Output nets */
wire t_798,    t_799,    t_800;
/* u2_281 Output nets */
wire t_801,    t_802,    t_803;
/* u2_282 Output nets */
wire t_804,    t_805,    t_806;
/* u2_283 Output nets */
wire t_807,    t_808,    t_809;
/* u2_284 Output nets */
wire t_810,    t_811,    t_812;
/* u2_285 Output nets */
wire t_813,    t_814,    t_815;
/* u2_286 Output nets */
wire t_816,    t_817,    t_818;
/* u2_287 Output nets */
wire t_819,    t_820,    t_821;
/* u2_288 Output nets */
wire t_822,    t_823,    t_824;
/* u2_289 Output nets */
wire t_825,    t_826,    t_827;
/* u2_290 Output nets */
wire t_828,    t_829,    t_830;
/* u2_291 Output nets */
wire t_831,    t_832,    t_833;
/* u2_292 Output nets */
wire t_834,    t_835,    t_836;
/* u2_293 Output nets */
wire t_837,    t_838,    t_839;
/* u2_294 Output nets */
wire t_840,    t_841,    t_842;
/* u2_295 Output nets */
wire t_843,    t_844,    t_845;
/* u2_296 Output nets */
wire t_846,    t_847,    t_848;
/* u2_297 Output nets */
wire t_849,    t_850,    t_851;
/* u2_298 Output nets */
wire t_852,    t_853,    t_854;
/* u2_299 Output nets */
wire t_855,    t_856,    t_857;
/* u2_300 Output nets */
wire t_858,    t_859,    t_860;
/* u2_301 Output nets */
wire t_861,    t_862,    t_863;
/* u2_302 Output nets */
wire t_864,    t_865,    t_866;
/* u2_303 Output nets */
wire t_867,    t_868,    t_869;
/* u2_304 Output nets */
wire t_870,    t_871,    t_872;
/* u2_305 Output nets */
wire t_873,    t_874,    t_875;
/* u2_306 Output nets */
wire t_876,    t_877,    t_878;
/* u2_307 Output nets */
wire t_879,    t_880,    t_881;
/* u2_308 Output nets */
wire t_882,    t_883,    t_884;
/* u2_309 Output nets */
wire t_885,    t_886,    t_887;
/* u2_310 Output nets */
wire t_888,    t_889,    t_890;
/* u2_311 Output nets */
wire t_891,    t_892,    t_893;
/* u2_312 Output nets */
wire t_894,    t_895,    t_896;
/* u2_313 Output nets */
wire t_897,    t_898,    t_899;
/* u2_314 Output nets */
wire t_900,    t_901,    t_902;
/* u2_315 Output nets */
wire t_903,    t_904,    t_905;
/* u2_316 Output nets */
wire t_906,    t_907,    t_908;
/* u2_317 Output nets */
wire t_909,    t_910,    t_911;
/* u2_318 Output nets */
wire t_912,    t_913,    t_914;
/* u2_319 Output nets */
wire t_915,    t_916,    t_917;
/* u2_320 Output nets */
wire t_918,    t_919,    t_920;
/* u2_321 Output nets */
wire t_921,    t_922,    t_923;
/* u2_322 Output nets */
wire t_924,    t_925,    t_926;
/* u2_323 Output nets */
wire t_927,    t_928,    t_929;
/* u2_324 Output nets */
wire t_930,    t_931,    t_932;
/* u2_325 Output nets */
wire t_933,    t_934,    t_935;
/* u2_326 Output nets */
wire t_936,    t_937,    t_938;
/* u1_327 Output nets */
wire t_939,    t_940;
/* u2_328 Output nets */
wire t_941,    t_942,    t_943;
/* u2_329 Output nets */
wire t_944,    t_945,    t_946;
/* u2_330 Output nets */
wire t_947,    t_948,    t_949;
/* u2_331 Output nets */
wire t_950,    t_951,    t_952;
/* u2_332 Output nets */
wire t_953,    t_954,    t_955;
/* u2_333 Output nets */
wire t_956,    t_957,    t_958;
/* u2_334 Output nets */
wire t_959,    t_960,    t_961;
/* u1_335 Output nets */
wire t_962,    t_963;
/* u2_336 Output nets */
wire t_964,    t_965,    t_966;
/* u2_337 Output nets */
wire t_967,    t_968,    t_969;
/* u2_338 Output nets */
wire t_970,    t_971,    t_972;
/* u2_339 Output nets */
wire t_973,    t_974,    t_975;
/* u2_340 Output nets */
wire t_976,    t_977,    t_978;
/* u2_341 Output nets */
wire t_979,    t_980,    t_981;
/* u2_342 Output nets */
wire t_982,    t_983,    t_984;
/* u1_343 Output nets */
wire t_985,    t_986;
/* u2_344 Output nets */
wire t_987,    t_988,    t_989;
/* u2_345 Output nets */
wire t_990,    t_991,    t_992;
/* u2_346 Output nets */
wire t_993,    t_994,    t_995;
/* u2_347 Output nets */
wire t_996,    t_997,    t_998;
/* u2_348 Output nets */
wire t_999,   t_1000,   t_1001;
/* u2_349 Output nets */
wire t_1002,   t_1003,   t_1004;
/* u2_350 Output nets */
wire t_1005,   t_1006,   t_1007;
/* u1_351 Output nets */
wire t_1008,   t_1009;
/* u2_352 Output nets */
wire t_1010,   t_1011,   t_1012;
/* u2_353 Output nets */
wire t_1013,   t_1014,   t_1015;
/* u2_354 Output nets */
wire t_1016,   t_1017,   t_1018;
/* u2_355 Output nets */
wire t_1019,   t_1020,   t_1021;
/* u2_356 Output nets */
wire t_1022,   t_1023,   t_1024;
/* u2_357 Output nets */
wire t_1025,   t_1026,   t_1027;
/* u2_358 Output nets */
wire t_1028,   t_1029,   t_1030;
/* u0_359 Output nets */
wire t_1031,   t_1032;
/* u2_360 Output nets */
wire t_1033,   t_1034,   t_1035;
/* u2_361 Output nets */
wire t_1036,   t_1037,   t_1038;
/* u2_362 Output nets */
wire t_1039,   t_1040,   t_1041;
/* u2_363 Output nets */
wire t_1042,   t_1043,   t_1044;
/* u2_364 Output nets */
wire t_1045,   t_1046,   t_1047;
/* u2_365 Output nets */
wire t_1048,   t_1049,   t_1050;
/* u2_366 Output nets */
wire t_1051,   t_1052,   t_1053;
/* u0_367 Output nets */
wire t_1054,   t_1055;
/* u2_368 Output nets */
wire t_1056,   t_1057,   t_1058;
/* u2_369 Output nets */
wire t_1059,   t_1060,   t_1061;
/* u2_370 Output nets */
wire t_1062,   t_1063,   t_1064;
/* u2_371 Output nets */
wire t_1065,   t_1066,   t_1067;
/* u2_372 Output nets */
wire t_1068,   t_1069,   t_1070;
/* u2_373 Output nets */
wire t_1071,   t_1072,   t_1073;
/* u2_374 Output nets */
wire t_1074,   t_1075,   t_1076;
/* u2_375 Output nets */
wire t_1077,   t_1078,   t_1079;
/* u2_376 Output nets */
wire t_1080,   t_1081,   t_1082;
/* u2_377 Output nets */
wire t_1083,   t_1084,   t_1085;
/* u2_378 Output nets */
wire t_1086,   t_1087,   t_1088;
/* u2_379 Output nets */
wire t_1089,   t_1090,   t_1091;
/* u2_380 Output nets */
wire t_1092,   t_1093,   t_1094;
/* u2_381 Output nets */
wire t_1095,   t_1096,   t_1097;
/* u2_382 Output nets */
wire t_1098,   t_1099,   t_1100;
/* u2_383 Output nets */
wire t_1101,   t_1102,   t_1103;
/* u2_384 Output nets */
wire t_1104,   t_1105,   t_1106;
/* u2_385 Output nets */
wire t_1107,   t_1108,   t_1109;
/* u2_386 Output nets */
wire t_1110,   t_1111,   t_1112;
/* u2_387 Output nets */
wire t_1113,   t_1114,   t_1115;
/* u1_388 Output nets */
wire t_1116,   t_1117;
/* u2_389 Output nets */
wire t_1118,   t_1119,   t_1120;
/* u2_390 Output nets */
wire t_1121,   t_1122,   t_1123;
/* u2_391 Output nets */
wire t_1124,   t_1125,   t_1126;
/* u2_392 Output nets */
wire t_1127,   t_1128,   t_1129;
/* u2_393 Output nets */
wire t_1130,   t_1131,   t_1132;
/* u2_394 Output nets */
wire t_1133,   t_1134,   t_1135;
/* u1_395 Output nets */
wire t_1136,   t_1137;
/* u2_396 Output nets */
wire t_1138,   t_1139,   t_1140;
/* u2_397 Output nets */
wire t_1141,   t_1142,   t_1143;
/* u2_398 Output nets */
wire t_1144,   t_1145,   t_1146;
/* u2_399 Output nets */
wire t_1147,   t_1148,   t_1149;
/* u2_400 Output nets */
wire t_1150,   t_1151,   t_1152;
/* u2_401 Output nets */
wire t_1153,   t_1154,   t_1155;
/* u1_402 Output nets */
wire t_1156,   t_1157;
/* u2_403 Output nets */
wire t_1158,   t_1159,   t_1160;
/* u2_404 Output nets */
wire t_1161,   t_1162,   t_1163;
/* u2_405 Output nets */
wire t_1164,   t_1165,   t_1166;
/* u2_406 Output nets */
wire t_1167,   t_1168,   t_1169;
/* u2_407 Output nets */
wire t_1170,   t_1171,   t_1172;
/* u2_408 Output nets */
wire t_1173,   t_1174,   t_1175;
/* u1_409 Output nets */
wire t_1176,   t_1177;
/* u2_410 Output nets */
wire t_1178,   t_1179,   t_1180;
/* u2_411 Output nets */
wire t_1181,   t_1182,   t_1183;
/* u2_412 Output nets */
wire t_1184,   t_1185,   t_1186;
/* u2_413 Output nets */
wire t_1187,   t_1188,   t_1189;
/* u2_414 Output nets */
wire t_1190,   t_1191,   t_1192;
/* u2_415 Output nets */
wire t_1193,   t_1194,   t_1195;
/* u0_416 Output nets */
wire t_1196,   t_1197;
/* u2_417 Output nets */
wire t_1198,   t_1199,   t_1200;
/* u2_418 Output nets */
wire t_1201,   t_1202,   t_1203;
/* u2_419 Output nets */
wire t_1204,   t_1205,   t_1206;
/* u2_420 Output nets */
wire t_1207,   t_1208,   t_1209;
/* u2_421 Output nets */
wire t_1210,   t_1211,   t_1212;
/* u2_422 Output nets */
wire t_1213,   t_1214,   t_1215;
/* u0_423 Output nets */
wire t_1216,   t_1217;
/* u2_424 Output nets */
wire t_1218,   t_1219,   t_1220;
/* u2_425 Output nets */
wire t_1221,   t_1222,   t_1223;
/* u2_426 Output nets */
wire t_1224,   t_1225,   t_1226;
/* u2_427 Output nets */
wire t_1227,   t_1228,   t_1229;
/* u2_428 Output nets */
wire t_1230,   t_1231,   t_1232;
/* u2_429 Output nets */
wire t_1233,   t_1234,   t_1235;
/* u2_430 Output nets */
wire t_1236,   t_1237,   t_1238;
/* u2_431 Output nets */
wire t_1239,   t_1240,   t_1241;
/* u2_432 Output nets */
wire t_1242,   t_1243,   t_1244;
/* u2_433 Output nets */
wire t_1245,   t_1246,   t_1247;
/* u2_434 Output nets */
wire t_1248,   t_1249,   t_1250;
/* u2_435 Output nets */
wire t_1251,   t_1252,   t_1253;
/* u2_436 Output nets */
wire t_1254,   t_1255,   t_1256;
/* u2_437 Output nets */
wire t_1257,   t_1258,   t_1259;
/* u2_438 Output nets */
wire t_1260,   t_1261,   t_1262;
/* u2_439 Output nets */
wire t_1263,   t_1264,   t_1265;
/* u2_440 Output nets */
wire t_1266,   t_1267,   t_1268;
/* u1_441 Output nets */
wire t_1269,   t_1270;
/* u2_442 Output nets */
wire t_1271,   t_1272,   t_1273;
/* u2_443 Output nets */
wire t_1274,   t_1275,   t_1276;
/* u2_444 Output nets */
wire t_1277,   t_1278,   t_1279;
/* u2_445 Output nets */
wire t_1280,   t_1281,   t_1282;
/* u2_446 Output nets */
wire t_1283,   t_1284,   t_1285;
/* u1_447 Output nets */
wire t_1286,   t_1287;
/* u2_448 Output nets */
wire t_1288,   t_1289,   t_1290;
/* u2_449 Output nets */
wire t_1291,   t_1292,   t_1293;
/* u2_450 Output nets */
wire t_1294,   t_1295,   t_1296;
/* u2_451 Output nets */
wire t_1297,   t_1298,   t_1299;
/* u2_452 Output nets */
wire t_1300,   t_1301,   t_1302;
/* u1_453 Output nets */
wire t_1303,   t_1304;
/* u2_454 Output nets */
wire t_1305,   t_1306,   t_1307;
/* u2_455 Output nets */
wire t_1308,   t_1309,   t_1310;
/* u2_456 Output nets */
wire t_1311,   t_1312,   t_1313;
/* u2_457 Output nets */
wire t_1314,   t_1315,   t_1316;
/* u2_458 Output nets */
wire t_1317,   t_1318,   t_1319;
/* u1_459 Output nets */
wire t_1320,   t_1321;
/* u2_460 Output nets */
wire t_1322,   t_1323,   t_1324;
/* u2_461 Output nets */
wire t_1325,   t_1326,   t_1327;
/* u2_462 Output nets */
wire t_1328,   t_1329,   t_1330;
/* u2_463 Output nets */
wire t_1331,   t_1332,   t_1333;
/* u2_464 Output nets */
wire t_1334,   t_1335,   t_1336;
/* u0_465 Output nets */
wire t_1337,   t_1338;
/* u2_466 Output nets */
wire t_1339,   t_1340,   t_1341;
/* u2_467 Output nets */
wire t_1342,   t_1343,   t_1344;
/* u2_468 Output nets */
wire t_1345,   t_1346,   t_1347;
/* u2_469 Output nets */
wire t_1348,   t_1349,   t_1350;
/* u2_470 Output nets */
wire t_1351,   t_1352,   t_1353;
/* u0_471 Output nets */
wire t_1354,   t_1355;
/* u2_472 Output nets */
wire t_1356,   t_1357,   t_1358;
/* u2_473 Output nets */
wire t_1359,   t_1360,   t_1361;
/* u2_474 Output nets */
wire t_1362,   t_1363,   t_1364;
/* u2_475 Output nets */
wire t_1365,   t_1366,   t_1367;
/* u2_476 Output nets */
wire t_1368,   t_1369,   t_1370;
/* u2_477 Output nets */
wire t_1371,   t_1372,   t_1373;
/* u2_478 Output nets */
wire t_1374,   t_1375,   t_1376;
/* u2_479 Output nets */
wire t_1377,   t_1378,   t_1379;
/* u2_480 Output nets */
wire t_1380,   t_1381,   t_1382;
/* u2_481 Output nets */
wire t_1383,   t_1384,   t_1385;
/* u2_482 Output nets */
wire t_1386,   t_1387,   t_1388;
/* u2_483 Output nets */
wire t_1389,   t_1390,   t_1391;
/* u2_484 Output nets */
wire t_1392,   t_1393,   t_1394;
/* u2_485 Output nets */
wire t_1395,   t_1396,   t_1397;
/* u1_486 Output nets */
wire t_1398,   t_1399;
/* u2_487 Output nets */
wire t_1400,   t_1401,   t_1402;
/* u2_488 Output nets */
wire t_1403,   t_1404,   t_1405;
/* u2_489 Output nets */
wire t_1406,   t_1407,   t_1408;
/* u2_490 Output nets */
wire t_1409,   t_1410,   t_1411;
/* u1_491 Output nets */
wire t_1412,   t_1413;
/* u2_492 Output nets */
wire t_1414,   t_1415,   t_1416;
/* u2_493 Output nets */
wire t_1417,   t_1418,   t_1419;
/* u2_494 Output nets */
wire t_1420,   t_1421,   t_1422;
/* u2_495 Output nets */
wire t_1423,   t_1424,   t_1425;
/* u1_496 Output nets */
wire t_1426,   t_1427;
/* u2_497 Output nets */
wire t_1428,   t_1429,   t_1430;
/* u2_498 Output nets */
wire t_1431,   t_1432,   t_1433;
/* u2_499 Output nets */
wire t_1434,   t_1435,   t_1436;
/* u2_500 Output nets */
wire t_1437,   t_1438,   t_1439;
/* u1_501 Output nets */
wire t_1440,   t_1441;
/* u2_502 Output nets */
wire t_1442,   t_1443,   t_1444;
/* u2_503 Output nets */
wire t_1445,   t_1446,   t_1447;
/* u2_504 Output nets */
wire t_1448,   t_1449,   t_1450;
/* u2_505 Output nets */
wire t_1451,   t_1452,   t_1453;
/* u0_506 Output nets */
wire t_1454,   t_1455;
/* u2_507 Output nets */
wire t_1456,   t_1457,   t_1458;
/* u2_508 Output nets */
wire t_1459,   t_1460,   t_1461;
/* u2_509 Output nets */
wire t_1462,   t_1463,   t_1464;
/* u2_510 Output nets */
wire t_1465,   t_1466,   t_1467;
/* u0_511 Output nets */
wire t_1468,   t_1469;
/* u2_512 Output nets */
wire t_1470,   t_1471,   t_1472;
/* u2_513 Output nets */
wire t_1473,   t_1474,   t_1475;
/* u2_514 Output nets */
wire t_1476,   t_1477,   t_1478;
/* u2_515 Output nets */
wire t_1479,   t_1480,   t_1481;
/* u2_516 Output nets */
wire t_1482,   t_1483,   t_1484;
/* u2_517 Output nets */
wire t_1485,   t_1486,   t_1487;
/* u2_518 Output nets */
wire t_1488,   t_1489,   t_1490;
/* u2_519 Output nets */
wire t_1491,   t_1492,   t_1493;
/* u2_520 Output nets */
wire t_1494,   t_1495,   t_1496;
/* u2_521 Output nets */
wire t_1497,   t_1498,   t_1499;
/* u2_522 Output nets */
wire t_1500,   t_1501,   t_1502;
/* u1_523 Output nets */
wire t_1503,   t_1504;
/* u2_524 Output nets */
wire t_1505,   t_1506,   t_1507;
/* u2_525 Output nets */
wire t_1508,   t_1509,   t_1510;
/* u2_526 Output nets */
wire t_1511,   t_1512,   t_1513;
/* u1_527 Output nets */
wire t_1514,   t_1515;
/* u2_528 Output nets */
wire t_1516,   t_1517,   t_1518;
/* u2_529 Output nets */
wire t_1519,   t_1520,   t_1521;
/* u2_530 Output nets */
wire t_1522,   t_1523,   t_1524;
/* u1_531 Output nets */
wire t_1525,   t_1526;
/* u2_532 Output nets */
wire t_1527,   t_1528,   t_1529;
/* u2_533 Output nets */
wire t_1530,   t_1531,   t_1532;
/* u2_534 Output nets */
wire t_1533,   t_1534,   t_1535;
/* u1_535 Output nets */
wire t_1536,   t_1537;
/* u2_536 Output nets */
wire t_1538,   t_1539,   t_1540;
/* u2_537 Output nets */
wire t_1541,   t_1542,   t_1543;
/* u2_538 Output nets */
wire t_1544,   t_1545,   t_1546;
/* u0_539 Output nets */
wire t_1547,   t_1548;
/* u2_540 Output nets */
wire t_1549,   t_1550,   t_1551;
/* u2_541 Output nets */
wire t_1552,   t_1553,   t_1554;
/* u2_542 Output nets */
wire t_1555,   t_1556,   t_1557;
/* u0_543 Output nets */
wire t_1558,   t_1559;
/* u2_544 Output nets */
wire t_1560,   t_1561,   t_1562;
/* u2_545 Output nets */
wire t_1563,   t_1564,   t_1565;
/* u2_546 Output nets */
wire t_1566,   t_1567,   t_1568;
/* u2_547 Output nets */
wire t_1569,   t_1570,   t_1571;
/* u2_548 Output nets */
wire t_1572,   t_1573,   t_1574;
/* u2_549 Output nets */
wire t_1575,   t_1576,   t_1577;
/* u2_550 Output nets */
wire t_1578,   t_1579,   t_1580;
/* u2_551 Output nets */
wire t_1581,   t_1582,   t_1583;
/* u1_552 Output nets */
wire t_1584,   t_1585;
/* u2_553 Output nets */
wire t_1586,   t_1587,   t_1588;
/* u2_554 Output nets */
wire t_1589,   t_1590,   t_1591;
/* u1_555 Output nets */
wire t_1592,   t_1593;
/* u2_556 Output nets */
wire t_1594,   t_1595,   t_1596;
/* u2_557 Output nets */
wire t_1597,   t_1598,   t_1599;
/* u1_558 Output nets */
wire t_1600,   t_1601;
/* u2_559 Output nets */
wire t_1602,   t_1603,   t_1604;
/* u2_560 Output nets */
wire t_1605,   t_1606,   t_1607;
/* u1_561 Output nets */
wire t_1608,   t_1609;
/* u2_562 Output nets */
wire t_1610,   t_1611,   t_1612;
/* u2_563 Output nets */
wire t_1613,   t_1614,   t_1615;
/* u0_564 Output nets */
wire t_1616,   t_1617;
/* u2_565 Output nets */
wire t_1618,   t_1619,   t_1620;
/* u2_566 Output nets */
wire t_1621,   t_1622,   t_1623;
/* u0_567 Output nets */
wire t_1624,   t_1625;
/* u2_568 Output nets */
wire t_1626,   t_1627,   t_1628;
/* u2_569 Output nets */
wire t_1629,   t_1630,   t_1631;
/* u2_570 Output nets */
wire t_1632,   t_1633,   t_1634;
/* u2_571 Output nets */
wire t_1635,   t_1636,   t_1637;
/* u2_572 Output nets */
wire t_1638,   t_1639,   t_1640;
/* u1_573 Output nets */
wire t_1641,   t_1642;
/* u2_574 Output nets */
wire t_1643,   t_1644,   t_1645;
/* u1_575 Output nets */
wire t_1646,   t_1647;
/* u2_576 Output nets */
wire t_1648,   t_1649,   t_1650;
/* u1_577 Output nets */
wire t_1651,   t_1652;
/* u2_578 Output nets */
wire t_1653,   t_1654,   t_1655;
/* u1_579 Output nets */
wire t_1656,   t_1657;
/* u2_580 Output nets */
wire t_1658,   t_1659,   t_1660;
/* u0_581 Output nets */
wire t_1661,   t_1662;
/* u2_582 Output nets */
wire t_1663,   t_1664,   t_1665;
/* u0_583 Output nets */
wire t_1666,   t_1667;
/* u2_584 Output nets */
wire t_1668,   t_1669,   t_1670;
/* u2_585 Output nets */
wire t_1671,   t_1672,   t_1673;
/* u1_586 Output nets */
wire t_1674,   t_1675;
/* u1_587 Output nets */
wire t_1676,   t_1677;
/* u0_588 Output nets */
wire t_1678,   t_1679;
/* u0_589 Output nets */
wire t_1680;

/* compress stage 1 */
half_adder u0_1(.a(s_0_1), .b(s_0_0), .o(t_0), .cout(t_1));
compressor_3_2 u1_2(.a(s_2_2), .b(s_2_1), .cin(s_2_0), .o(t_2), .cout(t_3));
half_adder u0_3(.a(s_3_1), .b(s_3_0), .o(t_4), .cout(t_5));
compressor_4_2 u2_4(.a(s_4_3), .b(s_4_2), .c(s_4_1), .d(s_4_0), .cin(t_5), .o(t_6), .co(t_7), .cout(t_8));
compressor_3_2 u1_5(.a(s_5_1), .b(s_5_0), .cin(t_8), .o(t_9), .cout(t_10));
compressor_4_2 u2_6(.a(s_6_4), .b(s_6_3), .c(s_6_2), .d(s_6_1), .cin(s_6_0), .o(t_11), .co(t_12), .cout(t_13));
compressor_4_2 u2_7(.a(s_7_3), .b(s_7_2), .c(s_7_1), .d(s_7_0), .cin(t_13), .o(t_14), .co(t_15), .cout(t_16));
compressor_4_2 u2_8(.a(s_8_3), .b(s_8_2), .c(s_8_1), .d(s_8_0), .cin(t_16), .o(t_17), .co(t_18), .cout(t_19));
half_adder u0_9(.a(s_8_5), .b(s_8_4), .o(t_20), .cout(t_21));
compressor_4_2 u2_10(.a(s_9_2), .b(s_9_1), .c(s_9_0), .d(t_19), .cin(t_21), .o(t_22), .co(t_23), .cout(t_24));
half_adder u0_11(.a(s_9_4), .b(s_9_3), .o(t_25), .cout(t_26));
compressor_4_2 u2_12(.a(s_10_2), .b(s_10_1), .c(s_10_0), .d(t_24), .cin(t_26), .o(t_27), .co(t_28), .cout(t_29));
compressor_3_2 u1_13(.a(s_10_5), .b(s_10_4), .cin(s_10_3), .o(t_30), .cout(t_31));
compressor_4_2 u2_14(.a(s_11_2), .b(s_11_1), .c(s_11_0), .d(t_29), .cin(t_31), .o(t_32), .co(t_33), .cout(t_34));
compressor_3_2 u1_15(.a(s_11_5), .b(s_11_4), .cin(s_11_3), .o(t_35), .cout(t_36));
compressor_4_2 u2_16(.a(s_12_2), .b(s_12_1), .c(s_12_0), .d(t_34), .cin(t_36), .o(t_37), .co(t_38), .cout(t_39));
compressor_4_2 u2_17(.a(s_12_7), .b(s_12_6), .c(s_12_5), .d(s_12_4), .cin(s_12_3), .o(t_40), .co(t_41), .cout(t_42));
compressor_4_2 u2_18(.a(s_13_2), .b(s_13_1), .c(s_13_0), .d(t_39), .cin(t_42), .o(t_43), .co(t_44), .cout(t_45));
compressor_3_2 u1_19(.a(s_13_5), .b(s_13_4), .cin(s_13_3), .o(t_46), .cout(t_47));
compressor_4_2 u2_20(.a(s_14_2), .b(s_14_1), .c(s_14_0), .d(t_45), .cin(t_47), .o(t_48), .co(t_49), .cout(t_50));
compressor_4_2 u2_21(.a(s_14_7), .b(s_14_6), .c(s_14_5), .d(s_14_4), .cin(s_14_3), .o(t_51), .co(t_52), .cout(t_53));
compressor_4_2 u2_22(.a(s_15_2), .b(s_15_1), .c(s_15_0), .d(t_50), .cin(t_53), .o(t_54), .co(t_55), .cout(t_56));
compressor_4_2 u2_23(.a(s_15_7), .b(s_15_6), .c(s_15_5), .d(s_15_4), .cin(s_15_3), .o(t_57), .co(t_58), .cout(t_59));
compressor_4_2 u2_24(.a(s_16_2), .b(s_16_1), .c(s_16_0), .d(t_56), .cin(t_59), .o(t_60), .co(t_61), .cout(t_62));
compressor_4_2 u2_25(.a(s_16_7), .b(s_16_6), .c(s_16_5), .d(s_16_4), .cin(s_16_3), .o(t_63), .co(t_64), .cout(t_65));
half_adder u0_26(.a(s_16_9), .b(s_16_8), .o(t_66), .cout(t_67));
compressor_4_2 u2_27(.a(s_17_2), .b(s_17_1), .c(s_17_0), .d(t_62), .cin(t_65), .o(t_68), .co(t_69), .cout(t_70));
compressor_4_2 u2_28(.a(s_17_6), .b(s_17_5), .c(s_17_4), .d(s_17_3), .cin(t_67), .o(t_71), .co(t_72), .cout(t_73));
half_adder u0_29(.a(s_17_8), .b(s_17_7), .o(t_74), .cout(t_75));
compressor_4_2 u2_30(.a(s_18_2), .b(s_18_1), .c(s_18_0), .d(t_70), .cin(t_73), .o(t_76), .co(t_77), .cout(t_78));
compressor_4_2 u2_31(.a(s_18_6), .b(s_18_5), .c(s_18_4), .d(s_18_3), .cin(t_75), .o(t_79), .co(t_80), .cout(t_81));
compressor_3_2 u1_32(.a(s_18_9), .b(s_18_8), .cin(s_18_7), .o(t_82), .cout(t_83));
compressor_4_2 u2_33(.a(s_19_2), .b(s_19_1), .c(s_19_0), .d(t_78), .cin(t_81), .o(t_84), .co(t_85), .cout(t_86));
compressor_4_2 u2_34(.a(s_19_6), .b(s_19_5), .c(s_19_4), .d(s_19_3), .cin(t_83), .o(t_87), .co(t_88), .cout(t_89));
compressor_3_2 u1_35(.a(s_19_9), .b(s_19_8), .cin(s_19_7), .o(t_90), .cout(t_91));
compressor_4_2 u2_36(.a(s_20_2), .b(s_20_1), .c(s_20_0), .d(t_86), .cin(t_89), .o(t_92), .co(t_93), .cout(t_94));
compressor_4_2 u2_37(.a(s_20_6), .b(s_20_5), .c(s_20_4), .d(s_20_3), .cin(t_91), .o(t_95), .co(t_96), .cout(t_97));
compressor_4_2 u2_38(.a(s_20_11), .b(s_20_10), .c(s_20_9), .d(s_20_8), .cin(s_20_7), .o(t_98), .co(t_99), .cout(t_100));
compressor_4_2 u2_39(.a(s_21_2), .b(s_21_1), .c(s_21_0), .d(t_94), .cin(t_97), .o(t_101), .co(t_102), .cout(t_103));
compressor_4_2 u2_40(.a(s_21_6), .b(s_21_5), .c(s_21_4), .d(s_21_3), .cin(t_100), .o(t_104), .co(t_105), .cout(t_106));
compressor_3_2 u1_41(.a(s_21_9), .b(s_21_8), .cin(s_21_7), .o(t_107), .cout(t_108));
compressor_4_2 u2_42(.a(s_22_2), .b(s_22_1), .c(s_22_0), .d(t_103), .cin(t_106), .o(t_109), .co(t_110), .cout(t_111));
compressor_4_2 u2_43(.a(s_22_6), .b(s_22_5), .c(s_22_4), .d(s_22_3), .cin(t_108), .o(t_112), .co(t_113), .cout(t_114));
compressor_4_2 u2_44(.a(s_22_11), .b(s_22_10), .c(s_22_9), .d(s_22_8), .cin(s_22_7), .o(t_115), .co(t_116), .cout(t_117));
compressor_4_2 u2_45(.a(s_23_2), .b(s_23_1), .c(s_23_0), .d(t_111), .cin(t_114), .o(t_118), .co(t_119), .cout(t_120));
compressor_4_2 u2_46(.a(s_23_6), .b(s_23_5), .c(s_23_4), .d(s_23_3), .cin(t_117), .o(t_121), .co(t_122), .cout(t_123));
compressor_4_2 u2_47(.a(s_23_11), .b(s_23_10), .c(s_23_9), .d(s_23_8), .cin(s_23_7), .o(t_124), .co(t_125), .cout(t_126));
compressor_4_2 u2_48(.a(s_24_2), .b(s_24_1), .c(s_24_0), .d(t_120), .cin(t_123), .o(t_127), .co(t_128), .cout(t_129));
compressor_4_2 u2_49(.a(s_24_6), .b(s_24_5), .c(s_24_4), .d(s_24_3), .cin(t_126), .o(t_130), .co(t_131), .cout(t_132));
compressor_4_2 u2_50(.a(s_24_11), .b(s_24_10), .c(s_24_9), .d(s_24_8), .cin(s_24_7), .o(t_133), .co(t_134), .cout(t_135));
half_adder u0_51(.a(s_24_13), .b(s_24_12), .o(t_136), .cout(t_137));
compressor_4_2 u2_52(.a(s_25_2), .b(s_25_1), .c(s_25_0), .d(t_129), .cin(t_132), .o(t_138), .co(t_139), .cout(t_140));
compressor_4_2 u2_53(.a(s_25_5), .b(s_25_4), .c(s_25_3), .d(t_135), .cin(t_137), .o(t_141), .co(t_142), .cout(t_143));
compressor_4_2 u2_54(.a(s_25_10), .b(s_25_9), .c(s_25_8), .d(s_25_7), .cin(s_25_6), .o(t_144), .co(t_145), .cout(t_146));
half_adder u0_55(.a(s_25_12), .b(s_25_11), .o(t_147), .cout(t_148));
compressor_4_2 u2_56(.a(s_26_2), .b(s_26_1), .c(s_26_0), .d(t_140), .cin(t_143), .o(t_149), .co(t_150), .cout(t_151));
compressor_4_2 u2_57(.a(s_26_5), .b(s_26_4), .c(s_26_3), .d(t_146), .cin(t_148), .o(t_152), .co(t_153), .cout(t_154));
compressor_4_2 u2_58(.a(s_26_10), .b(s_26_9), .c(s_26_8), .d(s_26_7), .cin(s_26_6), .o(t_155), .co(t_156), .cout(t_157));
compressor_3_2 u1_59(.a(s_26_13), .b(s_26_12), .cin(s_26_11), .o(t_158), .cout(t_159));
compressor_4_2 u2_60(.a(s_27_2), .b(s_27_1), .c(s_27_0), .d(t_151), .cin(t_154), .o(t_160), .co(t_161), .cout(t_162));
compressor_4_2 u2_61(.a(s_27_5), .b(s_27_4), .c(s_27_3), .d(t_157), .cin(t_159), .o(t_163), .co(t_164), .cout(t_165));
compressor_4_2 u2_62(.a(s_27_10), .b(s_27_9), .c(s_27_8), .d(s_27_7), .cin(s_27_6), .o(t_166), .co(t_167), .cout(t_168));
compressor_3_2 u1_63(.a(s_27_13), .b(s_27_12), .cin(s_27_11), .o(t_169), .cout(t_170));
compressor_4_2 u2_64(.a(s_28_2), .b(s_28_1), .c(s_28_0), .d(t_162), .cin(t_165), .o(t_171), .co(t_172), .cout(t_173));
compressor_4_2 u2_65(.a(s_28_5), .b(s_28_4), .c(s_28_3), .d(t_168), .cin(t_170), .o(t_174), .co(t_175), .cout(t_176));
compressor_4_2 u2_66(.a(s_28_10), .b(s_28_9), .c(s_28_8), .d(s_28_7), .cin(s_28_6), .o(t_177), .co(t_178), .cout(t_179));
compressor_4_2 u2_67(.a(s_28_15), .b(s_28_14), .c(s_28_13), .d(s_28_12), .cin(s_28_11), .o(t_180), .co(t_181), .cout(t_182));
compressor_4_2 u2_68(.a(s_29_2), .b(s_29_1), .c(s_29_0), .d(t_173), .cin(t_176), .o(t_183), .co(t_184), .cout(t_185));
compressor_4_2 u2_69(.a(s_29_5), .b(s_29_4), .c(s_29_3), .d(t_179), .cin(t_182), .o(t_186), .co(t_187), .cout(t_188));
compressor_4_2 u2_70(.a(s_29_10), .b(s_29_9), .c(s_29_8), .d(s_29_7), .cin(s_29_6), .o(t_189), .co(t_190), .cout(t_191));
compressor_3_2 u1_71(.a(s_29_13), .b(s_29_12), .cin(s_29_11), .o(t_192), .cout(t_193));
compressor_4_2 u2_72(.a(s_30_2), .b(s_30_1), .c(s_30_0), .d(t_185), .cin(t_188), .o(t_194), .co(t_195), .cout(t_196));
compressor_4_2 u2_73(.a(s_30_5), .b(s_30_4), .c(s_30_3), .d(t_191), .cin(t_193), .o(t_197), .co(t_198), .cout(t_199));
compressor_4_2 u2_74(.a(s_30_10), .b(s_30_9), .c(s_30_8), .d(s_30_7), .cin(s_30_6), .o(t_200), .co(t_201), .cout(t_202));
compressor_4_2 u2_75(.a(s_30_15), .b(s_30_14), .c(s_30_13), .d(s_30_12), .cin(s_30_11), .o(t_203), .co(t_204), .cout(t_205));
compressor_4_2 u2_76(.a(s_31_2), .b(s_31_1), .c(s_31_0), .d(t_196), .cin(t_199), .o(t_206), .co(t_207), .cout(t_208));
compressor_4_2 u2_77(.a(s_31_5), .b(s_31_4), .c(s_31_3), .d(t_202), .cin(t_205), .o(t_209), .co(t_210), .cout(t_211));
compressor_4_2 u2_78(.a(s_31_10), .b(s_31_9), .c(s_31_8), .d(s_31_7), .cin(s_31_6), .o(t_212), .co(t_213), .cout(t_214));
compressor_4_2 u2_79(.a(s_31_15), .b(s_31_14), .c(s_31_13), .d(s_31_12), .cin(s_31_11), .o(t_215), .co(t_216), .cout(t_217));
compressor_4_2 u2_80(.a(s_32_2), .b(s_32_1), .c(s_32_0), .d(t_208), .cin(t_211), .o(t_218), .co(t_219), .cout(t_220));
compressor_4_2 u2_81(.a(s_32_5), .b(s_32_4), .c(s_32_3), .d(t_214), .cin(t_217), .o(t_221), .co(t_222), .cout(t_223));
compressor_4_2 u2_82(.a(s_32_10), .b(s_32_9), .c(s_32_8), .d(s_32_7), .cin(s_32_6), .o(t_224), .co(t_225), .cout(t_226));
compressor_4_2 u2_83(.a(s_32_15), .b(s_32_14), .c(s_32_13), .d(s_32_12), .cin(s_32_11), .o(t_227), .co(t_228), .cout(t_229));
half_adder u0_84(.a(s_32_17), .b(s_32_16), .o(t_230), .cout(t_231));
compressor_4_2 u2_85(.a(s_33_2), .b(s_33_1), .c(s_33_0), .d(t_220), .cin(t_223), .o(t_232), .co(t_233), .cout(t_234));
compressor_4_2 u2_86(.a(s_33_5), .b(s_33_4), .c(s_33_3), .d(t_226), .cin(t_229), .o(t_235), .co(t_236), .cout(t_237));
compressor_4_2 u2_87(.a(s_33_9), .b(s_33_8), .c(s_33_7), .d(s_33_6), .cin(t_231), .o(t_238), .co(t_239), .cout(t_240));
compressor_4_2 u2_88(.a(s_33_14), .b(s_33_13), .c(s_33_12), .d(s_33_11), .cin(s_33_10), .o(t_241), .co(t_242), .cout(t_243));
half_adder u0_89(.a(s_33_16), .b(s_33_15), .o(t_244), .cout(t_245));
compressor_4_2 u2_90(.a(s_34_2), .b(s_34_1), .c(s_34_0), .d(t_234), .cin(t_237), .o(t_246), .co(t_247), .cout(t_248));
compressor_4_2 u2_91(.a(s_34_5), .b(s_34_4), .c(s_34_3), .d(t_240), .cin(t_243), .o(t_249), .co(t_250), .cout(t_251));
compressor_4_2 u2_92(.a(s_34_9), .b(s_34_8), .c(s_34_7), .d(s_34_6), .cin(t_245), .o(t_252), .co(t_253), .cout(t_254));
compressor_4_2 u2_93(.a(s_34_14), .b(s_34_13), .c(s_34_12), .d(s_34_11), .cin(s_34_10), .o(t_255), .co(t_256), .cout(t_257));
compressor_3_2 u1_94(.a(s_34_17), .b(s_34_16), .cin(s_34_15), .o(t_258), .cout(t_259));
compressor_4_2 u2_95(.a(s_35_2), .b(s_35_1), .c(s_35_0), .d(t_248), .cin(t_251), .o(t_260), .co(t_261), .cout(t_262));
compressor_4_2 u2_96(.a(s_35_5), .b(s_35_4), .c(s_35_3), .d(t_254), .cin(t_257), .o(t_263), .co(t_264), .cout(t_265));
compressor_4_2 u2_97(.a(s_35_9), .b(s_35_8), .c(s_35_7), .d(s_35_6), .cin(t_259), .o(t_266), .co(t_267), .cout(t_268));
compressor_4_2 u2_98(.a(s_35_14), .b(s_35_13), .c(s_35_12), .d(s_35_11), .cin(s_35_10), .o(t_269), .co(t_270), .cout(t_271));
compressor_3_2 u1_99(.a(s_35_17), .b(s_35_16), .cin(s_35_15), .o(t_272), .cout(t_273));
compressor_4_2 u2_100(.a(s_36_2), .b(s_36_1), .c(s_36_0), .d(t_262), .cin(t_265), .o(t_274), .co(t_275), .cout(t_276));
compressor_4_2 u2_101(.a(s_36_5), .b(s_36_4), .c(s_36_3), .d(t_268), .cin(t_271), .o(t_277), .co(t_278), .cout(t_279));
compressor_4_2 u2_102(.a(s_36_9), .b(s_36_8), .c(s_36_7), .d(s_36_6), .cin(t_273), .o(t_280), .co(t_281), .cout(t_282));
compressor_4_2 u2_103(.a(s_36_14), .b(s_36_13), .c(s_36_12), .d(s_36_11), .cin(s_36_10), .o(t_283), .co(t_284), .cout(t_285));
compressor_4_2 u2_104(.a(s_36_19), .b(s_36_18), .c(s_36_17), .d(s_36_16), .cin(s_36_15), .o(t_286), .co(t_287), .cout(t_288));
compressor_4_2 u2_105(.a(s_37_2), .b(s_37_1), .c(s_37_0), .d(t_276), .cin(t_279), .o(t_289), .co(t_290), .cout(t_291));
compressor_4_2 u2_106(.a(s_37_5), .b(s_37_4), .c(s_37_3), .d(t_282), .cin(t_285), .o(t_292), .co(t_293), .cout(t_294));
compressor_4_2 u2_107(.a(s_37_9), .b(s_37_8), .c(s_37_7), .d(s_37_6), .cin(t_288), .o(t_295), .co(t_296), .cout(t_297));
compressor_4_2 u2_108(.a(s_37_14), .b(s_37_13), .c(s_37_12), .d(s_37_11), .cin(s_37_10), .o(t_298), .co(t_299), .cout(t_300));
compressor_3_2 u1_109(.a(s_37_17), .b(s_37_16), .cin(s_37_15), .o(t_301), .cout(t_302));
compressor_4_2 u2_110(.a(s_38_2), .b(s_38_1), .c(s_38_0), .d(t_291), .cin(t_294), .o(t_303), .co(t_304), .cout(t_305));
compressor_4_2 u2_111(.a(s_38_5), .b(s_38_4), .c(s_38_3), .d(t_297), .cin(t_300), .o(t_306), .co(t_307), .cout(t_308));
compressor_4_2 u2_112(.a(s_38_9), .b(s_38_8), .c(s_38_7), .d(s_38_6), .cin(t_302), .o(t_309), .co(t_310), .cout(t_311));
compressor_4_2 u2_113(.a(s_38_14), .b(s_38_13), .c(s_38_12), .d(s_38_11), .cin(s_38_10), .o(t_312), .co(t_313), .cout(t_314));
compressor_4_2 u2_114(.a(s_38_19), .b(s_38_18), .c(s_38_17), .d(s_38_16), .cin(s_38_15), .o(t_315), .co(t_316), .cout(t_317));
compressor_4_2 u2_115(.a(s_39_2), .b(s_39_1), .c(s_39_0), .d(t_305), .cin(t_308), .o(t_318), .co(t_319), .cout(t_320));
compressor_4_2 u2_116(.a(s_39_5), .b(s_39_4), .c(s_39_3), .d(t_311), .cin(t_314), .o(t_321), .co(t_322), .cout(t_323));
compressor_4_2 u2_117(.a(s_39_9), .b(s_39_8), .c(s_39_7), .d(s_39_6), .cin(t_317), .o(t_324), .co(t_325), .cout(t_326));
compressor_4_2 u2_118(.a(s_39_14), .b(s_39_13), .c(s_39_12), .d(s_39_11), .cin(s_39_10), .o(t_327), .co(t_328), .cout(t_329));
compressor_4_2 u2_119(.a(s_39_19), .b(s_39_18), .c(s_39_17), .d(s_39_16), .cin(s_39_15), .o(t_330), .co(t_331), .cout(t_332));
compressor_4_2 u2_120(.a(s_40_2), .b(s_40_1), .c(s_40_0), .d(t_320), .cin(t_323), .o(t_333), .co(t_334), .cout(t_335));
compressor_4_2 u2_121(.a(s_40_5), .b(s_40_4), .c(s_40_3), .d(t_326), .cin(t_329), .o(t_336), .co(t_337), .cout(t_338));
compressor_4_2 u2_122(.a(s_40_9), .b(s_40_8), .c(s_40_7), .d(s_40_6), .cin(t_332), .o(t_339), .co(t_340), .cout(t_341));
compressor_4_2 u2_123(.a(s_40_14), .b(s_40_13), .c(s_40_12), .d(s_40_11), .cin(s_40_10), .o(t_342), .co(t_343), .cout(t_344));
compressor_4_2 u2_124(.a(s_40_19), .b(s_40_18), .c(s_40_17), .d(s_40_16), .cin(s_40_15), .o(t_345), .co(t_346), .cout(t_347));
half_adder u0_125(.a(s_40_21), .b(s_40_20), .o(t_348), .cout(t_349));
compressor_4_2 u2_126(.a(s_41_2), .b(s_41_1), .c(s_41_0), .d(t_335), .cin(t_338), .o(t_350), .co(t_351), .cout(t_352));
compressor_4_2 u2_127(.a(s_41_5), .b(s_41_4), .c(s_41_3), .d(t_341), .cin(t_344), .o(t_353), .co(t_354), .cout(t_355));
compressor_4_2 u2_128(.a(s_41_8), .b(s_41_7), .c(s_41_6), .d(t_347), .cin(t_349), .o(t_356), .co(t_357), .cout(t_358));
compressor_4_2 u2_129(.a(s_41_13), .b(s_41_12), .c(s_41_11), .d(s_41_10), .cin(s_41_9), .o(t_359), .co(t_360), .cout(t_361));
compressor_4_2 u2_130(.a(s_41_18), .b(s_41_17), .c(s_41_16), .d(s_41_15), .cin(s_41_14), .o(t_362), .co(t_363), .cout(t_364));
half_adder u0_131(.a(s_41_20), .b(s_41_19), .o(t_365), .cout(t_366));
compressor_4_2 u2_132(.a(s_42_2), .b(s_42_1), .c(s_42_0), .d(t_352), .cin(t_355), .o(t_367), .co(t_368), .cout(t_369));
compressor_4_2 u2_133(.a(s_42_5), .b(s_42_4), .c(s_42_3), .d(t_358), .cin(t_361), .o(t_370), .co(t_371), .cout(t_372));
compressor_4_2 u2_134(.a(s_42_8), .b(s_42_7), .c(s_42_6), .d(t_364), .cin(t_366), .o(t_373), .co(t_374), .cout(t_375));
compressor_4_2 u2_135(.a(s_42_13), .b(s_42_12), .c(s_42_11), .d(s_42_10), .cin(s_42_9), .o(t_376), .co(t_377), .cout(t_378));
compressor_4_2 u2_136(.a(s_42_18), .b(s_42_17), .c(s_42_16), .d(s_42_15), .cin(s_42_14), .o(t_379), .co(t_380), .cout(t_381));
compressor_3_2 u1_137(.a(s_42_21), .b(s_42_20), .cin(s_42_19), .o(t_382), .cout(t_383));
compressor_4_2 u2_138(.a(s_43_2), .b(s_43_1), .c(s_43_0), .d(t_369), .cin(t_372), .o(t_384), .co(t_385), .cout(t_386));
compressor_4_2 u2_139(.a(s_43_5), .b(s_43_4), .c(s_43_3), .d(t_375), .cin(t_378), .o(t_387), .co(t_388), .cout(t_389));
compressor_4_2 u2_140(.a(s_43_8), .b(s_43_7), .c(s_43_6), .d(t_381), .cin(t_383), .o(t_390), .co(t_391), .cout(t_392));
compressor_4_2 u2_141(.a(s_43_13), .b(s_43_12), .c(s_43_11), .d(s_43_10), .cin(s_43_9), .o(t_393), .co(t_394), .cout(t_395));
compressor_4_2 u2_142(.a(s_43_18), .b(s_43_17), .c(s_43_16), .d(s_43_15), .cin(s_43_14), .o(t_396), .co(t_397), .cout(t_398));
compressor_3_2 u1_143(.a(s_43_21), .b(s_43_20), .cin(s_43_19), .o(t_399), .cout(t_400));
compressor_4_2 u2_144(.a(s_44_2), .b(s_44_1), .c(s_44_0), .d(t_386), .cin(t_389), .o(t_401), .co(t_402), .cout(t_403));
compressor_4_2 u2_145(.a(s_44_5), .b(s_44_4), .c(s_44_3), .d(t_392), .cin(t_395), .o(t_404), .co(t_405), .cout(t_406));
compressor_4_2 u2_146(.a(s_44_8), .b(s_44_7), .c(s_44_6), .d(t_398), .cin(t_400), .o(t_407), .co(t_408), .cout(t_409));
compressor_4_2 u2_147(.a(s_44_13), .b(s_44_12), .c(s_44_11), .d(s_44_10), .cin(s_44_9), .o(t_410), .co(t_411), .cout(t_412));
compressor_4_2 u2_148(.a(s_44_18), .b(s_44_17), .c(s_44_16), .d(s_44_15), .cin(s_44_14), .o(t_413), .co(t_414), .cout(t_415));
compressor_4_2 u2_149(.a(s_44_23), .b(s_44_22), .c(s_44_21), .d(s_44_20), .cin(s_44_19), .o(t_416), .co(t_417), .cout(t_418));
compressor_4_2 u2_150(.a(s_45_2), .b(s_45_1), .c(s_45_0), .d(t_403), .cin(t_406), .o(t_419), .co(t_420), .cout(t_421));
compressor_4_2 u2_151(.a(s_45_5), .b(s_45_4), .c(s_45_3), .d(t_409), .cin(t_412), .o(t_422), .co(t_423), .cout(t_424));
compressor_4_2 u2_152(.a(s_45_8), .b(s_45_7), .c(s_45_6), .d(t_415), .cin(t_418), .o(t_425), .co(t_426), .cout(t_427));
compressor_4_2 u2_153(.a(s_45_13), .b(s_45_12), .c(s_45_11), .d(s_45_10), .cin(s_45_9), .o(t_428), .co(t_429), .cout(t_430));
compressor_4_2 u2_154(.a(s_45_18), .b(s_45_17), .c(s_45_16), .d(s_45_15), .cin(s_45_14), .o(t_431), .co(t_432), .cout(t_433));
compressor_3_2 u1_155(.a(s_45_21), .b(s_45_20), .cin(s_45_19), .o(t_434), .cout(t_435));
compressor_4_2 u2_156(.a(s_46_2), .b(s_46_1), .c(s_46_0), .d(t_421), .cin(t_424), .o(t_436), .co(t_437), .cout(t_438));
compressor_4_2 u2_157(.a(s_46_5), .b(s_46_4), .c(s_46_3), .d(t_427), .cin(t_430), .o(t_439), .co(t_440), .cout(t_441));
compressor_4_2 u2_158(.a(s_46_8), .b(s_46_7), .c(s_46_6), .d(t_433), .cin(t_435), .o(t_442), .co(t_443), .cout(t_444));
compressor_4_2 u2_159(.a(s_46_13), .b(s_46_12), .c(s_46_11), .d(s_46_10), .cin(s_46_9), .o(t_445), .co(t_446), .cout(t_447));
compressor_4_2 u2_160(.a(s_46_18), .b(s_46_17), .c(s_46_16), .d(s_46_15), .cin(s_46_14), .o(t_448), .co(t_449), .cout(t_450));
compressor_4_2 u2_161(.a(s_46_23), .b(s_46_22), .c(s_46_21), .d(s_46_20), .cin(s_46_19), .o(t_451), .co(t_452), .cout(t_453));
compressor_4_2 u2_162(.a(s_47_2), .b(s_47_1), .c(s_47_0), .d(t_438), .cin(t_441), .o(t_454), .co(t_455), .cout(t_456));
compressor_4_2 u2_163(.a(s_47_5), .b(s_47_4), .c(s_47_3), .d(t_444), .cin(t_447), .o(t_457), .co(t_458), .cout(t_459));
compressor_4_2 u2_164(.a(s_47_8), .b(s_47_7), .c(s_47_6), .d(t_450), .cin(t_453), .o(t_460), .co(t_461), .cout(t_462));
compressor_4_2 u2_165(.a(s_47_13), .b(s_47_12), .c(s_47_11), .d(s_47_10), .cin(s_47_9), .o(t_463), .co(t_464), .cout(t_465));
compressor_4_2 u2_166(.a(s_47_18), .b(s_47_17), .c(s_47_16), .d(s_47_15), .cin(s_47_14), .o(t_466), .co(t_467), .cout(t_468));
compressor_4_2 u2_167(.a(s_47_23), .b(s_47_22), .c(s_47_21), .d(s_47_20), .cin(s_47_19), .o(t_469), .co(t_470), .cout(t_471));
compressor_4_2 u2_168(.a(s_48_2), .b(s_48_1), .c(s_48_0), .d(t_456), .cin(t_459), .o(t_472), .co(t_473), .cout(t_474));
compressor_4_2 u2_169(.a(s_48_5), .b(s_48_4), .c(s_48_3), .d(t_462), .cin(t_465), .o(t_475), .co(t_476), .cout(t_477));
compressor_4_2 u2_170(.a(s_48_8), .b(s_48_7), .c(s_48_6), .d(t_468), .cin(t_471), .o(t_478), .co(t_479), .cout(t_480));
compressor_4_2 u2_171(.a(s_48_13), .b(s_48_12), .c(s_48_11), .d(s_48_10), .cin(s_48_9), .o(t_481), .co(t_482), .cout(t_483));
compressor_4_2 u2_172(.a(s_48_18), .b(s_48_17), .c(s_48_16), .d(s_48_15), .cin(s_48_14), .o(t_484), .co(t_485), .cout(t_486));
compressor_4_2 u2_173(.a(s_48_23), .b(s_48_22), .c(s_48_21), .d(s_48_20), .cin(s_48_19), .o(t_487), .co(t_488), .cout(t_489));
half_adder u0_174(.a(s_48_25), .b(s_48_24), .o(t_490), .cout(t_491));
compressor_4_2 u2_175(.a(s_49_2), .b(s_49_1), .c(s_49_0), .d(t_474), .cin(t_477), .o(t_492), .co(t_493), .cout(t_494));
compressor_4_2 u2_176(.a(s_49_5), .b(s_49_4), .c(s_49_3), .d(t_480), .cin(t_483), .o(t_495), .co(t_496), .cout(t_497));
compressor_4_2 u2_177(.a(s_49_8), .b(s_49_7), .c(s_49_6), .d(t_486), .cin(t_489), .o(t_498), .co(t_499), .cout(t_500));
compressor_4_2 u2_178(.a(s_49_12), .b(s_49_11), .c(s_49_10), .d(s_49_9), .cin(t_491), .o(t_501), .co(t_502), .cout(t_503));
compressor_4_2 u2_179(.a(s_49_17), .b(s_49_16), .c(s_49_15), .d(s_49_14), .cin(s_49_13), .o(t_504), .co(t_505), .cout(t_506));
compressor_4_2 u2_180(.a(s_49_22), .b(s_49_21), .c(s_49_20), .d(s_49_19), .cin(s_49_18), .o(t_507), .co(t_508), .cout(t_509));
half_adder u0_181(.a(s_49_24), .b(s_49_23), .o(t_510), .cout(t_511));
compressor_4_2 u2_182(.a(s_50_2), .b(s_50_1), .c(s_50_0), .d(t_494), .cin(t_497), .o(t_512), .co(t_513), .cout(t_514));
compressor_4_2 u2_183(.a(s_50_5), .b(s_50_4), .c(s_50_3), .d(t_500), .cin(t_503), .o(t_515), .co(t_516), .cout(t_517));
compressor_4_2 u2_184(.a(s_50_8), .b(s_50_7), .c(s_50_6), .d(t_506), .cin(t_509), .o(t_518), .co(t_519), .cout(t_520));
compressor_4_2 u2_185(.a(s_50_12), .b(s_50_11), .c(s_50_10), .d(s_50_9), .cin(t_511), .o(t_521), .co(t_522), .cout(t_523));
compressor_4_2 u2_186(.a(s_50_17), .b(s_50_16), .c(s_50_15), .d(s_50_14), .cin(s_50_13), .o(t_524), .co(t_525), .cout(t_526));
compressor_4_2 u2_187(.a(s_50_22), .b(s_50_21), .c(s_50_20), .d(s_50_19), .cin(s_50_18), .o(t_527), .co(t_528), .cout(t_529));
compressor_3_2 u1_188(.a(s_50_25), .b(s_50_24), .cin(s_50_23), .o(t_530), .cout(t_531));
compressor_4_2 u2_189(.a(s_51_2), .b(s_51_1), .c(s_51_0), .d(t_514), .cin(t_517), .o(t_532), .co(t_533), .cout(t_534));
compressor_4_2 u2_190(.a(s_51_5), .b(s_51_4), .c(s_51_3), .d(t_520), .cin(t_523), .o(t_535), .co(t_536), .cout(t_537));
compressor_4_2 u2_191(.a(s_51_8), .b(s_51_7), .c(s_51_6), .d(t_526), .cin(t_529), .o(t_538), .co(t_539), .cout(t_540));
compressor_4_2 u2_192(.a(s_51_12), .b(s_51_11), .c(s_51_10), .d(s_51_9), .cin(t_531), .o(t_541), .co(t_542), .cout(t_543));
compressor_4_2 u2_193(.a(s_51_17), .b(s_51_16), .c(s_51_15), .d(s_51_14), .cin(s_51_13), .o(t_544), .co(t_545), .cout(t_546));
compressor_4_2 u2_194(.a(s_51_22), .b(s_51_21), .c(s_51_20), .d(s_51_19), .cin(s_51_18), .o(t_547), .co(t_548), .cout(t_549));
compressor_3_2 u1_195(.a(s_51_25), .b(s_51_24), .cin(s_51_23), .o(t_550), .cout(t_551));
compressor_4_2 u2_196(.a(s_52_2), .b(s_52_1), .c(s_52_0), .d(t_534), .cin(t_537), .o(t_552), .co(t_553), .cout(t_554));
compressor_4_2 u2_197(.a(s_52_5), .b(s_52_4), .c(s_52_3), .d(t_540), .cin(t_543), .o(t_555), .co(t_556), .cout(t_557));
compressor_4_2 u2_198(.a(s_52_8), .b(s_52_7), .c(s_52_6), .d(t_546), .cin(t_549), .o(t_558), .co(t_559), .cout(t_560));
compressor_4_2 u2_199(.a(s_52_12), .b(s_52_11), .c(s_52_10), .d(s_52_9), .cin(t_551), .o(t_561), .co(t_562), .cout(t_563));
compressor_4_2 u2_200(.a(s_52_17), .b(s_52_16), .c(s_52_15), .d(s_52_14), .cin(s_52_13), .o(t_564), .co(t_565), .cout(t_566));
compressor_4_2 u2_201(.a(s_52_22), .b(s_52_21), .c(s_52_20), .d(s_52_19), .cin(s_52_18), .o(t_567), .co(t_568), .cout(t_569));
compressor_4_2 u2_202(.a(s_52_27), .b(s_52_26), .c(s_52_25), .d(s_52_24), .cin(s_52_23), .o(t_570), .co(t_571), .cout(t_572));
compressor_4_2 u2_203(.a(s_53_2), .b(s_53_1), .c(s_53_0), .d(t_554), .cin(t_557), .o(t_573), .co(t_574), .cout(t_575));
compressor_4_2 u2_204(.a(s_53_5), .b(s_53_4), .c(s_53_3), .d(t_560), .cin(t_563), .o(t_576), .co(t_577), .cout(t_578));
compressor_4_2 u2_205(.a(s_53_8), .b(s_53_7), .c(s_53_6), .d(t_566), .cin(t_569), .o(t_579), .co(t_580), .cout(t_581));
compressor_4_2 u2_206(.a(s_53_12), .b(s_53_11), .c(s_53_10), .d(s_53_9), .cin(t_572), .o(t_582), .co(t_583), .cout(t_584));
compressor_4_2 u2_207(.a(s_53_17), .b(s_53_16), .c(s_53_15), .d(s_53_14), .cin(s_53_13), .o(t_585), .co(t_586), .cout(t_587));
compressor_4_2 u2_208(.a(s_53_22), .b(s_53_21), .c(s_53_20), .d(s_53_19), .cin(s_53_18), .o(t_588), .co(t_589), .cout(t_590));
compressor_3_2 u1_209(.a(s_53_25), .b(s_53_24), .cin(s_53_23), .o(t_591), .cout(t_592));
compressor_4_2 u2_210(.a(s_54_2), .b(s_54_1), .c(s_54_0), .d(t_575), .cin(t_578), .o(t_593), .co(t_594), .cout(t_595));
compressor_4_2 u2_211(.a(s_54_5), .b(s_54_4), .c(s_54_3), .d(t_581), .cin(t_584), .o(t_596), .co(t_597), .cout(t_598));
compressor_4_2 u2_212(.a(s_54_8), .b(s_54_7), .c(s_54_6), .d(t_587), .cin(t_590), .o(t_599), .co(t_600), .cout(t_601));
compressor_4_2 u2_213(.a(s_54_12), .b(s_54_11), .c(s_54_10), .d(s_54_9), .cin(t_592), .o(t_602), .co(t_603), .cout(t_604));
compressor_4_2 u2_214(.a(s_54_17), .b(s_54_16), .c(s_54_15), .d(s_54_14), .cin(s_54_13), .o(t_605), .co(t_606), .cout(t_607));
compressor_4_2 u2_215(.a(s_54_22), .b(s_54_21), .c(s_54_20), .d(s_54_19), .cin(s_54_18), .o(t_608), .co(t_609), .cout(t_610));
compressor_4_2 u2_216(.a(s_54_27), .b(s_54_26), .c(s_54_25), .d(s_54_24), .cin(s_54_23), .o(t_611), .co(t_612), .cout(t_613));
compressor_4_2 u2_217(.a(s_55_2), .b(s_55_1), .c(s_55_0), .d(t_595), .cin(t_598), .o(t_614), .co(t_615), .cout(t_616));
compressor_4_2 u2_218(.a(s_55_5), .b(s_55_4), .c(s_55_3), .d(t_601), .cin(t_604), .o(t_617), .co(t_618), .cout(t_619));
compressor_4_2 u2_219(.a(s_55_8), .b(s_55_7), .c(s_55_6), .d(t_607), .cin(t_610), .o(t_620), .co(t_621), .cout(t_622));
compressor_4_2 u2_220(.a(s_55_12), .b(s_55_11), .c(s_55_10), .d(s_55_9), .cin(t_613), .o(t_623), .co(t_624), .cout(t_625));
compressor_4_2 u2_221(.a(s_55_17), .b(s_55_16), .c(s_55_15), .d(s_55_14), .cin(s_55_13), .o(t_626), .co(t_627), .cout(t_628));
compressor_4_2 u2_222(.a(s_55_22), .b(s_55_21), .c(s_55_20), .d(s_55_19), .cin(s_55_18), .o(t_629), .co(t_630), .cout(t_631));
compressor_4_2 u2_223(.a(s_55_27), .b(s_55_26), .c(s_55_25), .d(s_55_24), .cin(s_55_23), .o(t_632), .co(t_633), .cout(t_634));
compressor_4_2 u2_224(.a(s_56_2), .b(s_56_1), .c(s_56_0), .d(t_616), .cin(t_619), .o(t_635), .co(t_636), .cout(t_637));
compressor_4_2 u2_225(.a(s_56_5), .b(s_56_4), .c(s_56_3), .d(t_622), .cin(t_625), .o(t_638), .co(t_639), .cout(t_640));
compressor_4_2 u2_226(.a(s_56_8), .b(s_56_7), .c(s_56_6), .d(t_628), .cin(t_631), .o(t_641), .co(t_642), .cout(t_643));
compressor_4_2 u2_227(.a(s_56_12), .b(s_56_11), .c(s_56_10), .d(s_56_9), .cin(t_634), .o(t_644), .co(t_645), .cout(t_646));
compressor_4_2 u2_228(.a(s_56_17), .b(s_56_16), .c(s_56_15), .d(s_56_14), .cin(s_56_13), .o(t_647), .co(t_648), .cout(t_649));
compressor_4_2 u2_229(.a(s_56_22), .b(s_56_21), .c(s_56_20), .d(s_56_19), .cin(s_56_18), .o(t_650), .co(t_651), .cout(t_652));
compressor_4_2 u2_230(.a(s_56_27), .b(s_56_26), .c(s_56_25), .d(s_56_24), .cin(s_56_23), .o(t_653), .co(t_654), .cout(t_655));
half_adder u0_231(.a(s_56_29), .b(s_56_28), .o(t_656), .cout(t_657));
compressor_4_2 u2_232(.a(s_57_2), .b(s_57_1), .c(s_57_0), .d(t_637), .cin(t_640), .o(t_658), .co(t_659), .cout(t_660));
compressor_4_2 u2_233(.a(s_57_5), .b(s_57_4), .c(s_57_3), .d(t_643), .cin(t_646), .o(t_661), .co(t_662), .cout(t_663));
compressor_4_2 u2_234(.a(s_57_8), .b(s_57_7), .c(s_57_6), .d(t_649), .cin(t_652), .o(t_664), .co(t_665), .cout(t_666));
compressor_4_2 u2_235(.a(s_57_11), .b(s_57_10), .c(s_57_9), .d(t_655), .cin(t_657), .o(t_667), .co(t_668), .cout(t_669));
compressor_4_2 u2_236(.a(s_57_16), .b(s_57_15), .c(s_57_14), .d(s_57_13), .cin(s_57_12), .o(t_670), .co(t_671), .cout(t_672));
compressor_4_2 u2_237(.a(s_57_21), .b(s_57_20), .c(s_57_19), .d(s_57_18), .cin(s_57_17), .o(t_673), .co(t_674), .cout(t_675));
compressor_4_2 u2_238(.a(s_57_26), .b(s_57_25), .c(s_57_24), .d(s_57_23), .cin(s_57_22), .o(t_676), .co(t_677), .cout(t_678));
half_adder u0_239(.a(s_57_28), .b(s_57_27), .o(t_679), .cout(t_680));
compressor_4_2 u2_240(.a(s_58_2), .b(s_58_1), .c(s_58_0), .d(t_660), .cin(t_663), .o(t_681), .co(t_682), .cout(t_683));
compressor_4_2 u2_241(.a(s_58_5), .b(s_58_4), .c(s_58_3), .d(t_666), .cin(t_669), .o(t_684), .co(t_685), .cout(t_686));
compressor_4_2 u2_242(.a(s_58_8), .b(s_58_7), .c(s_58_6), .d(t_672), .cin(t_675), .o(t_687), .co(t_688), .cout(t_689));
compressor_4_2 u2_243(.a(s_58_11), .b(s_58_10), .c(s_58_9), .d(t_678), .cin(t_680), .o(t_690), .co(t_691), .cout(t_692));
compressor_4_2 u2_244(.a(s_58_16), .b(s_58_15), .c(s_58_14), .d(s_58_13), .cin(s_58_12), .o(t_693), .co(t_694), .cout(t_695));
compressor_4_2 u2_245(.a(s_58_21), .b(s_58_20), .c(s_58_19), .d(s_58_18), .cin(s_58_17), .o(t_696), .co(t_697), .cout(t_698));
compressor_4_2 u2_246(.a(s_58_26), .b(s_58_25), .c(s_58_24), .d(s_58_23), .cin(s_58_22), .o(t_699), .co(t_700), .cout(t_701));
compressor_3_2 u1_247(.a(s_58_29), .b(s_58_28), .cin(s_58_27), .o(t_702), .cout(t_703));
compressor_4_2 u2_248(.a(s_59_2), .b(s_59_1), .c(s_59_0), .d(t_683), .cin(t_686), .o(t_704), .co(t_705), .cout(t_706));
compressor_4_2 u2_249(.a(s_59_5), .b(s_59_4), .c(s_59_3), .d(t_689), .cin(t_692), .o(t_707), .co(t_708), .cout(t_709));
compressor_4_2 u2_250(.a(s_59_8), .b(s_59_7), .c(s_59_6), .d(t_695), .cin(t_698), .o(t_710), .co(t_711), .cout(t_712));
compressor_4_2 u2_251(.a(s_59_11), .b(s_59_10), .c(s_59_9), .d(t_701), .cin(t_703), .o(t_713), .co(t_714), .cout(t_715));
compressor_4_2 u2_252(.a(s_59_16), .b(s_59_15), .c(s_59_14), .d(s_59_13), .cin(s_59_12), .o(t_716), .co(t_717), .cout(t_718));
compressor_4_2 u2_253(.a(s_59_21), .b(s_59_20), .c(s_59_19), .d(s_59_18), .cin(s_59_17), .o(t_719), .co(t_720), .cout(t_721));
compressor_4_2 u2_254(.a(s_59_26), .b(s_59_25), .c(s_59_24), .d(s_59_23), .cin(s_59_22), .o(t_722), .co(t_723), .cout(t_724));
compressor_3_2 u1_255(.a(s_59_29), .b(s_59_28), .cin(s_59_27), .o(t_725), .cout(t_726));
compressor_4_2 u2_256(.a(s_60_2), .b(s_60_1), .c(s_60_0), .d(t_706), .cin(t_709), .o(t_727), .co(t_728), .cout(t_729));
compressor_4_2 u2_257(.a(s_60_5), .b(s_60_4), .c(s_60_3), .d(t_712), .cin(t_715), .o(t_730), .co(t_731), .cout(t_732));
compressor_4_2 u2_258(.a(s_60_8), .b(s_60_7), .c(s_60_6), .d(t_718), .cin(t_721), .o(t_733), .co(t_734), .cout(t_735));
compressor_4_2 u2_259(.a(s_60_11), .b(s_60_10), .c(s_60_9), .d(t_724), .cin(t_726), .o(t_736), .co(t_737), .cout(t_738));
compressor_4_2 u2_260(.a(s_60_16), .b(s_60_15), .c(s_60_14), .d(s_60_13), .cin(s_60_12), .o(t_739), .co(t_740), .cout(t_741));
compressor_4_2 u2_261(.a(s_60_21), .b(s_60_20), .c(s_60_19), .d(s_60_18), .cin(s_60_17), .o(t_742), .co(t_743), .cout(t_744));
compressor_4_2 u2_262(.a(s_60_26), .b(s_60_25), .c(s_60_24), .d(s_60_23), .cin(s_60_22), .o(t_745), .co(t_746), .cout(t_747));
compressor_4_2 u2_263(.a(s_60_31), .b(s_60_30), .c(s_60_29), .d(s_60_28), .cin(s_60_27), .o(t_748), .co(t_749), .cout(t_750));
compressor_4_2 u2_264(.a(s_61_2), .b(s_61_1), .c(s_61_0), .d(t_729), .cin(t_732), .o(t_751), .co(t_752), .cout(t_753));
compressor_4_2 u2_265(.a(s_61_5), .b(s_61_4), .c(s_61_3), .d(t_735), .cin(t_738), .o(t_754), .co(t_755), .cout(t_756));
compressor_4_2 u2_266(.a(s_61_8), .b(s_61_7), .c(s_61_6), .d(t_741), .cin(t_744), .o(t_757), .co(t_758), .cout(t_759));
compressor_4_2 u2_267(.a(s_61_11), .b(s_61_10), .c(s_61_9), .d(t_747), .cin(t_750), .o(t_760), .co(t_761), .cout(t_762));
compressor_4_2 u2_268(.a(s_61_16), .b(s_61_15), .c(s_61_14), .d(s_61_13), .cin(s_61_12), .o(t_763), .co(t_764), .cout(t_765));
compressor_4_2 u2_269(.a(s_61_21), .b(s_61_20), .c(s_61_19), .d(s_61_18), .cin(s_61_17), .o(t_766), .co(t_767), .cout(t_768));
compressor_4_2 u2_270(.a(s_61_26), .b(s_61_25), .c(s_61_24), .d(s_61_23), .cin(s_61_22), .o(t_769), .co(t_770), .cout(t_771));
compressor_3_2 u1_271(.a(s_61_29), .b(s_61_28), .cin(s_61_27), .o(t_772), .cout(t_773));
compressor_4_2 u2_272(.a(s_62_2), .b(s_62_1), .c(s_62_0), .d(t_753), .cin(t_756), .o(t_774), .co(t_775), .cout(t_776));
compressor_4_2 u2_273(.a(s_62_5), .b(s_62_4), .c(s_62_3), .d(t_759), .cin(t_762), .o(t_777), .co(t_778), .cout(t_779));
compressor_4_2 u2_274(.a(s_62_8), .b(s_62_7), .c(s_62_6), .d(t_765), .cin(t_768), .o(t_780), .co(t_781), .cout(t_782));
compressor_4_2 u2_275(.a(s_62_11), .b(s_62_10), .c(s_62_9), .d(t_771), .cin(t_773), .o(t_783), .co(t_784), .cout(t_785));
compressor_4_2 u2_276(.a(s_62_16), .b(s_62_15), .c(s_62_14), .d(s_62_13), .cin(s_62_12), .o(t_786), .co(t_787), .cout(t_788));
compressor_4_2 u2_277(.a(s_62_21), .b(s_62_20), .c(s_62_19), .d(s_62_18), .cin(s_62_17), .o(t_789), .co(t_790), .cout(t_791));
compressor_4_2 u2_278(.a(s_62_26), .b(s_62_25), .c(s_62_24), .d(s_62_23), .cin(s_62_22), .o(t_792), .co(t_793), .cout(t_794));
compressor_4_2 u2_279(.a(s_62_31), .b(s_62_30), .c(s_62_29), .d(s_62_28), .cin(s_62_27), .o(t_795), .co(t_796), .cout(t_797));
compressor_4_2 u2_280(.a(s_63_2), .b(s_63_1), .c(s_63_0), .d(t_776), .cin(t_779), .o(t_798), .co(t_799), .cout(t_800));
compressor_4_2 u2_281(.a(s_63_5), .b(s_63_4), .c(s_63_3), .d(t_782), .cin(t_785), .o(t_801), .co(t_802), .cout(t_803));
compressor_4_2 u2_282(.a(s_63_8), .b(s_63_7), .c(s_63_6), .d(t_788), .cin(t_791), .o(t_804), .co(t_805), .cout(t_806));
compressor_4_2 u2_283(.a(s_63_11), .b(s_63_10), .c(s_63_9), .d(t_794), .cin(t_797), .o(t_807), .co(t_808), .cout(t_809));
compressor_4_2 u2_284(.a(s_63_16), .b(s_63_15), .c(s_63_14), .d(s_63_13), .cin(s_63_12), .o(t_810), .co(t_811), .cout(t_812));
compressor_4_2 u2_285(.a(s_63_21), .b(s_63_20), .c(s_63_19), .d(s_63_18), .cin(s_63_17), .o(t_813), .co(t_814), .cout(t_815));
compressor_4_2 u2_286(.a(s_63_26), .b(s_63_25), .c(s_63_24), .d(s_63_23), .cin(s_63_22), .o(t_816), .co(t_817), .cout(t_818));
compressor_4_2 u2_287(.a(s_63_31), .b(s_63_30), .c(s_63_29), .d(s_63_28), .cin(s_63_27), .o(t_819), .co(t_820), .cout(t_821));
compressor_4_2 u2_288(.a(s_64_2), .b(s_64_1), .c(s_64_0), .d(t_800), .cin(t_803), .o(t_822), .co(t_823), .cout(t_824));
compressor_4_2 u2_289(.a(s_64_5), .b(s_64_4), .c(s_64_3), .d(t_806), .cin(t_809), .o(t_825), .co(t_826), .cout(t_827));
compressor_4_2 u2_290(.a(s_64_8), .b(s_64_7), .c(s_64_6), .d(t_812), .cin(t_815), .o(t_828), .co(t_829), .cout(t_830));
compressor_4_2 u2_291(.a(s_64_11), .b(s_64_10), .c(s_64_9), .d(t_818), .cin(t_821), .o(t_831), .co(t_832), .cout(t_833));
compressor_4_2 u2_292(.a(s_64_16), .b(s_64_15), .c(s_64_14), .d(s_64_13), .cin(s_64_12), .o(t_834), .co(t_835), .cout(t_836));
compressor_4_2 u2_293(.a(s_64_21), .b(s_64_20), .c(s_64_19), .d(s_64_18), .cin(s_64_17), .o(t_837), .co(t_838), .cout(t_839));
compressor_4_2 u2_294(.a(s_64_26), .b(s_64_25), .c(s_64_24), .d(s_64_23), .cin(s_64_22), .o(t_840), .co(t_841), .cout(t_842));
compressor_4_2 u2_295(.a(s_64_31), .b(s_64_30), .c(s_64_29), .d(s_64_28), .cin(s_64_27), .o(t_843), .co(t_844), .cout(t_845));
compressor_4_2 u2_296(.a(s_65_2), .b(s_65_1), .c(s_65_0), .d(t_824), .cin(t_827), .o(t_846), .co(t_847), .cout(t_848));
compressor_4_2 u2_297(.a(s_65_5), .b(s_65_4), .c(s_65_3), .d(t_830), .cin(t_833), .o(t_849), .co(t_850), .cout(t_851));
compressor_4_2 u2_298(.a(s_65_8), .b(s_65_7), .c(s_65_6), .d(t_836), .cin(t_839), .o(t_852), .co(t_853), .cout(t_854));
compressor_4_2 u2_299(.a(s_65_11), .b(s_65_10), .c(s_65_9), .d(t_842), .cin(t_845), .o(t_855), .co(t_856), .cout(t_857));
compressor_4_2 u2_300(.a(s_65_16), .b(s_65_15), .c(s_65_14), .d(s_65_13), .cin(s_65_12), .o(t_858), .co(t_859), .cout(t_860));
compressor_4_2 u2_301(.a(s_65_21), .b(s_65_20), .c(s_65_19), .d(s_65_18), .cin(s_65_17), .o(t_861), .co(t_862), .cout(t_863));
compressor_4_2 u2_302(.a(s_65_26), .b(s_65_25), .c(s_65_24), .d(s_65_23), .cin(s_65_22), .o(t_864), .co(t_865), .cout(t_866));
compressor_4_2 u2_303(.a(s_65_31), .b(s_65_30), .c(s_65_29), .d(s_65_28), .cin(s_65_27), .o(t_867), .co(t_868), .cout(t_869));
compressor_4_2 u2_304(.a(s_66_2), .b(s_66_1), .c(s_66_0), .d(t_848), .cin(t_851), .o(t_870), .co(t_871), .cout(t_872));
compressor_4_2 u2_305(.a(s_66_5), .b(s_66_4), .c(s_66_3), .d(t_854), .cin(t_857), .o(t_873), .co(t_874), .cout(t_875));
compressor_4_2 u2_306(.a(s_66_8), .b(s_66_7), .c(s_66_6), .d(t_860), .cin(t_863), .o(t_876), .co(t_877), .cout(t_878));
compressor_4_2 u2_307(.a(s_66_11), .b(s_66_10), .c(s_66_9), .d(t_866), .cin(t_869), .o(t_879), .co(t_880), .cout(t_881));
compressor_4_2 u2_308(.a(s_66_16), .b(s_66_15), .c(s_66_14), .d(s_66_13), .cin(s_66_12), .o(t_882), .co(t_883), .cout(t_884));
compressor_4_2 u2_309(.a(s_66_21), .b(s_66_20), .c(s_66_19), .d(s_66_18), .cin(s_66_17), .o(t_885), .co(t_886), .cout(t_887));
compressor_4_2 u2_310(.a(s_66_26), .b(s_66_25), .c(s_66_24), .d(s_66_23), .cin(s_66_22), .o(t_888), .co(t_889), .cout(t_890));
compressor_4_2 u2_311(.a(s_66_31), .b(s_66_30), .c(s_66_29), .d(s_66_28), .cin(s_66_27), .o(t_891), .co(t_892), .cout(t_893));
compressor_4_2 u2_312(.a(s_67_2), .b(s_67_1), .c(s_67_0), .d(t_872), .cin(t_875), .o(t_894), .co(t_895), .cout(t_896));
compressor_4_2 u2_313(.a(s_67_5), .b(s_67_4), .c(s_67_3), .d(t_878), .cin(t_881), .o(t_897), .co(t_898), .cout(t_899));
compressor_4_2 u2_314(.a(s_67_8), .b(s_67_7), .c(s_67_6), .d(t_884), .cin(t_887), .o(t_900), .co(t_901), .cout(t_902));
compressor_4_2 u2_315(.a(s_67_11), .b(s_67_10), .c(s_67_9), .d(t_890), .cin(t_893), .o(t_903), .co(t_904), .cout(t_905));
compressor_4_2 u2_316(.a(s_67_16), .b(s_67_15), .c(s_67_14), .d(s_67_13), .cin(s_67_12), .o(t_906), .co(t_907), .cout(t_908));
compressor_4_2 u2_317(.a(s_67_21), .b(s_67_20), .c(s_67_19), .d(s_67_18), .cin(s_67_17), .o(t_909), .co(t_910), .cout(t_911));
compressor_4_2 u2_318(.a(s_67_26), .b(s_67_25), .c(s_67_24), .d(s_67_23), .cin(s_67_22), .o(t_912), .co(t_913), .cout(t_914));
compressor_4_2 u2_319(.a(s_67_31), .b(s_67_30), .c(s_67_29), .d(s_67_28), .cin(s_67_27), .o(t_915), .co(t_916), .cout(t_917));
compressor_4_2 u2_320(.a(s_68_2), .b(s_68_1), .c(s_68_0), .d(t_896), .cin(t_899), .o(t_918), .co(t_919), .cout(t_920));
compressor_4_2 u2_321(.a(s_68_5), .b(s_68_4), .c(s_68_3), .d(t_902), .cin(t_905), .o(t_921), .co(t_922), .cout(t_923));
compressor_4_2 u2_322(.a(s_68_8), .b(s_68_7), .c(s_68_6), .d(t_908), .cin(t_911), .o(t_924), .co(t_925), .cout(t_926));
compressor_4_2 u2_323(.a(s_68_11), .b(s_68_10), .c(s_68_9), .d(t_914), .cin(t_917), .o(t_927), .co(t_928), .cout(t_929));
compressor_4_2 u2_324(.a(s_68_16), .b(s_68_15), .c(s_68_14), .d(s_68_13), .cin(s_68_12), .o(t_930), .co(t_931), .cout(t_932));
compressor_4_2 u2_325(.a(s_68_21), .b(s_68_20), .c(s_68_19), .d(s_68_18), .cin(s_68_17), .o(t_933), .co(t_934), .cout(t_935));
compressor_4_2 u2_326(.a(s_68_26), .b(s_68_25), .c(s_68_24), .d(s_68_23), .cin(s_68_22), .o(t_936), .co(t_937), .cout(t_938));
compressor_3_2 u1_327(.a(s_68_29), .b(s_68_28), .cin(s_68_27), .o(t_939), .cout(t_940));
compressor_4_2 u2_328(.a(s_69_2), .b(s_69_1), .c(s_69_0), .d(t_920), .cin(t_923), .o(t_941), .co(t_942), .cout(t_943));
compressor_4_2 u2_329(.a(s_69_5), .b(s_69_4), .c(s_69_3), .d(t_926), .cin(t_929), .o(t_944), .co(t_945), .cout(t_946));
compressor_4_2 u2_330(.a(s_69_8), .b(s_69_7), .c(s_69_6), .d(t_932), .cin(t_935), .o(t_947), .co(t_948), .cout(t_949));
compressor_4_2 u2_331(.a(s_69_11), .b(s_69_10), .c(s_69_9), .d(t_938), .cin(t_940), .o(t_950), .co(t_951), .cout(t_952));
compressor_4_2 u2_332(.a(s_69_16), .b(s_69_15), .c(s_69_14), .d(s_69_13), .cin(s_69_12), .o(t_953), .co(t_954), .cout(t_955));
compressor_4_2 u2_333(.a(s_69_21), .b(s_69_20), .c(s_69_19), .d(s_69_18), .cin(s_69_17), .o(t_956), .co(t_957), .cout(t_958));
compressor_4_2 u2_334(.a(s_69_26), .b(s_69_25), .c(s_69_24), .d(s_69_23), .cin(s_69_22), .o(t_959), .co(t_960), .cout(t_961));
compressor_3_2 u1_335(.a(s_69_29), .b(s_69_28), .cin(s_69_27), .o(t_962), .cout(t_963));
compressor_4_2 u2_336(.a(s_70_2), .b(s_70_1), .c(s_70_0), .d(t_943), .cin(t_946), .o(t_964), .co(t_965), .cout(t_966));
compressor_4_2 u2_337(.a(s_70_5), .b(s_70_4), .c(s_70_3), .d(t_949), .cin(t_952), .o(t_967), .co(t_968), .cout(t_969));
compressor_4_2 u2_338(.a(s_70_8), .b(s_70_7), .c(s_70_6), .d(t_955), .cin(t_958), .o(t_970), .co(t_971), .cout(t_972));
compressor_4_2 u2_339(.a(s_70_11), .b(s_70_10), .c(s_70_9), .d(t_961), .cin(t_963), .o(t_973), .co(t_974), .cout(t_975));
compressor_4_2 u2_340(.a(s_70_16), .b(s_70_15), .c(s_70_14), .d(s_70_13), .cin(s_70_12), .o(t_976), .co(t_977), .cout(t_978));
compressor_4_2 u2_341(.a(s_70_21), .b(s_70_20), .c(s_70_19), .d(s_70_18), .cin(s_70_17), .o(t_979), .co(t_980), .cout(t_981));
compressor_4_2 u2_342(.a(s_70_26), .b(s_70_25), .c(s_70_24), .d(s_70_23), .cin(s_70_22), .o(t_982), .co(t_983), .cout(t_984));
compressor_3_2 u1_343(.a(s_70_29), .b(s_70_28), .cin(s_70_27), .o(t_985), .cout(t_986));
compressor_4_2 u2_344(.a(s_71_2), .b(s_71_1), .c(s_71_0), .d(t_966), .cin(t_969), .o(t_987), .co(t_988), .cout(t_989));
compressor_4_2 u2_345(.a(s_71_5), .b(s_71_4), .c(s_71_3), .d(t_972), .cin(t_975), .o(t_990), .co(t_991), .cout(t_992));
compressor_4_2 u2_346(.a(s_71_8), .b(s_71_7), .c(s_71_6), .d(t_978), .cin(t_981), .o(t_993), .co(t_994), .cout(t_995));
compressor_4_2 u2_347(.a(s_71_11), .b(s_71_10), .c(s_71_9), .d(t_984), .cin(t_986), .o(t_996), .co(t_997), .cout(t_998));
compressor_4_2 u2_348(.a(s_71_16), .b(s_71_15), .c(s_71_14), .d(s_71_13), .cin(s_71_12), .o(t_999), .co(t_1000), .cout(t_1001));
compressor_4_2 u2_349(.a(s_71_21), .b(s_71_20), .c(s_71_19), .d(s_71_18), .cin(s_71_17), .o(t_1002), .co(t_1003), .cout(t_1004));
compressor_4_2 u2_350(.a(s_71_26), .b(s_71_25), .c(s_71_24), .d(s_71_23), .cin(s_71_22), .o(t_1005), .co(t_1006), .cout(t_1007));
compressor_3_2 u1_351(.a(s_71_29), .b(s_71_28), .cin(s_71_27), .o(t_1008), .cout(t_1009));
compressor_4_2 u2_352(.a(s_72_2), .b(s_72_1), .c(s_72_0), .d(t_989), .cin(t_992), .o(t_1010), .co(t_1011), .cout(t_1012));
compressor_4_2 u2_353(.a(s_72_5), .b(s_72_4), .c(s_72_3), .d(t_995), .cin(t_998), .o(t_1013), .co(t_1014), .cout(t_1015));
compressor_4_2 u2_354(.a(s_72_8), .b(s_72_7), .c(s_72_6), .d(t_1001), .cin(t_1004), .o(t_1016), .co(t_1017), .cout(t_1018));
compressor_4_2 u2_355(.a(s_72_11), .b(s_72_10), .c(s_72_9), .d(t_1007), .cin(t_1009), .o(t_1019), .co(t_1020), .cout(t_1021));
compressor_4_2 u2_356(.a(s_72_16), .b(s_72_15), .c(s_72_14), .d(s_72_13), .cin(s_72_12), .o(t_1022), .co(t_1023), .cout(t_1024));
compressor_4_2 u2_357(.a(s_72_21), .b(s_72_20), .c(s_72_19), .d(s_72_18), .cin(s_72_17), .o(t_1025), .co(t_1026), .cout(t_1027));
compressor_4_2 u2_358(.a(s_72_26), .b(s_72_25), .c(s_72_24), .d(s_72_23), .cin(s_72_22), .o(t_1028), .co(t_1029), .cout(t_1030));
half_adder u0_359(.a(s_72_28), .b(s_72_27), .o(t_1031), .cout(t_1032));
compressor_4_2 u2_360(.a(s_73_2), .b(s_73_1), .c(s_73_0), .d(t_1012), .cin(t_1015), .o(t_1033), .co(t_1034), .cout(t_1035));
compressor_4_2 u2_361(.a(s_73_5), .b(s_73_4), .c(s_73_3), .d(t_1018), .cin(t_1021), .o(t_1036), .co(t_1037), .cout(t_1038));
compressor_4_2 u2_362(.a(s_73_8), .b(s_73_7), .c(s_73_6), .d(t_1024), .cin(t_1027), .o(t_1039), .co(t_1040), .cout(t_1041));
compressor_4_2 u2_363(.a(s_73_11), .b(s_73_10), .c(s_73_9), .d(t_1030), .cin(t_1032), .o(t_1042), .co(t_1043), .cout(t_1044));
compressor_4_2 u2_364(.a(s_73_16), .b(s_73_15), .c(s_73_14), .d(s_73_13), .cin(s_73_12), .o(t_1045), .co(t_1046), .cout(t_1047));
compressor_4_2 u2_365(.a(s_73_21), .b(s_73_20), .c(s_73_19), .d(s_73_18), .cin(s_73_17), .o(t_1048), .co(t_1049), .cout(t_1050));
compressor_4_2 u2_366(.a(s_73_26), .b(s_73_25), .c(s_73_24), .d(s_73_23), .cin(s_73_22), .o(t_1051), .co(t_1052), .cout(t_1053));
half_adder u0_367(.a(s_73_28), .b(s_73_27), .o(t_1054), .cout(t_1055));
compressor_4_2 u2_368(.a(s_74_2), .b(s_74_1), .c(s_74_0), .d(t_1035), .cin(t_1038), .o(t_1056), .co(t_1057), .cout(t_1058));
compressor_4_2 u2_369(.a(s_74_5), .b(s_74_4), .c(s_74_3), .d(t_1041), .cin(t_1044), .o(t_1059), .co(t_1060), .cout(t_1061));
compressor_4_2 u2_370(.a(s_74_8), .b(s_74_7), .c(s_74_6), .d(t_1047), .cin(t_1050), .o(t_1062), .co(t_1063), .cout(t_1064));
compressor_4_2 u2_371(.a(s_74_11), .b(s_74_10), .c(s_74_9), .d(t_1053), .cin(t_1055), .o(t_1065), .co(t_1066), .cout(t_1067));
compressor_4_2 u2_372(.a(s_74_16), .b(s_74_15), .c(s_74_14), .d(s_74_13), .cin(s_74_12), .o(t_1068), .co(t_1069), .cout(t_1070));
compressor_4_2 u2_373(.a(s_74_21), .b(s_74_20), .c(s_74_19), .d(s_74_18), .cin(s_74_17), .o(t_1071), .co(t_1072), .cout(t_1073));
compressor_4_2 u2_374(.a(s_74_26), .b(s_74_25), .c(s_74_24), .d(s_74_23), .cin(s_74_22), .o(t_1074), .co(t_1075), .cout(t_1076));
compressor_4_2 u2_375(.a(s_75_2), .b(s_75_1), .c(s_75_0), .d(t_1058), .cin(t_1061), .o(t_1077), .co(t_1078), .cout(t_1079));
compressor_4_2 u2_376(.a(s_75_5), .b(s_75_4), .c(s_75_3), .d(t_1064), .cin(t_1067), .o(t_1080), .co(t_1081), .cout(t_1082));
compressor_4_2 u2_377(.a(s_75_8), .b(s_75_7), .c(s_75_6), .d(t_1070), .cin(t_1073), .o(t_1083), .co(t_1084), .cout(t_1085));
compressor_4_2 u2_378(.a(s_75_12), .b(s_75_11), .c(s_75_10), .d(s_75_9), .cin(t_1076), .o(t_1086), .co(t_1087), .cout(t_1088));
compressor_4_2 u2_379(.a(s_75_17), .b(s_75_16), .c(s_75_15), .d(s_75_14), .cin(s_75_13), .o(t_1089), .co(t_1090), .cout(t_1091));
compressor_4_2 u2_380(.a(s_75_22), .b(s_75_21), .c(s_75_20), .d(s_75_19), .cin(s_75_18), .o(t_1092), .co(t_1093), .cout(t_1094));
compressor_4_2 u2_381(.a(s_75_27), .b(s_75_26), .c(s_75_25), .d(s_75_24), .cin(s_75_23), .o(t_1095), .co(t_1096), .cout(t_1097));
compressor_4_2 u2_382(.a(s_76_2), .b(s_76_1), .c(s_76_0), .d(t_1079), .cin(t_1082), .o(t_1098), .co(t_1099), .cout(t_1100));
compressor_4_2 u2_383(.a(s_76_5), .b(s_76_4), .c(s_76_3), .d(t_1085), .cin(t_1088), .o(t_1101), .co(t_1102), .cout(t_1103));
compressor_4_2 u2_384(.a(s_76_8), .b(s_76_7), .c(s_76_6), .d(t_1091), .cin(t_1094), .o(t_1104), .co(t_1105), .cout(t_1106));
compressor_4_2 u2_385(.a(s_76_12), .b(s_76_11), .c(s_76_10), .d(s_76_9), .cin(t_1097), .o(t_1107), .co(t_1108), .cout(t_1109));
compressor_4_2 u2_386(.a(s_76_17), .b(s_76_16), .c(s_76_15), .d(s_76_14), .cin(s_76_13), .o(t_1110), .co(t_1111), .cout(t_1112));
compressor_4_2 u2_387(.a(s_76_22), .b(s_76_21), .c(s_76_20), .d(s_76_19), .cin(s_76_18), .o(t_1113), .co(t_1114), .cout(t_1115));
compressor_3_2 u1_388(.a(s_76_25), .b(s_76_24), .cin(s_76_23), .o(t_1116), .cout(t_1117));
compressor_4_2 u2_389(.a(s_77_2), .b(s_77_1), .c(s_77_0), .d(t_1100), .cin(t_1103), .o(t_1118), .co(t_1119), .cout(t_1120));
compressor_4_2 u2_390(.a(s_77_5), .b(s_77_4), .c(s_77_3), .d(t_1106), .cin(t_1109), .o(t_1121), .co(t_1122), .cout(t_1123));
compressor_4_2 u2_391(.a(s_77_8), .b(s_77_7), .c(s_77_6), .d(t_1112), .cin(t_1115), .o(t_1124), .co(t_1125), .cout(t_1126));
compressor_4_2 u2_392(.a(s_77_12), .b(s_77_11), .c(s_77_10), .d(s_77_9), .cin(t_1117), .o(t_1127), .co(t_1128), .cout(t_1129));
compressor_4_2 u2_393(.a(s_77_17), .b(s_77_16), .c(s_77_15), .d(s_77_14), .cin(s_77_13), .o(t_1130), .co(t_1131), .cout(t_1132));
compressor_4_2 u2_394(.a(s_77_22), .b(s_77_21), .c(s_77_20), .d(s_77_19), .cin(s_77_18), .o(t_1133), .co(t_1134), .cout(t_1135));
compressor_3_2 u1_395(.a(s_77_25), .b(s_77_24), .cin(s_77_23), .o(t_1136), .cout(t_1137));
compressor_4_2 u2_396(.a(s_78_2), .b(s_78_1), .c(s_78_0), .d(t_1120), .cin(t_1123), .o(t_1138), .co(t_1139), .cout(t_1140));
compressor_4_2 u2_397(.a(s_78_5), .b(s_78_4), .c(s_78_3), .d(t_1126), .cin(t_1129), .o(t_1141), .co(t_1142), .cout(t_1143));
compressor_4_2 u2_398(.a(s_78_8), .b(s_78_7), .c(s_78_6), .d(t_1132), .cin(t_1135), .o(t_1144), .co(t_1145), .cout(t_1146));
compressor_4_2 u2_399(.a(s_78_12), .b(s_78_11), .c(s_78_10), .d(s_78_9), .cin(t_1137), .o(t_1147), .co(t_1148), .cout(t_1149));
compressor_4_2 u2_400(.a(s_78_17), .b(s_78_16), .c(s_78_15), .d(s_78_14), .cin(s_78_13), .o(t_1150), .co(t_1151), .cout(t_1152));
compressor_4_2 u2_401(.a(s_78_22), .b(s_78_21), .c(s_78_20), .d(s_78_19), .cin(s_78_18), .o(t_1153), .co(t_1154), .cout(t_1155));
compressor_3_2 u1_402(.a(s_78_25), .b(s_78_24), .cin(s_78_23), .o(t_1156), .cout(t_1157));
compressor_4_2 u2_403(.a(s_79_2), .b(s_79_1), .c(s_79_0), .d(t_1140), .cin(t_1143), .o(t_1158), .co(t_1159), .cout(t_1160));
compressor_4_2 u2_404(.a(s_79_5), .b(s_79_4), .c(s_79_3), .d(t_1146), .cin(t_1149), .o(t_1161), .co(t_1162), .cout(t_1163));
compressor_4_2 u2_405(.a(s_79_8), .b(s_79_7), .c(s_79_6), .d(t_1152), .cin(t_1155), .o(t_1164), .co(t_1165), .cout(t_1166));
compressor_4_2 u2_406(.a(s_79_12), .b(s_79_11), .c(s_79_10), .d(s_79_9), .cin(t_1157), .o(t_1167), .co(t_1168), .cout(t_1169));
compressor_4_2 u2_407(.a(s_79_17), .b(s_79_16), .c(s_79_15), .d(s_79_14), .cin(s_79_13), .o(t_1170), .co(t_1171), .cout(t_1172));
compressor_4_2 u2_408(.a(s_79_22), .b(s_79_21), .c(s_79_20), .d(s_79_19), .cin(s_79_18), .o(t_1173), .co(t_1174), .cout(t_1175));
compressor_3_2 u1_409(.a(s_79_25), .b(s_79_24), .cin(s_79_23), .o(t_1176), .cout(t_1177));
compressor_4_2 u2_410(.a(s_80_2), .b(s_80_1), .c(s_80_0), .d(t_1160), .cin(t_1163), .o(t_1178), .co(t_1179), .cout(t_1180));
compressor_4_2 u2_411(.a(s_80_5), .b(s_80_4), .c(s_80_3), .d(t_1166), .cin(t_1169), .o(t_1181), .co(t_1182), .cout(t_1183));
compressor_4_2 u2_412(.a(s_80_8), .b(s_80_7), .c(s_80_6), .d(t_1172), .cin(t_1175), .o(t_1184), .co(t_1185), .cout(t_1186));
compressor_4_2 u2_413(.a(s_80_12), .b(s_80_11), .c(s_80_10), .d(s_80_9), .cin(t_1177), .o(t_1187), .co(t_1188), .cout(t_1189));
compressor_4_2 u2_414(.a(s_80_17), .b(s_80_16), .c(s_80_15), .d(s_80_14), .cin(s_80_13), .o(t_1190), .co(t_1191), .cout(t_1192));
compressor_4_2 u2_415(.a(s_80_22), .b(s_80_21), .c(s_80_20), .d(s_80_19), .cin(s_80_18), .o(t_1193), .co(t_1194), .cout(t_1195));
half_adder u0_416(.a(s_80_24), .b(s_80_23), .o(t_1196), .cout(t_1197));
compressor_4_2 u2_417(.a(s_81_2), .b(s_81_1), .c(s_81_0), .d(t_1180), .cin(t_1183), .o(t_1198), .co(t_1199), .cout(t_1200));
compressor_4_2 u2_418(.a(s_81_5), .b(s_81_4), .c(s_81_3), .d(t_1186), .cin(t_1189), .o(t_1201), .co(t_1202), .cout(t_1203));
compressor_4_2 u2_419(.a(s_81_8), .b(s_81_7), .c(s_81_6), .d(t_1192), .cin(t_1195), .o(t_1204), .co(t_1205), .cout(t_1206));
compressor_4_2 u2_420(.a(s_81_12), .b(s_81_11), .c(s_81_10), .d(s_81_9), .cin(t_1197), .o(t_1207), .co(t_1208), .cout(t_1209));
compressor_4_2 u2_421(.a(s_81_17), .b(s_81_16), .c(s_81_15), .d(s_81_14), .cin(s_81_13), .o(t_1210), .co(t_1211), .cout(t_1212));
compressor_4_2 u2_422(.a(s_81_22), .b(s_81_21), .c(s_81_20), .d(s_81_19), .cin(s_81_18), .o(t_1213), .co(t_1214), .cout(t_1215));
half_adder u0_423(.a(s_81_24), .b(s_81_23), .o(t_1216), .cout(t_1217));
compressor_4_2 u2_424(.a(s_82_2), .b(s_82_1), .c(s_82_0), .d(t_1200), .cin(t_1203), .o(t_1218), .co(t_1219), .cout(t_1220));
compressor_4_2 u2_425(.a(s_82_5), .b(s_82_4), .c(s_82_3), .d(t_1206), .cin(t_1209), .o(t_1221), .co(t_1222), .cout(t_1223));
compressor_4_2 u2_426(.a(s_82_8), .b(s_82_7), .c(s_82_6), .d(t_1212), .cin(t_1215), .o(t_1224), .co(t_1225), .cout(t_1226));
compressor_4_2 u2_427(.a(s_82_12), .b(s_82_11), .c(s_82_10), .d(s_82_9), .cin(t_1217), .o(t_1227), .co(t_1228), .cout(t_1229));
compressor_4_2 u2_428(.a(s_82_17), .b(s_82_16), .c(s_82_15), .d(s_82_14), .cin(s_82_13), .o(t_1230), .co(t_1231), .cout(t_1232));
compressor_4_2 u2_429(.a(s_82_22), .b(s_82_21), .c(s_82_20), .d(s_82_19), .cin(s_82_18), .o(t_1233), .co(t_1234), .cout(t_1235));
compressor_4_2 u2_430(.a(s_83_2), .b(s_83_1), .c(s_83_0), .d(t_1220), .cin(t_1223), .o(t_1236), .co(t_1237), .cout(t_1238));
compressor_4_2 u2_431(.a(s_83_5), .b(s_83_4), .c(s_83_3), .d(t_1226), .cin(t_1229), .o(t_1239), .co(t_1240), .cout(t_1241));
compressor_4_2 u2_432(.a(s_83_8), .b(s_83_7), .c(s_83_6), .d(t_1232), .cin(t_1235), .o(t_1242), .co(t_1243), .cout(t_1244));
compressor_4_2 u2_433(.a(s_83_13), .b(s_83_12), .c(s_83_11), .d(s_83_10), .cin(s_83_9), .o(t_1245), .co(t_1246), .cout(t_1247));
compressor_4_2 u2_434(.a(s_83_18), .b(s_83_17), .c(s_83_16), .d(s_83_15), .cin(s_83_14), .o(t_1248), .co(t_1249), .cout(t_1250));
compressor_4_2 u2_435(.a(s_83_23), .b(s_83_22), .c(s_83_21), .d(s_83_20), .cin(s_83_19), .o(t_1251), .co(t_1252), .cout(t_1253));
compressor_4_2 u2_436(.a(s_84_2), .b(s_84_1), .c(s_84_0), .d(t_1238), .cin(t_1241), .o(t_1254), .co(t_1255), .cout(t_1256));
compressor_4_2 u2_437(.a(s_84_5), .b(s_84_4), .c(s_84_3), .d(t_1244), .cin(t_1247), .o(t_1257), .co(t_1258), .cout(t_1259));
compressor_4_2 u2_438(.a(s_84_8), .b(s_84_7), .c(s_84_6), .d(t_1250), .cin(t_1253), .o(t_1260), .co(t_1261), .cout(t_1262));
compressor_4_2 u2_439(.a(s_84_13), .b(s_84_12), .c(s_84_11), .d(s_84_10), .cin(s_84_9), .o(t_1263), .co(t_1264), .cout(t_1265));
compressor_4_2 u2_440(.a(s_84_18), .b(s_84_17), .c(s_84_16), .d(s_84_15), .cin(s_84_14), .o(t_1266), .co(t_1267), .cout(t_1268));
compressor_3_2 u1_441(.a(s_84_21), .b(s_84_20), .cin(s_84_19), .o(t_1269), .cout(t_1270));
compressor_4_2 u2_442(.a(s_85_2), .b(s_85_1), .c(s_85_0), .d(t_1256), .cin(t_1259), .o(t_1271), .co(t_1272), .cout(t_1273));
compressor_4_2 u2_443(.a(s_85_5), .b(s_85_4), .c(s_85_3), .d(t_1262), .cin(t_1265), .o(t_1274), .co(t_1275), .cout(t_1276));
compressor_4_2 u2_444(.a(s_85_8), .b(s_85_7), .c(s_85_6), .d(t_1268), .cin(t_1270), .o(t_1277), .co(t_1278), .cout(t_1279));
compressor_4_2 u2_445(.a(s_85_13), .b(s_85_12), .c(s_85_11), .d(s_85_10), .cin(s_85_9), .o(t_1280), .co(t_1281), .cout(t_1282));
compressor_4_2 u2_446(.a(s_85_18), .b(s_85_17), .c(s_85_16), .d(s_85_15), .cin(s_85_14), .o(t_1283), .co(t_1284), .cout(t_1285));
compressor_3_2 u1_447(.a(s_85_21), .b(s_85_20), .cin(s_85_19), .o(t_1286), .cout(t_1287));
compressor_4_2 u2_448(.a(s_86_2), .b(s_86_1), .c(s_86_0), .d(t_1273), .cin(t_1276), .o(t_1288), .co(t_1289), .cout(t_1290));
compressor_4_2 u2_449(.a(s_86_5), .b(s_86_4), .c(s_86_3), .d(t_1279), .cin(t_1282), .o(t_1291), .co(t_1292), .cout(t_1293));
compressor_4_2 u2_450(.a(s_86_8), .b(s_86_7), .c(s_86_6), .d(t_1285), .cin(t_1287), .o(t_1294), .co(t_1295), .cout(t_1296));
compressor_4_2 u2_451(.a(s_86_13), .b(s_86_12), .c(s_86_11), .d(s_86_10), .cin(s_86_9), .o(t_1297), .co(t_1298), .cout(t_1299));
compressor_4_2 u2_452(.a(s_86_18), .b(s_86_17), .c(s_86_16), .d(s_86_15), .cin(s_86_14), .o(t_1300), .co(t_1301), .cout(t_1302));
compressor_3_2 u1_453(.a(s_86_21), .b(s_86_20), .cin(s_86_19), .o(t_1303), .cout(t_1304));
compressor_4_2 u2_454(.a(s_87_2), .b(s_87_1), .c(s_87_0), .d(t_1290), .cin(t_1293), .o(t_1305), .co(t_1306), .cout(t_1307));
compressor_4_2 u2_455(.a(s_87_5), .b(s_87_4), .c(s_87_3), .d(t_1296), .cin(t_1299), .o(t_1308), .co(t_1309), .cout(t_1310));
compressor_4_2 u2_456(.a(s_87_8), .b(s_87_7), .c(s_87_6), .d(t_1302), .cin(t_1304), .o(t_1311), .co(t_1312), .cout(t_1313));
compressor_4_2 u2_457(.a(s_87_13), .b(s_87_12), .c(s_87_11), .d(s_87_10), .cin(s_87_9), .o(t_1314), .co(t_1315), .cout(t_1316));
compressor_4_2 u2_458(.a(s_87_18), .b(s_87_17), .c(s_87_16), .d(s_87_15), .cin(s_87_14), .o(t_1317), .co(t_1318), .cout(t_1319));
compressor_3_2 u1_459(.a(s_87_21), .b(s_87_20), .cin(s_87_19), .o(t_1320), .cout(t_1321));
compressor_4_2 u2_460(.a(s_88_2), .b(s_88_1), .c(s_88_0), .d(t_1307), .cin(t_1310), .o(t_1322), .co(t_1323), .cout(t_1324));
compressor_4_2 u2_461(.a(s_88_5), .b(s_88_4), .c(s_88_3), .d(t_1313), .cin(t_1316), .o(t_1325), .co(t_1326), .cout(t_1327));
compressor_4_2 u2_462(.a(s_88_8), .b(s_88_7), .c(s_88_6), .d(t_1319), .cin(t_1321), .o(t_1328), .co(t_1329), .cout(t_1330));
compressor_4_2 u2_463(.a(s_88_13), .b(s_88_12), .c(s_88_11), .d(s_88_10), .cin(s_88_9), .o(t_1331), .co(t_1332), .cout(t_1333));
compressor_4_2 u2_464(.a(s_88_18), .b(s_88_17), .c(s_88_16), .d(s_88_15), .cin(s_88_14), .o(t_1334), .co(t_1335), .cout(t_1336));
half_adder u0_465(.a(s_88_20), .b(s_88_19), .o(t_1337), .cout(t_1338));
compressor_4_2 u2_466(.a(s_89_2), .b(s_89_1), .c(s_89_0), .d(t_1324), .cin(t_1327), .o(t_1339), .co(t_1340), .cout(t_1341));
compressor_4_2 u2_467(.a(s_89_5), .b(s_89_4), .c(s_89_3), .d(t_1330), .cin(t_1333), .o(t_1342), .co(t_1343), .cout(t_1344));
compressor_4_2 u2_468(.a(s_89_8), .b(s_89_7), .c(s_89_6), .d(t_1336), .cin(t_1338), .o(t_1345), .co(t_1346), .cout(t_1347));
compressor_4_2 u2_469(.a(s_89_13), .b(s_89_12), .c(s_89_11), .d(s_89_10), .cin(s_89_9), .o(t_1348), .co(t_1349), .cout(t_1350));
compressor_4_2 u2_470(.a(s_89_18), .b(s_89_17), .c(s_89_16), .d(s_89_15), .cin(s_89_14), .o(t_1351), .co(t_1352), .cout(t_1353));
half_adder u0_471(.a(s_89_20), .b(s_89_19), .o(t_1354), .cout(t_1355));
compressor_4_2 u2_472(.a(s_90_2), .b(s_90_1), .c(s_90_0), .d(t_1341), .cin(t_1344), .o(t_1356), .co(t_1357), .cout(t_1358));
compressor_4_2 u2_473(.a(s_90_5), .b(s_90_4), .c(s_90_3), .d(t_1347), .cin(t_1350), .o(t_1359), .co(t_1360), .cout(t_1361));
compressor_4_2 u2_474(.a(s_90_8), .b(s_90_7), .c(s_90_6), .d(t_1353), .cin(t_1355), .o(t_1362), .co(t_1363), .cout(t_1364));
compressor_4_2 u2_475(.a(s_90_13), .b(s_90_12), .c(s_90_11), .d(s_90_10), .cin(s_90_9), .o(t_1365), .co(t_1366), .cout(t_1367));
compressor_4_2 u2_476(.a(s_90_18), .b(s_90_17), .c(s_90_16), .d(s_90_15), .cin(s_90_14), .o(t_1368), .co(t_1369), .cout(t_1370));
compressor_4_2 u2_477(.a(s_91_2), .b(s_91_1), .c(s_91_0), .d(t_1358), .cin(t_1361), .o(t_1371), .co(t_1372), .cout(t_1373));
compressor_4_2 u2_478(.a(s_91_5), .b(s_91_4), .c(s_91_3), .d(t_1364), .cin(t_1367), .o(t_1374), .co(t_1375), .cout(t_1376));
compressor_4_2 u2_479(.a(s_91_9), .b(s_91_8), .c(s_91_7), .d(s_91_6), .cin(t_1370), .o(t_1377), .co(t_1378), .cout(t_1379));
compressor_4_2 u2_480(.a(s_91_14), .b(s_91_13), .c(s_91_12), .d(s_91_11), .cin(s_91_10), .o(t_1380), .co(t_1381), .cout(t_1382));
compressor_4_2 u2_481(.a(s_91_19), .b(s_91_18), .c(s_91_17), .d(s_91_16), .cin(s_91_15), .o(t_1383), .co(t_1384), .cout(t_1385));
compressor_4_2 u2_482(.a(s_92_2), .b(s_92_1), .c(s_92_0), .d(t_1373), .cin(t_1376), .o(t_1386), .co(t_1387), .cout(t_1388));
compressor_4_2 u2_483(.a(s_92_5), .b(s_92_4), .c(s_92_3), .d(t_1379), .cin(t_1382), .o(t_1389), .co(t_1390), .cout(t_1391));
compressor_4_2 u2_484(.a(s_92_9), .b(s_92_8), .c(s_92_7), .d(s_92_6), .cin(t_1385), .o(t_1392), .co(t_1393), .cout(t_1394));
compressor_4_2 u2_485(.a(s_92_14), .b(s_92_13), .c(s_92_12), .d(s_92_11), .cin(s_92_10), .o(t_1395), .co(t_1396), .cout(t_1397));
compressor_3_2 u1_486(.a(s_92_17), .b(s_92_16), .cin(s_92_15), .o(t_1398), .cout(t_1399));
compressor_4_2 u2_487(.a(s_93_2), .b(s_93_1), .c(s_93_0), .d(t_1388), .cin(t_1391), .o(t_1400), .co(t_1401), .cout(t_1402));
compressor_4_2 u2_488(.a(s_93_5), .b(s_93_4), .c(s_93_3), .d(t_1394), .cin(t_1397), .o(t_1403), .co(t_1404), .cout(t_1405));
compressor_4_2 u2_489(.a(s_93_9), .b(s_93_8), .c(s_93_7), .d(s_93_6), .cin(t_1399), .o(t_1406), .co(t_1407), .cout(t_1408));
compressor_4_2 u2_490(.a(s_93_14), .b(s_93_13), .c(s_93_12), .d(s_93_11), .cin(s_93_10), .o(t_1409), .co(t_1410), .cout(t_1411));
compressor_3_2 u1_491(.a(s_93_17), .b(s_93_16), .cin(s_93_15), .o(t_1412), .cout(t_1413));
compressor_4_2 u2_492(.a(s_94_2), .b(s_94_1), .c(s_94_0), .d(t_1402), .cin(t_1405), .o(t_1414), .co(t_1415), .cout(t_1416));
compressor_4_2 u2_493(.a(s_94_5), .b(s_94_4), .c(s_94_3), .d(t_1408), .cin(t_1411), .o(t_1417), .co(t_1418), .cout(t_1419));
compressor_4_2 u2_494(.a(s_94_9), .b(s_94_8), .c(s_94_7), .d(s_94_6), .cin(t_1413), .o(t_1420), .co(t_1421), .cout(t_1422));
compressor_4_2 u2_495(.a(s_94_14), .b(s_94_13), .c(s_94_12), .d(s_94_11), .cin(s_94_10), .o(t_1423), .co(t_1424), .cout(t_1425));
compressor_3_2 u1_496(.a(s_94_17), .b(s_94_16), .cin(s_94_15), .o(t_1426), .cout(t_1427));
compressor_4_2 u2_497(.a(s_95_2), .b(s_95_1), .c(s_95_0), .d(t_1416), .cin(t_1419), .o(t_1428), .co(t_1429), .cout(t_1430));
compressor_4_2 u2_498(.a(s_95_5), .b(s_95_4), .c(s_95_3), .d(t_1422), .cin(t_1425), .o(t_1431), .co(t_1432), .cout(t_1433));
compressor_4_2 u2_499(.a(s_95_9), .b(s_95_8), .c(s_95_7), .d(s_95_6), .cin(t_1427), .o(t_1434), .co(t_1435), .cout(t_1436));
compressor_4_2 u2_500(.a(s_95_14), .b(s_95_13), .c(s_95_12), .d(s_95_11), .cin(s_95_10), .o(t_1437), .co(t_1438), .cout(t_1439));
compressor_3_2 u1_501(.a(s_95_17), .b(s_95_16), .cin(s_95_15), .o(t_1440), .cout(t_1441));
compressor_4_2 u2_502(.a(s_96_2), .b(s_96_1), .c(s_96_0), .d(t_1430), .cin(t_1433), .o(t_1442), .co(t_1443), .cout(t_1444));
compressor_4_2 u2_503(.a(s_96_5), .b(s_96_4), .c(s_96_3), .d(t_1436), .cin(t_1439), .o(t_1445), .co(t_1446), .cout(t_1447));
compressor_4_2 u2_504(.a(s_96_9), .b(s_96_8), .c(s_96_7), .d(s_96_6), .cin(t_1441), .o(t_1448), .co(t_1449), .cout(t_1450));
compressor_4_2 u2_505(.a(s_96_14), .b(s_96_13), .c(s_96_12), .d(s_96_11), .cin(s_96_10), .o(t_1451), .co(t_1452), .cout(t_1453));
half_adder u0_506(.a(s_96_16), .b(s_96_15), .o(t_1454), .cout(t_1455));
compressor_4_2 u2_507(.a(s_97_2), .b(s_97_1), .c(s_97_0), .d(t_1444), .cin(t_1447), .o(t_1456), .co(t_1457), .cout(t_1458));
compressor_4_2 u2_508(.a(s_97_5), .b(s_97_4), .c(s_97_3), .d(t_1450), .cin(t_1453), .o(t_1459), .co(t_1460), .cout(t_1461));
compressor_4_2 u2_509(.a(s_97_9), .b(s_97_8), .c(s_97_7), .d(s_97_6), .cin(t_1455), .o(t_1462), .co(t_1463), .cout(t_1464));
compressor_4_2 u2_510(.a(s_97_14), .b(s_97_13), .c(s_97_12), .d(s_97_11), .cin(s_97_10), .o(t_1465), .co(t_1466), .cout(t_1467));
half_adder u0_511(.a(s_97_16), .b(s_97_15), .o(t_1468), .cout(t_1469));
compressor_4_2 u2_512(.a(s_98_2), .b(s_98_1), .c(s_98_0), .d(t_1458), .cin(t_1461), .o(t_1470), .co(t_1471), .cout(t_1472));
compressor_4_2 u2_513(.a(s_98_5), .b(s_98_4), .c(s_98_3), .d(t_1464), .cin(t_1467), .o(t_1473), .co(t_1474), .cout(t_1475));
compressor_4_2 u2_514(.a(s_98_9), .b(s_98_8), .c(s_98_7), .d(s_98_6), .cin(t_1469), .o(t_1476), .co(t_1477), .cout(t_1478));
compressor_4_2 u2_515(.a(s_98_14), .b(s_98_13), .c(s_98_12), .d(s_98_11), .cin(s_98_10), .o(t_1479), .co(t_1480), .cout(t_1481));
compressor_4_2 u2_516(.a(s_99_2), .b(s_99_1), .c(s_99_0), .d(t_1472), .cin(t_1475), .o(t_1482), .co(t_1483), .cout(t_1484));
compressor_4_2 u2_517(.a(s_99_5), .b(s_99_4), .c(s_99_3), .d(t_1478), .cin(t_1481), .o(t_1485), .co(t_1486), .cout(t_1487));
compressor_4_2 u2_518(.a(s_99_10), .b(s_99_9), .c(s_99_8), .d(s_99_7), .cin(s_99_6), .o(t_1488), .co(t_1489), .cout(t_1490));
compressor_4_2 u2_519(.a(s_99_15), .b(s_99_14), .c(s_99_13), .d(s_99_12), .cin(s_99_11), .o(t_1491), .co(t_1492), .cout(t_1493));
compressor_4_2 u2_520(.a(s_100_2), .b(s_100_1), .c(s_100_0), .d(t_1484), .cin(t_1487), .o(t_1494), .co(t_1495), .cout(t_1496));
compressor_4_2 u2_521(.a(s_100_5), .b(s_100_4), .c(s_100_3), .d(t_1490), .cin(t_1493), .o(t_1497), .co(t_1498), .cout(t_1499));
compressor_4_2 u2_522(.a(s_100_10), .b(s_100_9), .c(s_100_8), .d(s_100_7), .cin(s_100_6), .o(t_1500), .co(t_1501), .cout(t_1502));
compressor_3_2 u1_523(.a(s_100_13), .b(s_100_12), .cin(s_100_11), .o(t_1503), .cout(t_1504));
compressor_4_2 u2_524(.a(s_101_2), .b(s_101_1), .c(s_101_0), .d(t_1496), .cin(t_1499), .o(t_1505), .co(t_1506), .cout(t_1507));
compressor_4_2 u2_525(.a(s_101_5), .b(s_101_4), .c(s_101_3), .d(t_1502), .cin(t_1504), .o(t_1508), .co(t_1509), .cout(t_1510));
compressor_4_2 u2_526(.a(s_101_10), .b(s_101_9), .c(s_101_8), .d(s_101_7), .cin(s_101_6), .o(t_1511), .co(t_1512), .cout(t_1513));
compressor_3_2 u1_527(.a(s_101_13), .b(s_101_12), .cin(s_101_11), .o(t_1514), .cout(t_1515));
compressor_4_2 u2_528(.a(s_102_2), .b(s_102_1), .c(s_102_0), .d(t_1507), .cin(t_1510), .o(t_1516), .co(t_1517), .cout(t_1518));
compressor_4_2 u2_529(.a(s_102_5), .b(s_102_4), .c(s_102_3), .d(t_1513), .cin(t_1515), .o(t_1519), .co(t_1520), .cout(t_1521));
compressor_4_2 u2_530(.a(s_102_10), .b(s_102_9), .c(s_102_8), .d(s_102_7), .cin(s_102_6), .o(t_1522), .co(t_1523), .cout(t_1524));
compressor_3_2 u1_531(.a(s_102_13), .b(s_102_12), .cin(s_102_11), .o(t_1525), .cout(t_1526));
compressor_4_2 u2_532(.a(s_103_2), .b(s_103_1), .c(s_103_0), .d(t_1518), .cin(t_1521), .o(t_1527), .co(t_1528), .cout(t_1529));
compressor_4_2 u2_533(.a(s_103_5), .b(s_103_4), .c(s_103_3), .d(t_1524), .cin(t_1526), .o(t_1530), .co(t_1531), .cout(t_1532));
compressor_4_2 u2_534(.a(s_103_10), .b(s_103_9), .c(s_103_8), .d(s_103_7), .cin(s_103_6), .o(t_1533), .co(t_1534), .cout(t_1535));
compressor_3_2 u1_535(.a(s_103_13), .b(s_103_12), .cin(s_103_11), .o(t_1536), .cout(t_1537));
compressor_4_2 u2_536(.a(s_104_2), .b(s_104_1), .c(s_104_0), .d(t_1529), .cin(t_1532), .o(t_1538), .co(t_1539), .cout(t_1540));
compressor_4_2 u2_537(.a(s_104_5), .b(s_104_4), .c(s_104_3), .d(t_1535), .cin(t_1537), .o(t_1541), .co(t_1542), .cout(t_1543));
compressor_4_2 u2_538(.a(s_104_10), .b(s_104_9), .c(s_104_8), .d(s_104_7), .cin(s_104_6), .o(t_1544), .co(t_1545), .cout(t_1546));
half_adder u0_539(.a(s_104_12), .b(s_104_11), .o(t_1547), .cout(t_1548));
compressor_4_2 u2_540(.a(s_105_2), .b(s_105_1), .c(s_105_0), .d(t_1540), .cin(t_1543), .o(t_1549), .co(t_1550), .cout(t_1551));
compressor_4_2 u2_541(.a(s_105_5), .b(s_105_4), .c(s_105_3), .d(t_1546), .cin(t_1548), .o(t_1552), .co(t_1553), .cout(t_1554));
compressor_4_2 u2_542(.a(s_105_10), .b(s_105_9), .c(s_105_8), .d(s_105_7), .cin(s_105_6), .o(t_1555), .co(t_1556), .cout(t_1557));
half_adder u0_543(.a(s_105_12), .b(s_105_11), .o(t_1558), .cout(t_1559));
compressor_4_2 u2_544(.a(s_106_2), .b(s_106_1), .c(s_106_0), .d(t_1551), .cin(t_1554), .o(t_1560), .co(t_1561), .cout(t_1562));
compressor_4_2 u2_545(.a(s_106_5), .b(s_106_4), .c(s_106_3), .d(t_1557), .cin(t_1559), .o(t_1563), .co(t_1564), .cout(t_1565));
compressor_4_2 u2_546(.a(s_106_10), .b(s_106_9), .c(s_106_8), .d(s_106_7), .cin(s_106_6), .o(t_1566), .co(t_1567), .cout(t_1568));
compressor_4_2 u2_547(.a(s_107_2), .b(s_107_1), .c(s_107_0), .d(t_1562), .cin(t_1565), .o(t_1569), .co(t_1570), .cout(t_1571));
compressor_4_2 u2_548(.a(s_107_6), .b(s_107_5), .c(s_107_4), .d(s_107_3), .cin(t_1568), .o(t_1572), .co(t_1573), .cout(t_1574));
compressor_4_2 u2_549(.a(s_107_11), .b(s_107_10), .c(s_107_9), .d(s_107_8), .cin(s_107_7), .o(t_1575), .co(t_1576), .cout(t_1577));
compressor_4_2 u2_550(.a(s_108_2), .b(s_108_1), .c(s_108_0), .d(t_1571), .cin(t_1574), .o(t_1578), .co(t_1579), .cout(t_1580));
compressor_4_2 u2_551(.a(s_108_6), .b(s_108_5), .c(s_108_4), .d(s_108_3), .cin(t_1577), .o(t_1581), .co(t_1582), .cout(t_1583));
compressor_3_2 u1_552(.a(s_108_9), .b(s_108_8), .cin(s_108_7), .o(t_1584), .cout(t_1585));
compressor_4_2 u2_553(.a(s_109_2), .b(s_109_1), .c(s_109_0), .d(t_1580), .cin(t_1583), .o(t_1586), .co(t_1587), .cout(t_1588));
compressor_4_2 u2_554(.a(s_109_6), .b(s_109_5), .c(s_109_4), .d(s_109_3), .cin(t_1585), .o(t_1589), .co(t_1590), .cout(t_1591));
compressor_3_2 u1_555(.a(s_109_9), .b(s_109_8), .cin(s_109_7), .o(t_1592), .cout(t_1593));
compressor_4_2 u2_556(.a(s_110_2), .b(s_110_1), .c(s_110_0), .d(t_1588), .cin(t_1591), .o(t_1594), .co(t_1595), .cout(t_1596));
compressor_4_2 u2_557(.a(s_110_6), .b(s_110_5), .c(s_110_4), .d(s_110_3), .cin(t_1593), .o(t_1597), .co(t_1598), .cout(t_1599));
compressor_3_2 u1_558(.a(s_110_9), .b(s_110_8), .cin(s_110_7), .o(t_1600), .cout(t_1601));
compressor_4_2 u2_559(.a(s_111_2), .b(s_111_1), .c(s_111_0), .d(t_1596), .cin(t_1599), .o(t_1602), .co(t_1603), .cout(t_1604));
compressor_4_2 u2_560(.a(s_111_6), .b(s_111_5), .c(s_111_4), .d(s_111_3), .cin(t_1601), .o(t_1605), .co(t_1606), .cout(t_1607));
compressor_3_2 u1_561(.a(s_111_9), .b(s_111_8), .cin(s_111_7), .o(t_1608), .cout(t_1609));
compressor_4_2 u2_562(.a(s_112_2), .b(s_112_1), .c(s_112_0), .d(t_1604), .cin(t_1607), .o(t_1610), .co(t_1611), .cout(t_1612));
compressor_4_2 u2_563(.a(s_112_6), .b(s_112_5), .c(s_112_4), .d(s_112_3), .cin(t_1609), .o(t_1613), .co(t_1614), .cout(t_1615));
half_adder u0_564(.a(s_112_8), .b(s_112_7), .o(t_1616), .cout(t_1617));
compressor_4_2 u2_565(.a(s_113_2), .b(s_113_1), .c(s_113_0), .d(t_1612), .cin(t_1615), .o(t_1618), .co(t_1619), .cout(t_1620));
compressor_4_2 u2_566(.a(s_113_6), .b(s_113_5), .c(s_113_4), .d(s_113_3), .cin(t_1617), .o(t_1621), .co(t_1622), .cout(t_1623));
half_adder u0_567(.a(s_113_8), .b(s_113_7), .o(t_1624), .cout(t_1625));
compressor_4_2 u2_568(.a(s_114_2), .b(s_114_1), .c(s_114_0), .d(t_1620), .cin(t_1623), .o(t_1626), .co(t_1627), .cout(t_1628));
compressor_4_2 u2_569(.a(s_114_6), .b(s_114_5), .c(s_114_4), .d(s_114_3), .cin(t_1625), .o(t_1629), .co(t_1630), .cout(t_1631));
compressor_4_2 u2_570(.a(s_115_2), .b(s_115_1), .c(s_115_0), .d(t_1628), .cin(t_1631), .o(t_1632), .co(t_1633), .cout(t_1634));
compressor_4_2 u2_571(.a(s_115_7), .b(s_115_6), .c(s_115_5), .d(s_115_4), .cin(s_115_3), .o(t_1635), .co(t_1636), .cout(t_1637));
compressor_4_2 u2_572(.a(s_116_2), .b(s_116_1), .c(s_116_0), .d(t_1634), .cin(t_1637), .o(t_1638), .co(t_1639), .cout(t_1640));
compressor_3_2 u1_573(.a(s_116_5), .b(s_116_4), .cin(s_116_3), .o(t_1641), .cout(t_1642));
compressor_4_2 u2_574(.a(s_117_2), .b(s_117_1), .c(s_117_0), .d(t_1640), .cin(t_1642), .o(t_1643), .co(t_1644), .cout(t_1645));
compressor_3_2 u1_575(.a(s_117_5), .b(s_117_4), .cin(s_117_3), .o(t_1646), .cout(t_1647));
compressor_4_2 u2_576(.a(s_118_2), .b(s_118_1), .c(s_118_0), .d(t_1645), .cin(t_1647), .o(t_1648), .co(t_1649), .cout(t_1650));
compressor_3_2 u1_577(.a(s_118_5), .b(s_118_4), .cin(s_118_3), .o(t_1651), .cout(t_1652));
compressor_4_2 u2_578(.a(s_119_2), .b(s_119_1), .c(s_119_0), .d(t_1650), .cin(t_1652), .o(t_1653), .co(t_1654), .cout(t_1655));
compressor_3_2 u1_579(.a(s_119_5), .b(s_119_4), .cin(s_119_3), .o(t_1656), .cout(t_1657));
compressor_4_2 u2_580(.a(s_120_2), .b(s_120_1), .c(s_120_0), .d(t_1655), .cin(t_1657), .o(t_1658), .co(t_1659), .cout(t_1660));
half_adder u0_581(.a(s_120_4), .b(s_120_3), .o(t_1661), .cout(t_1662));
compressor_4_2 u2_582(.a(s_121_2), .b(s_121_1), .c(s_121_0), .d(t_1660), .cin(t_1662), .o(t_1663), .co(t_1664), .cout(t_1665));
half_adder u0_583(.a(s_121_4), .b(s_121_3), .o(t_1666), .cout(t_1667));
compressor_4_2 u2_584(.a(s_122_2), .b(s_122_1), .c(s_122_0), .d(t_1665), .cin(t_1667), .o(t_1668), .co(t_1669), .cout(t_1670));
compressor_4_2 u2_585(.a(s_123_3), .b(s_123_2), .c(s_123_1), .d(s_123_0), .cin(t_1670), .o(t_1671), .co(t_1672), .cout(t_1673));
compressor_3_2 u1_586(.a(s_124_1), .b(s_124_0), .cin(t_1673), .o(t_1674), .cout(t_1675));
compressor_3_2 u1_587(.a(s_125_2), .b(s_125_1), .cin(s_125_0), .o(t_1676), .cout(t_1677));
half_adder u0_588(.a(s_126_1), .b(s_126_0), .o(t_1678), .cout(t_1679));
half_adder u0_589(.a(s_127_1), .b(s_127_0), .o(t_1680), .cout());

/* u0_590 Output nets */
wire t_1681,   t_1682;
/* u0_591 Output nets */
wire t_1683,   t_1684;
/* u1_592 Output nets */
wire t_1685,   t_1686;
/* u0_593 Output nets */
wire t_1687,   t_1688;
/* u0_594 Output nets */
wire t_1689,   t_1690;
/* u1_595 Output nets */
wire t_1691,   t_1692;
/* u1_596 Output nets */
wire t_1693,   t_1694;
/* u2_597 Output nets */
wire t_1695,   t_1696,   t_1697;
/* u1_598 Output nets */
wire t_1698,   t_1699;
/* u1_599 Output nets */
wire t_1700,   t_1701;
/* u2_600 Output nets */
wire t_1702,   t_1703,   t_1704;
/* u2_601 Output nets */
wire t_1705,   t_1706,   t_1707;
/* u2_602 Output nets */
wire t_1708,   t_1709,   t_1710;
/* u2_603 Output nets */
wire t_1711,   t_1712,   t_1713;
/* u2_604 Output nets */
wire t_1714,   t_1715,   t_1716;
/* u2_605 Output nets */
wire t_1717,   t_1718,   t_1719;
/* u0_606 Output nets */
wire t_1720,   t_1721;
/* u2_607 Output nets */
wire t_1722,   t_1723,   t_1724;
/* u0_608 Output nets */
wire t_1725,   t_1726;
/* u2_609 Output nets */
wire t_1727,   t_1728,   t_1729;
/* u0_610 Output nets */
wire t_1730,   t_1731;
/* u2_611 Output nets */
wire t_1732,   t_1733,   t_1734;
/* u1_612 Output nets */
wire t_1735,   t_1736;
/* u2_613 Output nets */
wire t_1737,   t_1738,   t_1739;
/* u1_614 Output nets */
wire t_1740,   t_1741;
/* u2_615 Output nets */
wire t_1742,   t_1743,   t_1744;
/* u1_616 Output nets */
wire t_1745,   t_1746;
/* u2_617 Output nets */
wire t_1747,   t_1748,   t_1749;
/* u1_618 Output nets */
wire t_1750,   t_1751;
/* u2_619 Output nets */
wire t_1752,   t_1753,   t_1754;
/* u1_620 Output nets */
wire t_1755,   t_1756;
/* u2_621 Output nets */
wire t_1757,   t_1758,   t_1759;
/* u2_622 Output nets */
wire t_1760,   t_1761,   t_1762;
/* u2_623 Output nets */
wire t_1763,   t_1764,   t_1765;
/* u1_624 Output nets */
wire t_1766,   t_1767;
/* u2_625 Output nets */
wire t_1768,   t_1769,   t_1770;
/* u1_626 Output nets */
wire t_1771,   t_1772;
/* u2_627 Output nets */
wire t_1773,   t_1774,   t_1775;
/* u2_628 Output nets */
wire t_1776,   t_1777,   t_1778;
/* u2_629 Output nets */
wire t_1779,   t_1780,   t_1781;
/* u2_630 Output nets */
wire t_1782,   t_1783,   t_1784;
/* u2_631 Output nets */
wire t_1785,   t_1786,   t_1787;
/* u2_632 Output nets */
wire t_1788,   t_1789,   t_1790;
/* u2_633 Output nets */
wire t_1791,   t_1792,   t_1793;
/* u2_634 Output nets */
wire t_1794,   t_1795,   t_1796;
/* u2_635 Output nets */
wire t_1797,   t_1798,   t_1799;
/* u2_636 Output nets */
wire t_1800,   t_1801,   t_1802;
/* u2_637 Output nets */
wire t_1803,   t_1804,   t_1805;
/* u2_638 Output nets */
wire t_1806,   t_1807,   t_1808;
/* u0_639 Output nets */
wire t_1809,   t_1810;
/* u2_640 Output nets */
wire t_1811,   t_1812,   t_1813;
/* u2_641 Output nets */
wire t_1814,   t_1815,   t_1816;
/* u0_642 Output nets */
wire t_1817,   t_1818;
/* u2_643 Output nets */
wire t_1819,   t_1820,   t_1821;
/* u2_644 Output nets */
wire t_1822,   t_1823,   t_1824;
/* u0_645 Output nets */
wire t_1825,   t_1826;
/* u2_646 Output nets */
wire t_1827,   t_1828,   t_1829;
/* u2_647 Output nets */
wire t_1830,   t_1831,   t_1832;
/* u1_648 Output nets */
wire t_1833,   t_1834;
/* u2_649 Output nets */
wire t_1835,   t_1836,   t_1837;
/* u2_650 Output nets */
wire t_1838,   t_1839,   t_1840;
/* u1_651 Output nets */
wire t_1841,   t_1842;
/* u2_652 Output nets */
wire t_1843,   t_1844,   t_1845;
/* u2_653 Output nets */
wire t_1846,   t_1847,   t_1848;
/* u1_654 Output nets */
wire t_1849,   t_1850;
/* u2_655 Output nets */
wire t_1851,   t_1852,   t_1853;
/* u2_656 Output nets */
wire t_1854,   t_1855,   t_1856;
/* u1_657 Output nets */
wire t_1857,   t_1858;
/* u2_658 Output nets */
wire t_1859,   t_1860,   t_1861;
/* u2_659 Output nets */
wire t_1862,   t_1863,   t_1864;
/* u1_660 Output nets */
wire t_1865,   t_1866;
/* u2_661 Output nets */
wire t_1867,   t_1868,   t_1869;
/* u2_662 Output nets */
wire t_1870,   t_1871,   t_1872;
/* u2_663 Output nets */
wire t_1873,   t_1874,   t_1875;
/* u2_664 Output nets */
wire t_1876,   t_1877,   t_1878;
/* u2_665 Output nets */
wire t_1879,   t_1880,   t_1881;
/* u1_666 Output nets */
wire t_1882,   t_1883;
/* u2_667 Output nets */
wire t_1884,   t_1885,   t_1886;
/* u2_668 Output nets */
wire t_1887,   t_1888,   t_1889;
/* u1_669 Output nets */
wire t_1890,   t_1891;
/* u2_670 Output nets */
wire t_1892,   t_1893,   t_1894;
/* u2_671 Output nets */
wire t_1895,   t_1896,   t_1897;
/* u2_672 Output nets */
wire t_1898,   t_1899,   t_1900;
/* u2_673 Output nets */
wire t_1901,   t_1902,   t_1903;
/* u2_674 Output nets */
wire t_1904,   t_1905,   t_1906;
/* u2_675 Output nets */
wire t_1907,   t_1908,   t_1909;
/* u2_676 Output nets */
wire t_1910,   t_1911,   t_1912;
/* u2_677 Output nets */
wire t_1913,   t_1914,   t_1915;
/* u2_678 Output nets */
wire t_1916,   t_1917,   t_1918;
/* u2_679 Output nets */
wire t_1919,   t_1920,   t_1921;
/* u2_680 Output nets */
wire t_1922,   t_1923,   t_1924;
/* u2_681 Output nets */
wire t_1925,   t_1926,   t_1927;
/* u2_682 Output nets */
wire t_1928,   t_1929,   t_1930;
/* u2_683 Output nets */
wire t_1931,   t_1932,   t_1933;
/* u2_684 Output nets */
wire t_1934,   t_1935,   t_1936;
/* u2_685 Output nets */
wire t_1937,   t_1938,   t_1939;
/* u2_686 Output nets */
wire t_1940,   t_1941,   t_1942;
/* u2_687 Output nets */
wire t_1943,   t_1944,   t_1945;
/* u0_688 Output nets */
wire t_1946,   t_1947;
/* u2_689 Output nets */
wire t_1948,   t_1949,   t_1950;
/* u2_690 Output nets */
wire t_1951,   t_1952,   t_1953;
/* u2_691 Output nets */
wire t_1954,   t_1955,   t_1956;
/* u0_692 Output nets */
wire t_1957,   t_1958;
/* u2_693 Output nets */
wire t_1959,   t_1960,   t_1961;
/* u2_694 Output nets */
wire t_1962,   t_1963,   t_1964;
/* u2_695 Output nets */
wire t_1965,   t_1966,   t_1967;
/* u0_696 Output nets */
wire t_1968,   t_1969;
/* u2_697 Output nets */
wire t_1970,   t_1971,   t_1972;
/* u2_698 Output nets */
wire t_1973,   t_1974,   t_1975;
/* u2_699 Output nets */
wire t_1976,   t_1977,   t_1978;
/* u1_700 Output nets */
wire t_1979,   t_1980;
/* u2_701 Output nets */
wire t_1981,   t_1982,   t_1983;
/* u2_702 Output nets */
wire t_1984,   t_1985,   t_1986;
/* u2_703 Output nets */
wire t_1987,   t_1988,   t_1989;
/* u1_704 Output nets */
wire t_1990,   t_1991;
/* u2_705 Output nets */
wire t_1992,   t_1993,   t_1994;
/* u2_706 Output nets */
wire t_1995,   t_1996,   t_1997;
/* u2_707 Output nets */
wire t_1998,   t_1999,   t_2000;
/* u1_708 Output nets */
wire t_2001,   t_2002;
/* u2_709 Output nets */
wire t_2003,   t_2004,   t_2005;
/* u2_710 Output nets */
wire t_2006,   t_2007,   t_2008;
/* u2_711 Output nets */
wire t_2009,   t_2010,   t_2011;
/* u1_712 Output nets */
wire t_2012,   t_2013;
/* u2_713 Output nets */
wire t_2014,   t_2015,   t_2016;
/* u2_714 Output nets */
wire t_2017,   t_2018,   t_2019;
/* u2_715 Output nets */
wire t_2020,   t_2021,   t_2022;
/* u1_716 Output nets */
wire t_2023,   t_2024;
/* u2_717 Output nets */
wire t_2025,   t_2026,   t_2027;
/* u2_718 Output nets */
wire t_2028,   t_2029,   t_2030;
/* u2_719 Output nets */
wire t_2031,   t_2032,   t_2033;
/* u2_720 Output nets */
wire t_2034,   t_2035,   t_2036;
/* u2_721 Output nets */
wire t_2037,   t_2038,   t_2039;
/* u2_722 Output nets */
wire t_2040,   t_2041,   t_2042;
/* u2_723 Output nets */
wire t_2043,   t_2044,   t_2045;
/* u1_724 Output nets */
wire t_2046,   t_2047;
/* u2_725 Output nets */
wire t_2048,   t_2049,   t_2050;
/* u2_726 Output nets */
wire t_2051,   t_2052,   t_2053;
/* u2_727 Output nets */
wire t_2054,   t_2055,   t_2056;
/* u1_728 Output nets */
wire t_2057,   t_2058;
/* u2_729 Output nets */
wire t_2059,   t_2060,   t_2061;
/* u2_730 Output nets */
wire t_2062,   t_2063,   t_2064;
/* u2_731 Output nets */
wire t_2065,   t_2066,   t_2067;
/* u2_732 Output nets */
wire t_2068,   t_2069,   t_2070;
/* u2_733 Output nets */
wire t_2071,   t_2072,   t_2073;
/* u2_734 Output nets */
wire t_2074,   t_2075,   t_2076;
/* u2_735 Output nets */
wire t_2077,   t_2078,   t_2079;
/* u2_736 Output nets */
wire t_2080,   t_2081,   t_2082;
/* u2_737 Output nets */
wire t_2083,   t_2084,   t_2085;
/* u2_738 Output nets */
wire t_2086,   t_2087,   t_2088;
/* u2_739 Output nets */
wire t_2089,   t_2090,   t_2091;
/* u2_740 Output nets */
wire t_2092,   t_2093,   t_2094;
/* u2_741 Output nets */
wire t_2095,   t_2096,   t_2097;
/* u2_742 Output nets */
wire t_2098,   t_2099,   t_2100;
/* u2_743 Output nets */
wire t_2101,   t_2102,   t_2103;
/* u2_744 Output nets */
wire t_2104,   t_2105,   t_2106;
/* u2_745 Output nets */
wire t_2107,   t_2108,   t_2109;
/* u2_746 Output nets */
wire t_2110,   t_2111,   t_2112;
/* u2_747 Output nets */
wire t_2113,   t_2114,   t_2115;
/* u2_748 Output nets */
wire t_2116,   t_2117,   t_2118;
/* u2_749 Output nets */
wire t_2119,   t_2120,   t_2121;
/* u2_750 Output nets */
wire t_2122,   t_2123,   t_2124;
/* u2_751 Output nets */
wire t_2125,   t_2126,   t_2127;
/* u2_752 Output nets */
wire t_2128,   t_2129,   t_2130;
/* u2_753 Output nets */
wire t_2131,   t_2132,   t_2133;
/* u2_754 Output nets */
wire t_2134,   t_2135,   t_2136;
/* u2_755 Output nets */
wire t_2137,   t_2138,   t_2139;
/* u2_756 Output nets */
wire t_2140,   t_2141,   t_2142;
/* u2_757 Output nets */
wire t_2143,   t_2144,   t_2145;
/* u2_758 Output nets */
wire t_2146,   t_2147,   t_2148;
/* u2_759 Output nets */
wire t_2149,   t_2150,   t_2151;
/* u2_760 Output nets */
wire t_2152,   t_2153,   t_2154;
/* u2_761 Output nets */
wire t_2155,   t_2156,   t_2157;
/* u2_762 Output nets */
wire t_2158,   t_2159,   t_2160;
/* u2_763 Output nets */
wire t_2161,   t_2162,   t_2163;
/* u2_764 Output nets */
wire t_2164,   t_2165,   t_2166;
/* u2_765 Output nets */
wire t_2167,   t_2168,   t_2169;
/* u2_766 Output nets */
wire t_2170,   t_2171,   t_2172;
/* u2_767 Output nets */
wire t_2173,   t_2174,   t_2175;
/* u1_768 Output nets */
wire t_2176,   t_2177;
/* u2_769 Output nets */
wire t_2178,   t_2179,   t_2180;
/* u2_770 Output nets */
wire t_2181,   t_2182,   t_2183;
/* u2_771 Output nets */
wire t_2184,   t_2185,   t_2186;
/* u1_772 Output nets */
wire t_2187,   t_2188;
/* u2_773 Output nets */
wire t_2189,   t_2190,   t_2191;
/* u2_774 Output nets */
wire t_2192,   t_2193,   t_2194;
/* u2_775 Output nets */
wire t_2195,   t_2196,   t_2197;
/* u1_776 Output nets */
wire t_2198,   t_2199;
/* u2_777 Output nets */
wire t_2200,   t_2201,   t_2202;
/* u2_778 Output nets */
wire t_2203,   t_2204,   t_2205;
/* u2_779 Output nets */
wire t_2206,   t_2207,   t_2208;
/* u1_780 Output nets */
wire t_2209,   t_2210;
/* u2_781 Output nets */
wire t_2211,   t_2212,   t_2213;
/* u2_782 Output nets */
wire t_2214,   t_2215,   t_2216;
/* u2_783 Output nets */
wire t_2217,   t_2218,   t_2219;
/* u1_784 Output nets */
wire t_2220,   t_2221;
/* u2_785 Output nets */
wire t_2222,   t_2223,   t_2224;
/* u2_786 Output nets */
wire t_2225,   t_2226,   t_2227;
/* u2_787 Output nets */
wire t_2228,   t_2229,   t_2230;
/* u1_788 Output nets */
wire t_2231,   t_2232;
/* u2_789 Output nets */
wire t_2233,   t_2234,   t_2235;
/* u2_790 Output nets */
wire t_2236,   t_2237,   t_2238;
/* u2_791 Output nets */
wire t_2239,   t_2240,   t_2241;
/* u1_792 Output nets */
wire t_2242,   t_2243;
/* u2_793 Output nets */
wire t_2244,   t_2245,   t_2246;
/* u2_794 Output nets */
wire t_2247,   t_2248,   t_2249;
/* u2_795 Output nets */
wire t_2250,   t_2251,   t_2252;
/* u1_796 Output nets */
wire t_2253,   t_2254;
/* u2_797 Output nets */
wire t_2255,   t_2256,   t_2257;
/* u2_798 Output nets */
wire t_2258,   t_2259,   t_2260;
/* u2_799 Output nets */
wire t_2261,   t_2262,   t_2263;
/* u0_800 Output nets */
wire t_2264,   t_2265;
/* u2_801 Output nets */
wire t_2266,   t_2267,   t_2268;
/* u2_802 Output nets */
wire t_2269,   t_2270,   t_2271;
/* u2_803 Output nets */
wire t_2272,   t_2273,   t_2274;
/* u0_804 Output nets */
wire t_2275,   t_2276;
/* u2_805 Output nets */
wire t_2277,   t_2278,   t_2279;
/* u2_806 Output nets */
wire t_2280,   t_2281,   t_2282;
/* u2_807 Output nets */
wire t_2283,   t_2284,   t_2285;
/* u0_808 Output nets */
wire t_2286,   t_2287;
/* u2_809 Output nets */
wire t_2288,   t_2289,   t_2290;
/* u2_810 Output nets */
wire t_2291,   t_2292,   t_2293;
/* u2_811 Output nets */
wire t_2294,   t_2295,   t_2296;
/* u0_812 Output nets */
wire t_2297,   t_2298;
/* u2_813 Output nets */
wire t_2299,   t_2300,   t_2301;
/* u2_814 Output nets */
wire t_2302,   t_2303,   t_2304;
/* u2_815 Output nets */
wire t_2305,   t_2306,   t_2307;
/* u0_816 Output nets */
wire t_2308,   t_2309;
/* u2_817 Output nets */
wire t_2310,   t_2311,   t_2312;
/* u2_818 Output nets */
wire t_2313,   t_2314,   t_2315;
/* u2_819 Output nets */
wire t_2316,   t_2317,   t_2318;
/* u2_820 Output nets */
wire t_2319,   t_2320,   t_2321;
/* u2_821 Output nets */
wire t_2322,   t_2323,   t_2324;
/* u2_822 Output nets */
wire t_2325,   t_2326,   t_2327;
/* u2_823 Output nets */
wire t_2328,   t_2329,   t_2330;
/* u2_824 Output nets */
wire t_2331,   t_2332,   t_2333;
/* u2_825 Output nets */
wire t_2334,   t_2335,   t_2336;
/* u2_826 Output nets */
wire t_2337,   t_2338,   t_2339;
/* u2_827 Output nets */
wire t_2340,   t_2341,   t_2342;
/* u1_828 Output nets */
wire t_2343,   t_2344;
/* u2_829 Output nets */
wire t_2345,   t_2346,   t_2347;
/* u2_830 Output nets */
wire t_2348,   t_2349,   t_2350;
/* u1_831 Output nets */
wire t_2351,   t_2352;
/* u2_832 Output nets */
wire t_2353,   t_2354,   t_2355;
/* u2_833 Output nets */
wire t_2356,   t_2357,   t_2358;
/* u1_834 Output nets */
wire t_2359,   t_2360;
/* u2_835 Output nets */
wire t_2361,   t_2362,   t_2363;
/* u2_836 Output nets */
wire t_2364,   t_2365,   t_2366;
/* u1_837 Output nets */
wire t_2367,   t_2368;
/* u2_838 Output nets */
wire t_2369,   t_2370,   t_2371;
/* u2_839 Output nets */
wire t_2372,   t_2373,   t_2374;
/* u1_840 Output nets */
wire t_2375,   t_2376;
/* u2_841 Output nets */
wire t_2377,   t_2378,   t_2379;
/* u2_842 Output nets */
wire t_2380,   t_2381,   t_2382;
/* u1_843 Output nets */
wire t_2383,   t_2384;
/* u2_844 Output nets */
wire t_2385,   t_2386,   t_2387;
/* u2_845 Output nets */
wire t_2388,   t_2389,   t_2390;
/* u1_846 Output nets */
wire t_2391,   t_2392;
/* u2_847 Output nets */
wire t_2393,   t_2394,   t_2395;
/* u2_848 Output nets */
wire t_2396,   t_2397,   t_2398;
/* u1_849 Output nets */
wire t_2399,   t_2400;
/* u2_850 Output nets */
wire t_2401,   t_2402,   t_2403;
/* u2_851 Output nets */
wire t_2404,   t_2405,   t_2406;
/* u0_852 Output nets */
wire t_2407,   t_2408;
/* u2_853 Output nets */
wire t_2409,   t_2410,   t_2411;
/* u2_854 Output nets */
wire t_2412,   t_2413,   t_2414;
/* u0_855 Output nets */
wire t_2415,   t_2416;
/* u2_856 Output nets */
wire t_2417,   t_2418,   t_2419;
/* u2_857 Output nets */
wire t_2420,   t_2421,   t_2422;
/* u0_858 Output nets */
wire t_2423,   t_2424;
/* u2_859 Output nets */
wire t_2425,   t_2426,   t_2427;
/* u2_860 Output nets */
wire t_2428,   t_2429,   t_2430;
/* u0_861 Output nets */
wire t_2431,   t_2432;
/* u2_862 Output nets */
wire t_2433,   t_2434,   t_2435;
/* u2_863 Output nets */
wire t_2436,   t_2437,   t_2438;
/* u0_864 Output nets */
wire t_2439,   t_2440;
/* u2_865 Output nets */
wire t_2441,   t_2442,   t_2443;
/* u2_866 Output nets */
wire t_2444,   t_2445,   t_2446;
/* u2_867 Output nets */
wire t_2447,   t_2448,   t_2449;
/* u2_868 Output nets */
wire t_2450,   t_2451,   t_2452;
/* u2_869 Output nets */
wire t_2453,   t_2454,   t_2455;
/* u2_870 Output nets */
wire t_2456,   t_2457,   t_2458;
/* u2_871 Output nets */
wire t_2459,   t_2460,   t_2461;
/* u1_872 Output nets */
wire t_2462,   t_2463;
/* u2_873 Output nets */
wire t_2464,   t_2465,   t_2466;
/* u1_874 Output nets */
wire t_2467,   t_2468;
/* u2_875 Output nets */
wire t_2469,   t_2470,   t_2471;
/* u1_876 Output nets */
wire t_2472,   t_2473;
/* u2_877 Output nets */
wire t_2474,   t_2475,   t_2476;
/* u1_878 Output nets */
wire t_2477,   t_2478;
/* u2_879 Output nets */
wire t_2479,   t_2480,   t_2481;
/* u1_880 Output nets */
wire t_2482,   t_2483;
/* u2_881 Output nets */
wire t_2484,   t_2485,   t_2486;
/* u1_882 Output nets */
wire t_2487,   t_2488;
/* u2_883 Output nets */
wire t_2489,   t_2490,   t_2491;
/* u1_884 Output nets */
wire t_2492,   t_2493;
/* u2_885 Output nets */
wire t_2494,   t_2495,   t_2496;
/* u1_886 Output nets */
wire t_2497,   t_2498;
/* u2_887 Output nets */
wire t_2499,   t_2500,   t_2501;
/* u0_888 Output nets */
wire t_2502,   t_2503;
/* u2_889 Output nets */
wire t_2504,   t_2505,   t_2506;
/* u0_890 Output nets */
wire t_2507,   t_2508;
/* u2_891 Output nets */
wire t_2509,   t_2510,   t_2511;
/* u0_892 Output nets */
wire t_2512,   t_2513;
/* u2_893 Output nets */
wire t_2514,   t_2515,   t_2516;
/* u0_894 Output nets */
wire t_2517,   t_2518;
/* u2_895 Output nets */
wire t_2519,   t_2520,   t_2521;
/* u0_896 Output nets */
wire t_2522,   t_2523;
/* u2_897 Output nets */
wire t_2524,   t_2525,   t_2526;
/* u2_898 Output nets */
wire t_2527,   t_2528,   t_2529;
/* u2_899 Output nets */
wire t_2530,   t_2531,   t_2532;
/* u1_900 Output nets */
wire t_2533,   t_2534;
/* u1_901 Output nets */
wire t_2535,   t_2536;
/* u1_902 Output nets */
wire t_2537,   t_2538;
/* u1_903 Output nets */
wire t_2539,   t_2540;
/* u1_904 Output nets */
wire t_2541,   t_2542;
/* u0_905 Output nets */
wire t_2543,   t_2544;
/* u1_906 Output nets */
wire t_2545,   t_2546;
/* u0_907 Output nets */
wire t_2547,   t_2548;
/* u0_908 Output nets */
wire t_2549,   t_2550;
/* u0_909 Output nets */
wire t_2551;

/* compress stage 2 */
half_adder u0_590(.a(t_1), .b(s_1_0), .o(t_1681), .cout(t_1682));
half_adder u0_591(.a(t_3), .b(t_4), .o(t_1683), .cout(t_1684));
compressor_3_2 u1_592(.a(t_7), .b(t_9), .cin(s_5_2), .o(t_1685), .cout(t_1686));
half_adder u0_593(.a(t_10), .b(t_11), .o(t_1687), .cout(t_1688));
half_adder u0_594(.a(t_12), .b(t_14), .o(t_1689), .cout(t_1690));
compressor_3_2 u1_595(.a(t_15), .b(t_20), .cin(t_17), .o(t_1691), .cout(t_1692));
compressor_3_2 u1_596(.a(t_18), .b(t_25), .cin(t_22), .o(t_1693), .cout(t_1694));
compressor_4_2 u2_597(.a(t_23), .b(t_30), .c(t_27), .d(s_10_6), .cin(t_1694), .o(t_1695), .co(t_1696), .cout(t_1697));
compressor_3_2 u1_598(.a(t_35), .b(t_32), .cin(t_1697), .o(t_1698), .cout(t_1699));
compressor_3_2 u1_599(.a(t_33), .b(t_40), .cin(t_37), .o(t_1700), .cout(t_1701));
compressor_4_2 u2_600(.a(t_38), .b(t_46), .c(t_43), .d(s_13_6), .cin(t_1701), .o(t_1702), .co(t_1703), .cout(t_1704));
compressor_4_2 u2_601(.a(t_44), .b(t_51), .c(t_48), .d(s_14_8), .cin(t_1704), .o(t_1705), .co(t_1706), .cout(t_1707));
compressor_4_2 u2_602(.a(t_52), .b(t_49), .c(t_57), .d(t_54), .cin(t_1707), .o(t_1708), .co(t_1709), .cout(t_1710));
compressor_4_2 u2_603(.a(t_55), .b(t_66), .c(t_63), .d(t_60), .cin(t_1710), .o(t_1711), .co(t_1712), .cout(t_1713));
compressor_4_2 u2_604(.a(t_61), .b(t_74), .c(t_71), .d(t_68), .cin(t_1713), .o(t_1714), .co(t_1715), .cout(t_1716));
compressor_4_2 u2_605(.a(t_82), .b(t_79), .c(t_76), .d(s_18_10), .cin(t_1716), .o(t_1717), .co(t_1718), .cout(t_1719));
half_adder u0_606(.a(t_72), .b(t_69), .o(t_1720), .cout(t_1721));
compressor_4_2 u2_607(.a(t_90), .b(t_87), .c(t_84), .d(t_1719), .cin(t_1721), .o(t_1722), .co(t_1723), .cout(t_1724));
half_adder u0_608(.a(t_80), .b(t_77), .o(t_1725), .cout(t_1726));
compressor_4_2 u2_609(.a(t_98), .b(t_95), .c(t_92), .d(t_1724), .cin(t_1726), .o(t_1727), .co(t_1728), .cout(t_1729));
half_adder u0_610(.a(t_88), .b(t_85), .o(t_1730), .cout(t_1731));
compressor_4_2 u2_611(.a(t_104), .b(t_101), .c(s_21_10), .d(t_1729), .cin(t_1731), .o(t_1732), .co(t_1733), .cout(t_1734));
compressor_3_2 u1_612(.a(t_96), .b(t_93), .cin(t_107), .o(t_1735), .cout(t_1736));
compressor_4_2 u2_613(.a(t_112), .b(t_109), .c(s_22_12), .d(t_1734), .cin(t_1736), .o(t_1737), .co(t_1738), .cout(t_1739));
compressor_3_2 u1_614(.a(t_105), .b(t_102), .cin(t_115), .o(t_1740), .cout(t_1741));
compressor_4_2 u2_615(.a(t_124), .b(t_121), .c(t_118), .d(t_1739), .cin(t_1741), .o(t_1742), .co(t_1743), .cout(t_1744));
compressor_3_2 u1_616(.a(t_116), .b(t_113), .cin(t_110), .o(t_1745), .cout(t_1746));
compressor_4_2 u2_617(.a(t_133), .b(t_130), .c(t_127), .d(t_1744), .cin(t_1746), .o(t_1747), .co(t_1748), .cout(t_1749));
compressor_3_2 u1_618(.a(t_122), .b(t_119), .cin(t_136), .o(t_1750), .cout(t_1751));
compressor_4_2 u2_619(.a(t_144), .b(t_141), .c(t_138), .d(t_1749), .cin(t_1751), .o(t_1752), .co(t_1753), .cout(t_1754));
compressor_3_2 u1_620(.a(t_131), .b(t_128), .cin(t_147), .o(t_1755), .cout(t_1756));
compressor_4_2 u2_621(.a(t_152), .b(t_149), .c(s_26_14), .d(t_1754), .cin(t_1756), .o(t_1757), .co(t_1758), .cout(t_1759));
compressor_4_2 u2_622(.a(t_145), .b(t_142), .c(t_139), .d(t_158), .cin(t_155), .o(t_1760), .co(t_1761), .cout(t_1762));
compressor_4_2 u2_623(.a(t_166), .b(t_163), .c(t_160), .d(t_1759), .cin(t_1762), .o(t_1763), .co(t_1764), .cout(t_1765));
compressor_3_2 u1_624(.a(t_153), .b(t_150), .cin(t_169), .o(t_1766), .cout(t_1767));
compressor_4_2 u2_625(.a(t_177), .b(t_174), .c(t_171), .d(t_1765), .cin(t_1767), .o(t_1768), .co(t_1769), .cout(t_1770));
compressor_3_2 u1_626(.a(t_164), .b(t_161), .cin(t_180), .o(t_1771), .cout(t_1772));
compressor_4_2 u2_627(.a(t_186), .b(t_183), .c(s_29_14), .d(t_1770), .cin(t_1772), .o(t_1773), .co(t_1774), .cout(t_1775));
compressor_4_2 u2_628(.a(t_178), .b(t_175), .c(t_172), .d(t_192), .cin(t_189), .o(t_1776), .co(t_1777), .cout(t_1778));
compressor_4_2 u2_629(.a(t_197), .b(t_194), .c(s_30_16), .d(t_1775), .cin(t_1778), .o(t_1779), .co(t_1780), .cout(t_1781));
compressor_4_2 u2_630(.a(t_190), .b(t_187), .c(t_184), .d(t_203), .cin(t_200), .o(t_1782), .co(t_1783), .cout(t_1784));
compressor_4_2 u2_631(.a(t_212), .b(t_209), .c(t_206), .d(t_1781), .cin(t_1784), .o(t_1785), .co(t_1786), .cout(t_1787));
compressor_4_2 u2_632(.a(t_204), .b(t_201), .c(t_198), .d(t_195), .cin(t_215), .o(t_1788), .co(t_1789), .cout(t_1790));
compressor_4_2 u2_633(.a(t_224), .b(t_221), .c(t_218), .d(t_1787), .cin(t_1790), .o(t_1791), .co(t_1792), .cout(t_1793));
compressor_4_2 u2_634(.a(t_213), .b(t_210), .c(t_207), .d(t_230), .cin(t_227), .o(t_1794), .co(t_1795), .cout(t_1796));
compressor_4_2 u2_635(.a(t_238), .b(t_235), .c(t_232), .d(t_1793), .cin(t_1796), .o(t_1797), .co(t_1798), .cout(t_1799));
compressor_4_2 u2_636(.a(t_225), .b(t_222), .c(t_219), .d(t_244), .cin(t_241), .o(t_1800), .co(t_1801), .cout(t_1802));
compressor_4_2 u2_637(.a(t_249), .b(t_246), .c(s_34_18), .d(t_1799), .cin(t_1802), .o(t_1803), .co(t_1804), .cout(t_1805));
compressor_4_2 u2_638(.a(t_236), .b(t_233), .c(t_258), .d(t_255), .cin(t_252), .o(t_1806), .co(t_1807), .cout(t_1808));
half_adder u0_639(.a(t_242), .b(t_239), .o(t_1809), .cout(t_1810));
compressor_4_2 u2_640(.a(t_266), .b(t_263), .c(t_260), .d(t_1805), .cin(t_1808), .o(t_1811), .co(t_1812), .cout(t_1813));
compressor_4_2 u2_641(.a(t_250), .b(t_247), .c(t_272), .d(t_269), .cin(t_1810), .o(t_1814), .co(t_1815), .cout(t_1816));
half_adder u0_642(.a(t_256), .b(t_253), .o(t_1817), .cout(t_1818));
compressor_4_2 u2_643(.a(t_280), .b(t_277), .c(t_274), .d(t_1813), .cin(t_1816), .o(t_1819), .co(t_1820), .cout(t_1821));
compressor_4_2 u2_644(.a(t_264), .b(t_261), .c(t_286), .d(t_283), .cin(t_1818), .o(t_1822), .co(t_1823), .cout(t_1824));
half_adder u0_645(.a(t_270), .b(t_267), .o(t_1825), .cout(t_1826));
compressor_4_2 u2_646(.a(t_292), .b(t_289), .c(s_37_18), .d(t_1821), .cin(t_1824), .o(t_1827), .co(t_1828), .cout(t_1829));
compressor_4_2 u2_647(.a(t_275), .b(t_301), .c(t_298), .d(t_295), .cin(t_1826), .o(t_1830), .co(t_1831), .cout(t_1832));
compressor_3_2 u1_648(.a(t_284), .b(t_281), .cin(t_278), .o(t_1833), .cout(t_1834));
compressor_4_2 u2_649(.a(t_306), .b(t_303), .c(s_38_20), .d(t_1829), .cin(t_1832), .o(t_1835), .co(t_1836), .cout(t_1837));
compressor_4_2 u2_650(.a(t_290), .b(t_315), .c(t_312), .d(t_309), .cin(t_1834), .o(t_1838), .co(t_1839), .cout(t_1840));
compressor_3_2 u1_651(.a(t_299), .b(t_296), .cin(t_293), .o(t_1841), .cout(t_1842));
compressor_4_2 u2_652(.a(t_324), .b(t_321), .c(t_318), .d(t_1837), .cin(t_1840), .o(t_1843), .co(t_1844), .cout(t_1845));
compressor_4_2 u2_653(.a(t_307), .b(t_304), .c(t_330), .d(t_327), .cin(t_1842), .o(t_1846), .co(t_1847), .cout(t_1848));
compressor_3_2 u1_654(.a(t_316), .b(t_313), .cin(t_310), .o(t_1849), .cout(t_1850));
compressor_4_2 u2_655(.a(t_339), .b(t_336), .c(t_333), .d(t_1845), .cin(t_1848), .o(t_1851), .co(t_1852), .cout(t_1853));
compressor_4_2 u2_656(.a(t_319), .b(t_348), .c(t_345), .d(t_342), .cin(t_1850), .o(t_1854), .co(t_1855), .cout(t_1856));
compressor_3_2 u1_657(.a(t_328), .b(t_325), .cin(t_322), .o(t_1857), .cout(t_1858));
compressor_4_2 u2_658(.a(t_356), .b(t_353), .c(t_350), .d(t_1853), .cin(t_1856), .o(t_1859), .co(t_1860), .cout(t_1861));
compressor_4_2 u2_659(.a(t_334), .b(t_365), .c(t_362), .d(t_359), .cin(t_1858), .o(t_1862), .co(t_1863), .cout(t_1864));
compressor_3_2 u1_660(.a(t_343), .b(t_340), .cin(t_337), .o(t_1865), .cout(t_1866));
compressor_4_2 u2_661(.a(t_370), .b(t_367), .c(s_42_22), .d(t_1861), .cin(t_1864), .o(t_1867), .co(t_1868), .cout(t_1869));
compressor_4_2 u2_662(.a(t_382), .b(t_379), .c(t_376), .d(t_373), .cin(t_1866), .o(t_1870), .co(t_1871), .cout(t_1872));
compressor_4_2 u2_663(.a(t_363), .b(t_360), .c(t_357), .d(t_354), .cin(t_351), .o(t_1873), .co(t_1874), .cout(t_1875));
compressor_4_2 u2_664(.a(t_390), .b(t_387), .c(t_384), .d(t_1869), .cin(t_1872), .o(t_1876), .co(t_1877), .cout(t_1878));
compressor_4_2 u2_665(.a(t_368), .b(t_399), .c(t_396), .d(t_393), .cin(t_1875), .o(t_1879), .co(t_1880), .cout(t_1881));
compressor_3_2 u1_666(.a(t_377), .b(t_374), .cin(t_371), .o(t_1882), .cout(t_1883));
compressor_4_2 u2_667(.a(t_407), .b(t_404), .c(t_401), .d(t_1878), .cin(t_1881), .o(t_1884), .co(t_1885), .cout(t_1886));
compressor_4_2 u2_668(.a(t_385), .b(t_416), .c(t_413), .d(t_410), .cin(t_1883), .o(t_1887), .co(t_1888), .cout(t_1889));
compressor_3_2 u1_669(.a(t_394), .b(t_391), .cin(t_388), .o(t_1890), .cout(t_1891));
compressor_4_2 u2_670(.a(t_422), .b(t_419), .c(s_45_22), .d(t_1886), .cin(t_1889), .o(t_1892), .co(t_1893), .cout(t_1894));
compressor_4_2 u2_671(.a(t_434), .b(t_431), .c(t_428), .d(t_425), .cin(t_1891), .o(t_1895), .co(t_1896), .cout(t_1897));
compressor_4_2 u2_672(.a(t_414), .b(t_411), .c(t_408), .d(t_405), .cin(t_402), .o(t_1898), .co(t_1899), .cout(t_1900));
compressor_4_2 u2_673(.a(t_439), .b(t_436), .c(s_46_24), .d(t_1894), .cin(t_1897), .o(t_1901), .co(t_1902), .cout(t_1903));
compressor_4_2 u2_674(.a(t_451), .b(t_448), .c(t_445), .d(t_442), .cin(t_1900), .o(t_1904), .co(t_1905), .cout(t_1906));
compressor_4_2 u2_675(.a(t_432), .b(t_429), .c(t_426), .d(t_423), .cin(t_420), .o(t_1907), .co(t_1908), .cout(t_1909));
compressor_4_2 u2_676(.a(t_460), .b(t_457), .c(t_454), .d(t_1903), .cin(t_1906), .o(t_1910), .co(t_1911), .cout(t_1912));
compressor_4_2 u2_677(.a(t_437), .b(t_469), .c(t_466), .d(t_463), .cin(t_1909), .o(t_1913), .co(t_1914), .cout(t_1915));
compressor_4_2 u2_678(.a(t_452), .b(t_449), .c(t_446), .d(t_443), .cin(t_440), .o(t_1916), .co(t_1917), .cout(t_1918));
compressor_4_2 u2_679(.a(t_478), .b(t_475), .c(t_472), .d(t_1912), .cin(t_1915), .o(t_1919), .co(t_1920), .cout(t_1921));
compressor_4_2 u2_680(.a(t_490), .b(t_487), .c(t_484), .d(t_481), .cin(t_1918), .o(t_1922), .co(t_1923), .cout(t_1924));
compressor_4_2 u2_681(.a(t_467), .b(t_464), .c(t_461), .d(t_458), .cin(t_455), .o(t_1925), .co(t_1926), .cout(t_1927));
compressor_4_2 u2_682(.a(t_498), .b(t_495), .c(t_492), .d(t_1921), .cin(t_1924), .o(t_1928), .co(t_1929), .cout(t_1930));
compressor_4_2 u2_683(.a(t_510), .b(t_507), .c(t_504), .d(t_501), .cin(t_1927), .o(t_1931), .co(t_1932), .cout(t_1933));
compressor_4_2 u2_684(.a(t_485), .b(t_482), .c(t_479), .d(t_476), .cin(t_473), .o(t_1934), .co(t_1935), .cout(t_1936));
compressor_4_2 u2_685(.a(t_515), .b(t_512), .c(s_50_26), .d(t_1930), .cin(t_1933), .o(t_1937), .co(t_1938), .cout(t_1939));
compressor_4_2 u2_686(.a(t_527), .b(t_524), .c(t_521), .d(t_518), .cin(t_1936), .o(t_1940), .co(t_1941), .cout(t_1942));
compressor_4_2 u2_687(.a(t_502), .b(t_499), .c(t_496), .d(t_493), .cin(t_530), .o(t_1943), .co(t_1944), .cout(t_1945));
half_adder u0_688(.a(t_508), .b(t_505), .o(t_1946), .cout(t_1947));
compressor_4_2 u2_689(.a(t_538), .b(t_535), .c(t_532), .d(t_1939), .cin(t_1942), .o(t_1948), .co(t_1949), .cout(t_1950));
compressor_4_2 u2_690(.a(t_547), .b(t_544), .c(t_541), .d(t_1945), .cin(t_1947), .o(t_1951), .co(t_1952), .cout(t_1953));
compressor_4_2 u2_691(.a(t_522), .b(t_519), .c(t_516), .d(t_513), .cin(t_550), .o(t_1954), .co(t_1955), .cout(t_1956));
half_adder u0_692(.a(t_528), .b(t_525), .o(t_1957), .cout(t_1958));
compressor_4_2 u2_693(.a(t_558), .b(t_555), .c(t_552), .d(t_1950), .cin(t_1953), .o(t_1959), .co(t_1960), .cout(t_1961));
compressor_4_2 u2_694(.a(t_567), .b(t_564), .c(t_561), .d(t_1956), .cin(t_1958), .o(t_1962), .co(t_1963), .cout(t_1964));
compressor_4_2 u2_695(.a(t_542), .b(t_539), .c(t_536), .d(t_533), .cin(t_570), .o(t_1965), .co(t_1966), .cout(t_1967));
half_adder u0_696(.a(t_548), .b(t_545), .o(t_1968), .cout(t_1969));
compressor_4_2 u2_697(.a(t_576), .b(t_573), .c(s_53_26), .d(t_1961), .cin(t_1964), .o(t_1970), .co(t_1971), .cout(t_1972));
compressor_4_2 u2_698(.a(t_585), .b(t_582), .c(t_579), .d(t_1967), .cin(t_1969), .o(t_1973), .co(t_1974), .cout(t_1975));
compressor_4_2 u2_699(.a(t_559), .b(t_556), .c(t_553), .d(t_591), .cin(t_588), .o(t_1976), .co(t_1977), .cout(t_1978));
compressor_3_2 u1_700(.a(t_568), .b(t_565), .cin(t_562), .o(t_1979), .cout(t_1980));
compressor_4_2 u2_701(.a(t_596), .b(t_593), .c(s_54_28), .d(t_1972), .cin(t_1975), .o(t_1981), .co(t_1982), .cout(t_1983));
compressor_4_2 u2_702(.a(t_605), .b(t_602), .c(t_599), .d(t_1978), .cin(t_1980), .o(t_1984), .co(t_1985), .cout(t_1986));
compressor_4_2 u2_703(.a(t_580), .b(t_577), .c(t_574), .d(t_611), .cin(t_608), .o(t_1987), .co(t_1988), .cout(t_1989));
compressor_3_2 u1_704(.a(t_589), .b(t_586), .cin(t_583), .o(t_1990), .cout(t_1991));
compressor_4_2 u2_705(.a(t_620), .b(t_617), .c(t_614), .d(t_1983), .cin(t_1986), .o(t_1992), .co(t_1993), .cout(t_1994));
compressor_4_2 u2_706(.a(t_629), .b(t_626), .c(t_623), .d(t_1989), .cin(t_1991), .o(t_1995), .co(t_1996), .cout(t_1997));
compressor_4_2 u2_707(.a(t_603), .b(t_600), .c(t_597), .d(t_594), .cin(t_632), .o(t_1998), .co(t_1999), .cout(t_2000));
compressor_3_2 u1_708(.a(t_612), .b(t_609), .cin(t_606), .o(t_2001), .cout(t_2002));
compressor_4_2 u2_709(.a(t_641), .b(t_638), .c(t_635), .d(t_1994), .cin(t_1997), .o(t_2003), .co(t_2004), .cout(t_2005));
compressor_4_2 u2_710(.a(t_650), .b(t_647), .c(t_644), .d(t_2000), .cin(t_2002), .o(t_2006), .co(t_2007), .cout(t_2008));
compressor_4_2 u2_711(.a(t_621), .b(t_618), .c(t_615), .d(t_656), .cin(t_653), .o(t_2009), .co(t_2010), .cout(t_2011));
compressor_3_2 u1_712(.a(t_630), .b(t_627), .cin(t_624), .o(t_2012), .cout(t_2013));
compressor_4_2 u2_713(.a(t_664), .b(t_661), .c(t_658), .d(t_2005), .cin(t_2008), .o(t_2014), .co(t_2015), .cout(t_2016));
compressor_4_2 u2_714(.a(t_673), .b(t_670), .c(t_667), .d(t_2011), .cin(t_2013), .o(t_2017), .co(t_2018), .cout(t_2019));
compressor_4_2 u2_715(.a(t_642), .b(t_639), .c(t_636), .d(t_679), .cin(t_676), .o(t_2020), .co(t_2021), .cout(t_2022));
compressor_3_2 u1_716(.a(t_651), .b(t_648), .cin(t_645), .o(t_2023), .cout(t_2024));
compressor_4_2 u2_717(.a(t_684), .b(t_681), .c(s_58_30), .d(t_2016), .cin(t_2019), .o(t_2025), .co(t_2026), .cout(t_2027));
compressor_4_2 u2_718(.a(t_693), .b(t_690), .c(t_687), .d(t_2022), .cin(t_2024), .o(t_2028), .co(t_2029), .cout(t_2030));
compressor_4_2 u2_719(.a(t_662), .b(t_659), .c(t_702), .d(t_699), .cin(t_696), .o(t_2031), .co(t_2032), .cout(t_2033));
compressor_4_2 u2_720(.a(t_677), .b(t_674), .c(t_671), .d(t_668), .cin(t_665), .o(t_2034), .co(t_2035), .cout(t_2036));
compressor_4_2 u2_721(.a(t_710), .b(t_707), .c(t_704), .d(t_2027), .cin(t_2030), .o(t_2037), .co(t_2038), .cout(t_2039));
compressor_4_2 u2_722(.a(t_719), .b(t_716), .c(t_713), .d(t_2033), .cin(t_2036), .o(t_2040), .co(t_2041), .cout(t_2042));
compressor_4_2 u2_723(.a(t_688), .b(t_685), .c(t_682), .d(t_725), .cin(t_722), .o(t_2043), .co(t_2044), .cout(t_2045));
compressor_3_2 u1_724(.a(t_697), .b(t_694), .cin(t_691), .o(t_2046), .cout(t_2047));
compressor_4_2 u2_725(.a(t_733), .b(t_730), .c(t_727), .d(t_2039), .cin(t_2042), .o(t_2048), .co(t_2049), .cout(t_2050));
compressor_4_2 u2_726(.a(t_742), .b(t_739), .c(t_736), .d(t_2045), .cin(t_2047), .o(t_2051), .co(t_2052), .cout(t_2053));
compressor_4_2 u2_727(.a(t_711), .b(t_708), .c(t_705), .d(t_748), .cin(t_745), .o(t_2054), .co(t_2055), .cout(t_2056));
compressor_3_2 u1_728(.a(t_720), .b(t_717), .cin(t_714), .o(t_2057), .cout(t_2058));
compressor_4_2 u2_729(.a(t_754), .b(t_751), .c(s_61_30), .d(t_2050), .cin(t_2053), .o(t_2059), .co(t_2060), .cout(t_2061));
compressor_4_2 u2_730(.a(t_763), .b(t_760), .c(t_757), .d(t_2056), .cin(t_2058), .o(t_2062), .co(t_2063), .cout(t_2064));
compressor_4_2 u2_731(.a(t_731), .b(t_728), .c(t_772), .d(t_769), .cin(t_766), .o(t_2065), .co(t_2066), .cout(t_2067));
compressor_4_2 u2_732(.a(t_746), .b(t_743), .c(t_740), .d(t_737), .cin(t_734), .o(t_2068), .co(t_2069), .cout(t_2070));
compressor_4_2 u2_733(.a(t_777), .b(t_774), .c(s_62_32), .d(t_2061), .cin(t_2064), .o(t_2071), .co(t_2072), .cout(t_2073));
compressor_4_2 u2_734(.a(t_786), .b(t_783), .c(t_780), .d(t_2067), .cin(t_2070), .o(t_2074), .co(t_2075), .cout(t_2076));
compressor_4_2 u2_735(.a(t_755), .b(t_752), .c(t_795), .d(t_792), .cin(t_789), .o(t_2077), .co(t_2078), .cout(t_2079));
compressor_4_2 u2_736(.a(t_770), .b(t_767), .c(t_764), .d(t_761), .cin(t_758), .o(t_2080), .co(t_2081), .cout(t_2082));
compressor_4_2 u2_737(.a(t_804), .b(t_801), .c(t_798), .d(t_2073), .cin(t_2076), .o(t_2083), .co(t_2084), .cout(t_2085));
compressor_4_2 u2_738(.a(t_813), .b(t_810), .c(t_807), .d(t_2079), .cin(t_2082), .o(t_2086), .co(t_2087), .cout(t_2088));
compressor_4_2 u2_739(.a(t_781), .b(t_778), .c(t_775), .d(t_819), .cin(t_816), .o(t_2089), .co(t_2090), .cout(t_2091));
compressor_4_2 u2_740(.a(t_796), .b(t_793), .c(t_790), .d(t_787), .cin(t_784), .o(t_2092), .co(t_2093), .cout(t_2094));
compressor_4_2 u2_741(.a(t_825), .b(t_822), .c(s_64_32), .d(t_2085), .cin(t_2088), .o(t_2095), .co(t_2096), .cout(t_2097));
compressor_4_2 u2_742(.a(t_834), .b(t_831), .c(t_828), .d(t_2091), .cin(t_2094), .o(t_2098), .co(t_2099), .cout(t_2100));
compressor_4_2 u2_743(.a(t_802), .b(t_799), .c(t_843), .d(t_840), .cin(t_837), .o(t_2101), .co(t_2102), .cout(t_2103));
compressor_4_2 u2_744(.a(t_817), .b(t_814), .c(t_811), .d(t_808), .cin(t_805), .o(t_2104), .co(t_2105), .cout(t_2106));
compressor_4_2 u2_745(.a(t_849), .b(t_846), .c(s_65_32), .d(t_2097), .cin(t_2100), .o(t_2107), .co(t_2108), .cout(t_2109));
compressor_4_2 u2_746(.a(t_858), .b(t_855), .c(t_852), .d(t_2103), .cin(t_2106), .o(t_2110), .co(t_2111), .cout(t_2112));
compressor_4_2 u2_747(.a(t_826), .b(t_823), .c(t_867), .d(t_864), .cin(t_861), .o(t_2113), .co(t_2114), .cout(t_2115));
compressor_4_2 u2_748(.a(t_841), .b(t_838), .c(t_835), .d(t_832), .cin(t_829), .o(t_2116), .co(t_2117), .cout(t_2118));
compressor_4_2 u2_749(.a(t_876), .b(t_873), .c(t_870), .d(t_2109), .cin(t_2112), .o(t_2119), .co(t_2120), .cout(t_2121));
compressor_4_2 u2_750(.a(t_885), .b(t_882), .c(t_879), .d(t_2115), .cin(t_2118), .o(t_2122), .co(t_2123), .cout(t_2124));
compressor_4_2 u2_751(.a(t_853), .b(t_850), .c(t_847), .d(t_891), .cin(t_888), .o(t_2125), .co(t_2126), .cout(t_2127));
compressor_4_2 u2_752(.a(t_868), .b(t_865), .c(t_862), .d(t_859), .cin(t_856), .o(t_2128), .co(t_2129), .cout(t_2130));
compressor_4_2 u2_753(.a(t_900), .b(t_897), .c(t_894), .d(t_2121), .cin(t_2124), .o(t_2131), .co(t_2132), .cout(t_2133));
compressor_4_2 u2_754(.a(t_909), .b(t_906), .c(t_903), .d(t_2127), .cin(t_2130), .o(t_2134), .co(t_2135), .cout(t_2136));
compressor_4_2 u2_755(.a(t_877), .b(t_874), .c(t_871), .d(t_915), .cin(t_912), .o(t_2137), .co(t_2138), .cout(t_2139));
compressor_4_2 u2_756(.a(t_892), .b(t_889), .c(t_886), .d(t_883), .cin(t_880), .o(t_2140), .co(t_2141), .cout(t_2142));
compressor_4_2 u2_757(.a(t_921), .b(t_918), .c(s_68_30), .d(t_2133), .cin(t_2136), .o(t_2143), .co(t_2144), .cout(t_2145));
compressor_4_2 u2_758(.a(t_930), .b(t_927), .c(t_924), .d(t_2139), .cin(t_2142), .o(t_2146), .co(t_2147), .cout(t_2148));
compressor_4_2 u2_759(.a(t_898), .b(t_895), .c(t_939), .d(t_936), .cin(t_933), .o(t_2149), .co(t_2150), .cout(t_2151));
compressor_4_2 u2_760(.a(t_913), .b(t_910), .c(t_907), .d(t_904), .cin(t_901), .o(t_2152), .co(t_2153), .cout(t_2154));
compressor_4_2 u2_761(.a(t_944), .b(t_941), .c(s_69_30), .d(t_2145), .cin(t_2148), .o(t_2155), .co(t_2156), .cout(t_2157));
compressor_4_2 u2_762(.a(t_953), .b(t_950), .c(t_947), .d(t_2151), .cin(t_2154), .o(t_2158), .co(t_2159), .cout(t_2160));
compressor_4_2 u2_763(.a(t_922), .b(t_919), .c(t_962), .d(t_959), .cin(t_956), .o(t_2161), .co(t_2162), .cout(t_2163));
compressor_4_2 u2_764(.a(t_937), .b(t_934), .c(t_931), .d(t_928), .cin(t_925), .o(t_2164), .co(t_2165), .cout(t_2166));
compressor_4_2 u2_765(.a(t_970), .b(t_967), .c(t_964), .d(t_2157), .cin(t_2160), .o(t_2167), .co(t_2168), .cout(t_2169));
compressor_4_2 u2_766(.a(t_979), .b(t_976), .c(t_973), .d(t_2163), .cin(t_2166), .o(t_2170), .co(t_2171), .cout(t_2172));
compressor_4_2 u2_767(.a(t_948), .b(t_945), .c(t_942), .d(t_985), .cin(t_982), .o(t_2173), .co(t_2174), .cout(t_2175));
compressor_3_2 u1_768(.a(t_957), .b(t_954), .cin(t_951), .o(t_2176), .cout(t_2177));
compressor_4_2 u2_769(.a(t_993), .b(t_990), .c(t_987), .d(t_2169), .cin(t_2172), .o(t_2178), .co(t_2179), .cout(t_2180));
compressor_4_2 u2_770(.a(t_1002), .b(t_999), .c(t_996), .d(t_2175), .cin(t_2177), .o(t_2181), .co(t_2182), .cout(t_2183));
compressor_4_2 u2_771(.a(t_971), .b(t_968), .c(t_965), .d(t_1008), .cin(t_1005), .o(t_2184), .co(t_2185), .cout(t_2186));
compressor_3_2 u1_772(.a(t_980), .b(t_977), .cin(t_974), .o(t_2187), .cout(t_2188));
compressor_4_2 u2_773(.a(t_1016), .b(t_1013), .c(t_1010), .d(t_2180), .cin(t_2183), .o(t_2189), .co(t_2190), .cout(t_2191));
compressor_4_2 u2_774(.a(t_1025), .b(t_1022), .c(t_1019), .d(t_2186), .cin(t_2188), .o(t_2192), .co(t_2193), .cout(t_2194));
compressor_4_2 u2_775(.a(t_994), .b(t_991), .c(t_988), .d(t_1031), .cin(t_1028), .o(t_2195), .co(t_2196), .cout(t_2197));
compressor_3_2 u1_776(.a(t_1003), .b(t_1000), .cin(t_997), .o(t_2198), .cout(t_2199));
compressor_4_2 u2_777(.a(t_1039), .b(t_1036), .c(t_1033), .d(t_2191), .cin(t_2194), .o(t_2200), .co(t_2201), .cout(t_2202));
compressor_4_2 u2_778(.a(t_1048), .b(t_1045), .c(t_1042), .d(t_2197), .cin(t_2199), .o(t_2203), .co(t_2204), .cout(t_2205));
compressor_4_2 u2_779(.a(t_1017), .b(t_1014), .c(t_1011), .d(t_1054), .cin(t_1051), .o(t_2206), .co(t_2207), .cout(t_2208));
compressor_3_2 u1_780(.a(t_1026), .b(t_1023), .cin(t_1020), .o(t_2209), .cout(t_2210));
compressor_4_2 u2_781(.a(t_1059), .b(t_1056), .c(s_74_27), .d(t_2202), .cin(t_2205), .o(t_2211), .co(t_2212), .cout(t_2213));
compressor_4_2 u2_782(.a(t_1068), .b(t_1065), .c(t_1062), .d(t_2208), .cin(t_2210), .o(t_2214), .co(t_2215), .cout(t_2216));
compressor_4_2 u2_783(.a(t_1040), .b(t_1037), .c(t_1034), .d(t_1074), .cin(t_1071), .o(t_2217), .co(t_2218), .cout(t_2219));
compressor_3_2 u1_784(.a(t_1049), .b(t_1046), .cin(t_1043), .o(t_2220), .cout(t_2221));
compressor_4_2 u2_785(.a(t_1083), .b(t_1080), .c(t_1077), .d(t_2213), .cin(t_2216), .o(t_2222), .co(t_2223), .cout(t_2224));
compressor_4_2 u2_786(.a(t_1092), .b(t_1089), .c(t_1086), .d(t_2219), .cin(t_2221), .o(t_2225), .co(t_2226), .cout(t_2227));
compressor_4_2 u2_787(.a(t_1066), .b(t_1063), .c(t_1060), .d(t_1057), .cin(t_1095), .o(t_2228), .co(t_2229), .cout(t_2230));
compressor_3_2 u1_788(.a(t_1075), .b(t_1072), .cin(t_1069), .o(t_2231), .cout(t_2232));
compressor_4_2 u2_789(.a(t_1101), .b(t_1098), .c(s_76_26), .d(t_2224), .cin(t_2227), .o(t_2233), .co(t_2234), .cout(t_2235));
compressor_4_2 u2_790(.a(t_1110), .b(t_1107), .c(t_1104), .d(t_2230), .cin(t_2232), .o(t_2236), .co(t_2237), .cout(t_2238));
compressor_4_2 u2_791(.a(t_1084), .b(t_1081), .c(t_1078), .d(t_1116), .cin(t_1113), .o(t_2239), .co(t_2240), .cout(t_2241));
compressor_3_2 u1_792(.a(t_1093), .b(t_1090), .cin(t_1087), .o(t_2242), .cout(t_2243));
compressor_4_2 u2_793(.a(t_1121), .b(t_1118), .c(s_77_26), .d(t_2235), .cin(t_2238), .o(t_2244), .co(t_2245), .cout(t_2246));
compressor_4_2 u2_794(.a(t_1130), .b(t_1127), .c(t_1124), .d(t_2241), .cin(t_2243), .o(t_2247), .co(t_2248), .cout(t_2249));
compressor_4_2 u2_795(.a(t_1105), .b(t_1102), .c(t_1099), .d(t_1136), .cin(t_1133), .o(t_2250), .co(t_2251), .cout(t_2252));
compressor_3_2 u1_796(.a(t_1114), .b(t_1111), .cin(t_1108), .o(t_2253), .cout(t_2254));
compressor_4_2 u2_797(.a(t_1144), .b(t_1141), .c(t_1138), .d(t_2246), .cin(t_2249), .o(t_2255), .co(t_2256), .cout(t_2257));
compressor_4_2 u2_798(.a(t_1153), .b(t_1150), .c(t_1147), .d(t_2252), .cin(t_2254), .o(t_2258), .co(t_2259), .cout(t_2260));
compressor_4_2 u2_799(.a(t_1128), .b(t_1125), .c(t_1122), .d(t_1119), .cin(t_1156), .o(t_2261), .co(t_2262), .cout(t_2263));
half_adder u0_800(.a(t_1134), .b(t_1131), .o(t_2264), .cout(t_2265));
compressor_4_2 u2_801(.a(t_1164), .b(t_1161), .c(t_1158), .d(t_2257), .cin(t_2260), .o(t_2266), .co(t_2267), .cout(t_2268));
compressor_4_2 u2_802(.a(t_1173), .b(t_1170), .c(t_1167), .d(t_2263), .cin(t_2265), .o(t_2269), .co(t_2270), .cout(t_2271));
compressor_4_2 u2_803(.a(t_1148), .b(t_1145), .c(t_1142), .d(t_1139), .cin(t_1176), .o(t_2272), .co(t_2273), .cout(t_2274));
half_adder u0_804(.a(t_1154), .b(t_1151), .o(t_2275), .cout(t_2276));
compressor_4_2 u2_805(.a(t_1184), .b(t_1181), .c(t_1178), .d(t_2268), .cin(t_2271), .o(t_2277), .co(t_2278), .cout(t_2279));
compressor_4_2 u2_806(.a(t_1193), .b(t_1190), .c(t_1187), .d(t_2274), .cin(t_2276), .o(t_2280), .co(t_2281), .cout(t_2282));
compressor_4_2 u2_807(.a(t_1168), .b(t_1165), .c(t_1162), .d(t_1159), .cin(t_1196), .o(t_2283), .co(t_2284), .cout(t_2285));
half_adder u0_808(.a(t_1174), .b(t_1171), .o(t_2286), .cout(t_2287));
compressor_4_2 u2_809(.a(t_1204), .b(t_1201), .c(t_1198), .d(t_2279), .cin(t_2282), .o(t_2288), .co(t_2289), .cout(t_2290));
compressor_4_2 u2_810(.a(t_1213), .b(t_1210), .c(t_1207), .d(t_2285), .cin(t_2287), .o(t_2291), .co(t_2292), .cout(t_2293));
compressor_4_2 u2_811(.a(t_1188), .b(t_1185), .c(t_1182), .d(t_1179), .cin(t_1216), .o(t_2294), .co(t_2295), .cout(t_2296));
half_adder u0_812(.a(t_1194), .b(t_1191), .o(t_2297), .cout(t_2298));
compressor_4_2 u2_813(.a(t_1221), .b(t_1218), .c(s_82_23), .d(t_2290), .cin(t_2293), .o(t_2299), .co(t_2300), .cout(t_2301));
compressor_4_2 u2_814(.a(t_1230), .b(t_1227), .c(t_1224), .d(t_2296), .cin(t_2298), .o(t_2302), .co(t_2303), .cout(t_2304));
compressor_4_2 u2_815(.a(t_1208), .b(t_1205), .c(t_1202), .d(t_1199), .cin(t_1233), .o(t_2305), .co(t_2306), .cout(t_2307));
half_adder u0_816(.a(t_1214), .b(t_1211), .o(t_2308), .cout(t_2309));
compressor_4_2 u2_817(.a(t_1242), .b(t_1239), .c(t_1236), .d(t_2301), .cin(t_2304), .o(t_2310), .co(t_2311), .cout(t_2312));
compressor_4_2 u2_818(.a(t_1251), .b(t_1248), .c(t_1245), .d(t_2307), .cin(t_2309), .o(t_2313), .co(t_2314), .cout(t_2315));
compressor_4_2 u2_819(.a(t_1231), .b(t_1228), .c(t_1225), .d(t_1222), .cin(t_1219), .o(t_2316), .co(t_2317), .cout(t_2318));
compressor_4_2 u2_820(.a(t_1257), .b(t_1254), .c(s_84_22), .d(t_2312), .cin(t_2315), .o(t_2319), .co(t_2320), .cout(t_2321));
compressor_4_2 u2_821(.a(t_1269), .b(t_1266), .c(t_1263), .d(t_1260), .cin(t_2318), .o(t_2322), .co(t_2323), .cout(t_2324));
compressor_4_2 u2_822(.a(t_1249), .b(t_1246), .c(t_1243), .d(t_1240), .cin(t_1237), .o(t_2325), .co(t_2326), .cout(t_2327));
compressor_4_2 u2_823(.a(t_1274), .b(t_1271), .c(s_85_22), .d(t_2321), .cin(t_2324), .o(t_2328), .co(t_2329), .cout(t_2330));
compressor_4_2 u2_824(.a(t_1286), .b(t_1283), .c(t_1280), .d(t_1277), .cin(t_2327), .o(t_2331), .co(t_2332), .cout(t_2333));
compressor_4_2 u2_825(.a(t_1267), .b(t_1264), .c(t_1261), .d(t_1258), .cin(t_1255), .o(t_2334), .co(t_2335), .cout(t_2336));
compressor_4_2 u2_826(.a(t_1294), .b(t_1291), .c(t_1288), .d(t_2330), .cin(t_2333), .o(t_2337), .co(t_2338), .cout(t_2339));
compressor_4_2 u2_827(.a(t_1272), .b(t_1303), .c(t_1300), .d(t_1297), .cin(t_2336), .o(t_2340), .co(t_2341), .cout(t_2342));
compressor_3_2 u1_828(.a(t_1281), .b(t_1278), .cin(t_1275), .o(t_2343), .cout(t_2344));
compressor_4_2 u2_829(.a(t_1311), .b(t_1308), .c(t_1305), .d(t_2339), .cin(t_2342), .o(t_2345), .co(t_2346), .cout(t_2347));
compressor_4_2 u2_830(.a(t_1289), .b(t_1320), .c(t_1317), .d(t_1314), .cin(t_2344), .o(t_2348), .co(t_2349), .cout(t_2350));
compressor_3_2 u1_831(.a(t_1298), .b(t_1295), .cin(t_1292), .o(t_2351), .cout(t_2352));
compressor_4_2 u2_832(.a(t_1328), .b(t_1325), .c(t_1322), .d(t_2347), .cin(t_2350), .o(t_2353), .co(t_2354), .cout(t_2355));
compressor_4_2 u2_833(.a(t_1306), .b(t_1337), .c(t_1334), .d(t_1331), .cin(t_2352), .o(t_2356), .co(t_2357), .cout(t_2358));
compressor_3_2 u1_834(.a(t_1315), .b(t_1312), .cin(t_1309), .o(t_2359), .cout(t_2360));
compressor_4_2 u2_835(.a(t_1345), .b(t_1342), .c(t_1339), .d(t_2355), .cin(t_2358), .o(t_2361), .co(t_2362), .cout(t_2363));
compressor_4_2 u2_836(.a(t_1323), .b(t_1354), .c(t_1351), .d(t_1348), .cin(t_2360), .o(t_2364), .co(t_2365), .cout(t_2366));
compressor_3_2 u1_837(.a(t_1332), .b(t_1329), .cin(t_1326), .o(t_2367), .cout(t_2368));
compressor_4_2 u2_838(.a(t_1359), .b(t_1356), .c(s_90_19), .d(t_2363), .cin(t_2366), .o(t_2369), .co(t_2370), .cout(t_2371));
compressor_4_2 u2_839(.a(t_1340), .b(t_1368), .c(t_1365), .d(t_1362), .cin(t_2368), .o(t_2372), .co(t_2373), .cout(t_2374));
compressor_3_2 u1_840(.a(t_1349), .b(t_1346), .cin(t_1343), .o(t_2375), .cout(t_2376));
compressor_4_2 u2_841(.a(t_1377), .b(t_1374), .c(t_1371), .d(t_2371), .cin(t_2374), .o(t_2377), .co(t_2378), .cout(t_2379));
compressor_4_2 u2_842(.a(t_1360), .b(t_1357), .c(t_1383), .d(t_1380), .cin(t_2376), .o(t_2380), .co(t_2381), .cout(t_2382));
compressor_3_2 u1_843(.a(t_1369), .b(t_1366), .cin(t_1363), .o(t_2383), .cout(t_2384));
compressor_4_2 u2_844(.a(t_1389), .b(t_1386), .c(s_92_18), .d(t_2379), .cin(t_2382), .o(t_2385), .co(t_2386), .cout(t_2387));
compressor_4_2 u2_845(.a(t_1372), .b(t_1398), .c(t_1395), .d(t_1392), .cin(t_2384), .o(t_2388), .co(t_2389), .cout(t_2390));
compressor_3_2 u1_846(.a(t_1381), .b(t_1378), .cin(t_1375), .o(t_2391), .cout(t_2392));
compressor_4_2 u2_847(.a(t_1403), .b(t_1400), .c(s_93_18), .d(t_2387), .cin(t_2390), .o(t_2393), .co(t_2394), .cout(t_2395));
compressor_4_2 u2_848(.a(t_1387), .b(t_1412), .c(t_1409), .d(t_1406), .cin(t_2392), .o(t_2396), .co(t_2397), .cout(t_2398));
compressor_3_2 u1_849(.a(t_1396), .b(t_1393), .cin(t_1390), .o(t_2399), .cout(t_2400));
compressor_4_2 u2_850(.a(t_1420), .b(t_1417), .c(t_1414), .d(t_2395), .cin(t_2398), .o(t_2401), .co(t_2402), .cout(t_2403));
compressor_4_2 u2_851(.a(t_1404), .b(t_1401), .c(t_1426), .d(t_1423), .cin(t_2400), .o(t_2404), .co(t_2405), .cout(t_2406));
half_adder u0_852(.a(t_1410), .b(t_1407), .o(t_2407), .cout(t_2408));
compressor_4_2 u2_853(.a(t_1434), .b(t_1431), .c(t_1428), .d(t_2403), .cin(t_2406), .o(t_2409), .co(t_2410), .cout(t_2411));
compressor_4_2 u2_854(.a(t_1418), .b(t_1415), .c(t_1440), .d(t_1437), .cin(t_2408), .o(t_2412), .co(t_2413), .cout(t_2414));
half_adder u0_855(.a(t_1424), .b(t_1421), .o(t_2415), .cout(t_2416));
compressor_4_2 u2_856(.a(t_1448), .b(t_1445), .c(t_1442), .d(t_2411), .cin(t_2414), .o(t_2417), .co(t_2418), .cout(t_2419));
compressor_4_2 u2_857(.a(t_1432), .b(t_1429), .c(t_1454), .d(t_1451), .cin(t_2416), .o(t_2420), .co(t_2421), .cout(t_2422));
half_adder u0_858(.a(t_1438), .b(t_1435), .o(t_2423), .cout(t_2424));
compressor_4_2 u2_859(.a(t_1462), .b(t_1459), .c(t_1456), .d(t_2419), .cin(t_2422), .o(t_2425), .co(t_2426), .cout(t_2427));
compressor_4_2 u2_860(.a(t_1446), .b(t_1443), .c(t_1468), .d(t_1465), .cin(t_2424), .o(t_2428), .co(t_2429), .cout(t_2430));
half_adder u0_861(.a(t_1452), .b(t_1449), .o(t_2431), .cout(t_2432));
compressor_4_2 u2_862(.a(t_1473), .b(t_1470), .c(s_98_15), .d(t_2427), .cin(t_2430), .o(t_2433), .co(t_2434), .cout(t_2435));
compressor_4_2 u2_863(.a(t_1460), .b(t_1457), .c(t_1479), .d(t_1476), .cin(t_2432), .o(t_2436), .co(t_2437), .cout(t_2438));
half_adder u0_864(.a(t_1466), .b(t_1463), .o(t_2439), .cout(t_2440));
compressor_4_2 u2_865(.a(t_1488), .b(t_1485), .c(t_1482), .d(t_2435), .cin(t_2438), .o(t_2441), .co(t_2442), .cout(t_2443));
compressor_4_2 u2_866(.a(t_1477), .b(t_1474), .c(t_1471), .d(t_1491), .cin(t_2440), .o(t_2444), .co(t_2445), .cout(t_2446));
compressor_4_2 u2_867(.a(t_1497), .b(t_1494), .c(s_100_14), .d(t_2443), .cin(t_2446), .o(t_2447), .co(t_2448), .cout(t_2449));
compressor_4_2 u2_868(.a(t_1489), .b(t_1486), .c(t_1483), .d(t_1503), .cin(t_1500), .o(t_2450), .co(t_2451), .cout(t_2452));
compressor_4_2 u2_869(.a(t_1508), .b(t_1505), .c(s_101_14), .d(t_2449), .cin(t_2452), .o(t_2453), .co(t_2454), .cout(t_2455));
compressor_4_2 u2_870(.a(t_1501), .b(t_1498), .c(t_1495), .d(t_1514), .cin(t_1511), .o(t_2456), .co(t_2457), .cout(t_2458));
compressor_4_2 u2_871(.a(t_1522), .b(t_1519), .c(t_1516), .d(t_2455), .cin(t_2458), .o(t_2459), .co(t_2460), .cout(t_2461));
compressor_3_2 u1_872(.a(t_1509), .b(t_1506), .cin(t_1525), .o(t_2462), .cout(t_2463));
compressor_4_2 u2_873(.a(t_1533), .b(t_1530), .c(t_1527), .d(t_2461), .cin(t_2463), .o(t_2464), .co(t_2465), .cout(t_2466));
compressor_3_2 u1_874(.a(t_1520), .b(t_1517), .cin(t_1536), .o(t_2467), .cout(t_2468));
compressor_4_2 u2_875(.a(t_1544), .b(t_1541), .c(t_1538), .d(t_2466), .cin(t_2468), .o(t_2469), .co(t_2470), .cout(t_2471));
compressor_3_2 u1_876(.a(t_1531), .b(t_1528), .cin(t_1547), .o(t_2472), .cout(t_2473));
compressor_4_2 u2_877(.a(t_1555), .b(t_1552), .c(t_1549), .d(t_2471), .cin(t_2473), .o(t_2474), .co(t_2475), .cout(t_2476));
compressor_3_2 u1_878(.a(t_1542), .b(t_1539), .cin(t_1558), .o(t_2477), .cout(t_2478));
compressor_4_2 u2_879(.a(t_1563), .b(t_1560), .c(s_106_11), .d(t_2476), .cin(t_2478), .o(t_2479), .co(t_2480), .cout(t_2481));
compressor_3_2 u1_880(.a(t_1553), .b(t_1550), .cin(t_1566), .o(t_2482), .cout(t_2483));
compressor_4_2 u2_881(.a(t_1575), .b(t_1572), .c(t_1569), .d(t_2481), .cin(t_2483), .o(t_2484), .co(t_2485), .cout(t_2486));
compressor_3_2 u1_882(.a(t_1567), .b(t_1564), .cin(t_1561), .o(t_2487), .cout(t_2488));
compressor_4_2 u2_883(.a(t_1581), .b(t_1578), .c(s_108_10), .d(t_2486), .cin(t_2488), .o(t_2489), .co(t_2490), .cout(t_2491));
compressor_3_2 u1_884(.a(t_1573), .b(t_1570), .cin(t_1584), .o(t_2492), .cout(t_2493));
compressor_4_2 u2_885(.a(t_1589), .b(t_1586), .c(s_109_10), .d(t_2491), .cin(t_2493), .o(t_2494), .co(t_2495), .cout(t_2496));
compressor_3_2 u1_886(.a(t_1582), .b(t_1579), .cin(t_1592), .o(t_2497), .cout(t_2498));
compressor_4_2 u2_887(.a(t_1600), .b(t_1597), .c(t_1594), .d(t_2496), .cin(t_2498), .o(t_2499), .co(t_2500), .cout(t_2501));
half_adder u0_888(.a(t_1590), .b(t_1587), .o(t_2502), .cout(t_2503));
compressor_4_2 u2_889(.a(t_1608), .b(t_1605), .c(t_1602), .d(t_2501), .cin(t_2503), .o(t_2504), .co(t_2505), .cout(t_2506));
half_adder u0_890(.a(t_1598), .b(t_1595), .o(t_2507), .cout(t_2508));
compressor_4_2 u2_891(.a(t_1616), .b(t_1613), .c(t_1610), .d(t_2506), .cin(t_2508), .o(t_2509), .co(t_2510), .cout(t_2511));
half_adder u0_892(.a(t_1606), .b(t_1603), .o(t_2512), .cout(t_2513));
compressor_4_2 u2_893(.a(t_1624), .b(t_1621), .c(t_1618), .d(t_2511), .cin(t_2513), .o(t_2514), .co(t_2515), .cout(t_2516));
half_adder u0_894(.a(t_1614), .b(t_1611), .o(t_2517), .cout(t_2518));
compressor_4_2 u2_895(.a(t_1629), .b(t_1626), .c(s_114_7), .d(t_2516), .cin(t_2518), .o(t_2519), .co(t_2520), .cout(t_2521));
half_adder u0_896(.a(t_1622), .b(t_1619), .o(t_2522), .cout(t_2523));
compressor_4_2 u2_897(.a(t_1627), .b(t_1635), .c(t_1632), .d(t_2521), .cin(t_2523), .o(t_2524), .co(t_2525), .cout(t_2526));
compressor_4_2 u2_898(.a(t_1633), .b(t_1641), .c(t_1638), .d(s_116_6), .cin(t_2526), .o(t_2527), .co(t_2528), .cout(t_2529));
compressor_4_2 u2_899(.a(t_1639), .b(t_1646), .c(t_1643), .d(s_117_6), .cin(t_2529), .o(t_2530), .co(t_2531), .cout(t_2532));
compressor_3_2 u1_900(.a(t_1651), .b(t_1648), .cin(t_2532), .o(t_2533), .cout(t_2534));
compressor_3_2 u1_901(.a(t_1649), .b(t_1656), .cin(t_1653), .o(t_2535), .cout(t_2536));
compressor_3_2 u1_902(.a(t_1654), .b(t_1661), .cin(t_1658), .o(t_2537), .cout(t_2538));
compressor_3_2 u1_903(.a(t_1659), .b(t_1666), .cin(t_1663), .o(t_2539), .cout(t_2540));
compressor_3_2 u1_904(.a(t_1664), .b(t_1668), .cin(s_122_3), .o(t_2541), .cout(t_2542));
half_adder u0_905(.a(t_1669), .b(t_1671), .o(t_2543), .cout(t_2544));
compressor_3_2 u1_906(.a(t_1672), .b(t_1674), .cin(s_124_2), .o(t_2545), .cout(t_2546));
half_adder u0_907(.a(t_1675), .b(t_1676), .o(t_2547), .cout(t_2548));
half_adder u0_908(.a(t_1677), .b(t_1678), .o(t_2549), .cout(t_2550));
half_adder u0_909(.a(t_1679), .b(t_1680), .o(t_2551), .cout());

/* u0_910 Output nets */
wire t_2552,   t_2553;
/* u0_911 Output nets */
wire t_2554,   t_2555;
/* u0_912 Output nets */
wire t_2556,   t_2557;
/* u0_913 Output nets */
wire t_2558,   t_2559;
/* u0_914 Output nets */
wire t_2560,   t_2561;
/* u0_915 Output nets */
wire t_2562,   t_2563;
/* u1_916 Output nets */
wire t_2564,   t_2565;
/* u0_917 Output nets */
wire t_2566,   t_2567;
/* u0_918 Output nets */
wire t_2568,   t_2569;
/* u0_919 Output nets */
wire t_2570,   t_2571;
/* u0_920 Output nets */
wire t_2572,   t_2573;
/* u1_921 Output nets */
wire t_2574,   t_2575;
/* u1_922 Output nets */
wire t_2576,   t_2577;
/* u1_923 Output nets */
wire t_2578,   t_2579;
/* u1_924 Output nets */
wire t_2580,   t_2581;
/* u1_925 Output nets */
wire t_2582,   t_2583;
/* u2_926 Output nets */
wire t_2584,   t_2585,   t_2586;
/* u1_927 Output nets */
wire t_2587,   t_2588;
/* u1_928 Output nets */
wire t_2589,   t_2590;
/* u2_929 Output nets */
wire t_2591,   t_2592,   t_2593;
/* u2_930 Output nets */
wire t_2594,   t_2595,   t_2596;
/* u1_931 Output nets */
wire t_2597,   t_2598;
/* u2_932 Output nets */
wire t_2599,   t_2600,   t_2601;
/* u2_933 Output nets */
wire t_2602,   t_2603,   t_2604;
/* u2_934 Output nets */
wire t_2605,   t_2606,   t_2607;
/* u2_935 Output nets */
wire t_2608,   t_2609,   t_2610;
/* u2_936 Output nets */
wire t_2611,   t_2612,   t_2613;
/* u2_937 Output nets */
wire t_2614,   t_2615,   t_2616;
/* u2_938 Output nets */
wire t_2617,   t_2618,   t_2619;
/* u2_939 Output nets */
wire t_2620,   t_2621,   t_2622;
/* u2_940 Output nets */
wire t_2623,   t_2624,   t_2625;
/* u2_941 Output nets */
wire t_2626,   t_2627,   t_2628;
/* u2_942 Output nets */
wire t_2629,   t_2630,   t_2631;
/* u0_943 Output nets */
wire t_2632,   t_2633;
/* u2_944 Output nets */
wire t_2634,   t_2635,   t_2636;
/* u0_945 Output nets */
wire t_2637,   t_2638;
/* u2_946 Output nets */
wire t_2639,   t_2640,   t_2641;
/* u0_947 Output nets */
wire t_2642,   t_2643;
/* u2_948 Output nets */
wire t_2644,   t_2645,   t_2646;
/* u1_949 Output nets */
wire t_2647,   t_2648;
/* u2_950 Output nets */
wire t_2649,   t_2650,   t_2651;
/* u1_951 Output nets */
wire t_2652,   t_2653;
/* u2_952 Output nets */
wire t_2654,   t_2655,   t_2656;
/* u0_953 Output nets */
wire t_2657,   t_2658;
/* u2_954 Output nets */
wire t_2659,   t_2660,   t_2661;
/* u1_955 Output nets */
wire t_2662,   t_2663;
/* u2_956 Output nets */
wire t_2664,   t_2665,   t_2666;
/* u1_957 Output nets */
wire t_2667,   t_2668;
/* u2_958 Output nets */
wire t_2669,   t_2670,   t_2671;
/* u1_959 Output nets */
wire t_2672,   t_2673;
/* u2_960 Output nets */
wire t_2674,   t_2675,   t_2676;
/* u1_961 Output nets */
wire t_2677,   t_2678;
/* u2_962 Output nets */
wire t_2679,   t_2680,   t_2681;
/* u1_963 Output nets */
wire t_2682,   t_2683;
/* u2_964 Output nets */
wire t_2684,   t_2685,   t_2686;
/* u1_965 Output nets */
wire t_2687,   t_2688;
/* u2_966 Output nets */
wire t_2689,   t_2690,   t_2691;
/* u1_967 Output nets */
wire t_2692,   t_2693;
/* u2_968 Output nets */
wire t_2694,   t_2695,   t_2696;
/* u1_969 Output nets */
wire t_2697,   t_2698;
/* u2_970 Output nets */
wire t_2699,   t_2700,   t_2701;
/* u1_971 Output nets */
wire t_2702,   t_2703;
/* u2_972 Output nets */
wire t_2704,   t_2705,   t_2706;
/* u1_973 Output nets */
wire t_2707,   t_2708;
/* u2_974 Output nets */
wire t_2709,   t_2710,   t_2711;
/* u2_975 Output nets */
wire t_2712,   t_2713,   t_2714;
/* u2_976 Output nets */
wire t_2715,   t_2716,   t_2717;
/* u1_977 Output nets */
wire t_2718,   t_2719;
/* u2_978 Output nets */
wire t_2720,   t_2721,   t_2722;
/* u1_979 Output nets */
wire t_2723,   t_2724;
/* u2_980 Output nets */
wire t_2725,   t_2726,   t_2727;
/* u2_981 Output nets */
wire t_2728,   t_2729,   t_2730;
/* u2_982 Output nets */
wire t_2731,   t_2732,   t_2733;
/* u2_983 Output nets */
wire t_2734,   t_2735,   t_2736;
/* u2_984 Output nets */
wire t_2737,   t_2738,   t_2739;
/* u1_985 Output nets */
wire t_2740,   t_2741;
/* u2_986 Output nets */
wire t_2742,   t_2743,   t_2744;
/* u2_987 Output nets */
wire t_2745,   t_2746,   t_2747;
/* u2_988 Output nets */
wire t_2748,   t_2749,   t_2750;
/* u2_989 Output nets */
wire t_2751,   t_2752,   t_2753;
/* u2_990 Output nets */
wire t_2754,   t_2755,   t_2756;
/* u2_991 Output nets */
wire t_2757,   t_2758,   t_2759;
/* u2_992 Output nets */
wire t_2760,   t_2761,   t_2762;
/* u2_993 Output nets */
wire t_2763,   t_2764,   t_2765;
/* u2_994 Output nets */
wire t_2766,   t_2767,   t_2768;
/* u2_995 Output nets */
wire t_2769,   t_2770,   t_2771;
/* u2_996 Output nets */
wire t_2772,   t_2773,   t_2774;
/* u2_997 Output nets */
wire t_2775,   t_2776,   t_2777;
/* u2_998 Output nets */
wire t_2778,   t_2779,   t_2780;
/* u2_999 Output nets */
wire t_2781,   t_2782,   t_2783;
/* u2_1000 Output nets */
wire t_2784,   t_2785,   t_2786;
/* u2_1001 Output nets */
wire t_2787,   t_2788,   t_2789;
/* u2_1002 Output nets */
wire t_2790,   t_2791,   t_2792;
/* u2_1003 Output nets */
wire t_2793,   t_2794,   t_2795;
/* u2_1004 Output nets */
wire t_2796,   t_2797,   t_2798;
/* u2_1005 Output nets */
wire t_2799,   t_2800,   t_2801;
/* u2_1006 Output nets */
wire t_2802,   t_2803,   t_2804;
/* u2_1007 Output nets */
wire t_2805,   t_2806,   t_2807;
/* u2_1008 Output nets */
wire t_2808,   t_2809,   t_2810;
/* u2_1009 Output nets */
wire t_2811,   t_2812,   t_2813;
/* u2_1010 Output nets */
wire t_2814,   t_2815,   t_2816;
/* u2_1011 Output nets */
wire t_2817,   t_2818,   t_2819;
/* u2_1012 Output nets */
wire t_2820,   t_2821,   t_2822;
/* u2_1013 Output nets */
wire t_2823,   t_2824,   t_2825;
/* u2_1014 Output nets */
wire t_2826,   t_2827,   t_2828;
/* u2_1015 Output nets */
wire t_2829,   t_2830,   t_2831;
/* u2_1016 Output nets */
wire t_2832,   t_2833,   t_2834;
/* u2_1017 Output nets */
wire t_2835,   t_2836,   t_2837;
/* u2_1018 Output nets */
wire t_2838,   t_2839,   t_2840;
/* u1_1019 Output nets */
wire t_2841,   t_2842;
/* u2_1020 Output nets */
wire t_2843,   t_2844,   t_2845;
/* u2_1021 Output nets */
wire t_2846,   t_2847,   t_2848;
/* u2_1022 Output nets */
wire t_2849,   t_2850,   t_2851;
/* u1_1023 Output nets */
wire t_2852,   t_2853;
/* u2_1024 Output nets */
wire t_2854,   t_2855,   t_2856;
/* u1_1025 Output nets */
wire t_2857,   t_2858;
/* u2_1026 Output nets */
wire t_2859,   t_2860,   t_2861;
/* u1_1027 Output nets */
wire t_2862,   t_2863;
/* u2_1028 Output nets */
wire t_2864,   t_2865,   t_2866;
/* u1_1029 Output nets */
wire t_2867,   t_2868;
/* u2_1030 Output nets */
wire t_2869,   t_2870,   t_2871;
/* u1_1031 Output nets */
wire t_2872,   t_2873;
/* u2_1032 Output nets */
wire t_2874,   t_2875,   t_2876;
/* u1_1033 Output nets */
wire t_2877,   t_2878;
/* u2_1034 Output nets */
wire t_2879,   t_2880,   t_2881;
/* u1_1035 Output nets */
wire t_2882,   t_2883;
/* u2_1036 Output nets */
wire t_2884,   t_2885,   t_2886;
/* u1_1037 Output nets */
wire t_2887,   t_2888;
/* u2_1038 Output nets */
wire t_2889,   t_2890,   t_2891;
/* u1_1039 Output nets */
wire t_2892,   t_2893;
/* u2_1040 Output nets */
wire t_2894,   t_2895,   t_2896;
/* u1_1041 Output nets */
wire t_2897,   t_2898;
/* u2_1042 Output nets */
wire t_2899,   t_2900,   t_2901;
/* u1_1043 Output nets */
wire t_2902,   t_2903;
/* u2_1044 Output nets */
wire t_2904,   t_2905,   t_2906;
/* u1_1045 Output nets */
wire t_2907,   t_2908;
/* u2_1046 Output nets */
wire t_2909,   t_2910,   t_2911;
/* u1_1047 Output nets */
wire t_2912,   t_2913;
/* u2_1048 Output nets */
wire t_2914,   t_2915,   t_2916;
/* u1_1049 Output nets */
wire t_2917,   t_2918;
/* u2_1050 Output nets */
wire t_2919,   t_2920,   t_2921;
/* u0_1051 Output nets */
wire t_2922,   t_2923;
/* u2_1052 Output nets */
wire t_2924,   t_2925,   t_2926;
/* u1_1053 Output nets */
wire t_2927,   t_2928;
/* u2_1054 Output nets */
wire t_2929,   t_2930,   t_2931;
/* u0_1055 Output nets */
wire t_2932,   t_2933;
/* u2_1056 Output nets */
wire t_2934,   t_2935,   t_2936;
/* u0_1057 Output nets */
wire t_2937,   t_2938;
/* u2_1058 Output nets */
wire t_2939,   t_2940,   t_2941;
/* u0_1059 Output nets */
wire t_2942,   t_2943;
/* u2_1060 Output nets */
wire t_2944,   t_2945,   t_2946;
/* u0_1061 Output nets */
wire t_2947,   t_2948;
/* u2_1062 Output nets */
wire t_2949,   t_2950,   t_2951;
/* u0_1063 Output nets */
wire t_2952,   t_2953;
/* u2_1064 Output nets */
wire t_2954,   t_2955,   t_2956;
/* u0_1065 Output nets */
wire t_2957,   t_2958;
/* u2_1066 Output nets */
wire t_2959,   t_2960,   t_2961;
/* u0_1067 Output nets */
wire t_2962,   t_2963;
/* u2_1068 Output nets */
wire t_2964,   t_2965,   t_2966;
/* u0_1069 Output nets */
wire t_2967,   t_2968;
/* u2_1070 Output nets */
wire t_2969,   t_2970,   t_2971;
/* u2_1071 Output nets */
wire t_2972,   t_2973,   t_2974;
/* u2_1072 Output nets */
wire t_2975,   t_2976,   t_2977;
/* u2_1073 Output nets */
wire t_2978,   t_2979,   t_2980;
/* u2_1074 Output nets */
wire t_2981,   t_2982,   t_2983;
/* u2_1075 Output nets */
wire t_2984,   t_2985,   t_2986;
/* u1_1076 Output nets */
wire t_2987,   t_2988;
/* u1_1077 Output nets */
wire t_2989,   t_2990;
/* u1_1078 Output nets */
wire t_2991,   t_2992;
/* u1_1079 Output nets */
wire t_2993,   t_2994;
/* u1_1080 Output nets */
wire t_2995,   t_2996;
/* u1_1081 Output nets */
wire t_2997,   t_2998;
/* u1_1082 Output nets */
wire t_2999,   t_3000;
/* u1_1083 Output nets */
wire t_3001,   t_3002;
/* u1_1084 Output nets */
wire t_3003,   t_3004;
/* u1_1085 Output nets */
wire t_3005,   t_3006;
/* u0_1086 Output nets */
wire t_3007,   t_3008;
/* u1_1087 Output nets */
wire t_3009,   t_3010;
/* u0_1088 Output nets */
wire t_3011,   t_3012;
/* u0_1089 Output nets */
wire t_3013,   t_3014;
/* u0_1090 Output nets */
wire t_3015,   t_3016;
/* u0_1091 Output nets */
wire t_3017,   t_3018;
/* u0_1092 Output nets */
wire t_3019,   t_3020;
/* u0_1093 Output nets */
wire t_3021,   t_3022;
/* u0_1094 Output nets */
wire t_3023,   t_3024;
/* u0_1095 Output nets */
wire t_3025,   t_3026;
/* u0_1096 Output nets */
wire t_3027;

/* compress stage 3 */
half_adder u0_910(.a(t_1682), .b(t_2), .o(t_2552), .cout(t_2553));
half_adder u0_911(.a(t_1684), .b(t_6), .o(t_2554), .cout(t_2555));
half_adder u0_912(.a(t_1686), .b(t_1687), .o(t_2556), .cout(t_2557));
half_adder u0_913(.a(t_1688), .b(t_1689), .o(t_2558), .cout(t_2559));
half_adder u0_914(.a(t_1690), .b(t_1691), .o(t_2560), .cout(t_2561));
half_adder u0_915(.a(t_1692), .b(t_1693), .o(t_2562), .cout(t_2563));
compressor_3_2 u1_916(.a(t_1696), .b(t_1698), .cin(t_28), .o(t_2564), .cout(t_2565));
half_adder u0_917(.a(t_1699), .b(t_1700), .o(t_2566), .cout(t_2567));
half_adder u0_918(.a(t_1702), .b(t_41), .o(t_2568), .cout(t_2569));
half_adder u0_919(.a(t_1703), .b(t_1705), .o(t_2570), .cout(t_2571));
half_adder u0_920(.a(t_1706), .b(t_1708), .o(t_2572), .cout(t_2573));
compressor_3_2 u1_921(.a(t_1709), .b(t_1711), .cin(t_58), .o(t_2574), .cout(t_2575));
compressor_3_2 u1_922(.a(t_1712), .b(t_1714), .cin(t_64), .o(t_2576), .cout(t_2577));
compressor_3_2 u1_923(.a(t_1715), .b(t_1720), .cin(t_1717), .o(t_2578), .cout(t_2579));
compressor_3_2 u1_924(.a(t_1718), .b(t_1725), .cin(t_1722), .o(t_2580), .cout(t_2581));
compressor_3_2 u1_925(.a(t_1723), .b(t_1730), .cin(t_1727), .o(t_2582), .cout(t_2583));
compressor_4_2 u2_926(.a(t_1728), .b(t_1735), .c(t_1732), .d(t_99), .cin(t_2583), .o(t_2584), .co(t_2585), .cout(t_2586));
compressor_3_2 u1_927(.a(t_1740), .b(t_1737), .cin(t_2586), .o(t_2587), .cout(t_2588));
compressor_3_2 u1_928(.a(t_1738), .b(t_1745), .cin(t_1742), .o(t_2589), .cout(t_2590));
compressor_4_2 u2_929(.a(t_1743), .b(t_1750), .c(t_1747), .d(t_125), .cin(t_2590), .o(t_2591), .co(t_2592), .cout(t_2593));
compressor_4_2 u2_930(.a(t_1748), .b(t_1755), .c(t_1752), .d(t_134), .cin(t_2593), .o(t_2594), .co(t_2595), .cout(t_2596));
compressor_3_2 u1_931(.a(t_1760), .b(t_1757), .cin(t_2596), .o(t_2597), .cout(t_2598));
compressor_4_2 u2_932(.a(t_1761), .b(t_1758), .c(t_1766), .d(t_1763), .cin(t_156), .o(t_2599), .co(t_2600), .cout(t_2601));
compressor_4_2 u2_933(.a(t_1764), .b(t_1771), .c(t_1768), .d(t_167), .cin(t_2601), .o(t_2602), .co(t_2603), .cout(t_2604));
compressor_4_2 u2_934(.a(t_1769), .b(t_1776), .c(t_1773), .d(t_181), .cin(t_2604), .o(t_2605), .co(t_2606), .cout(t_2607));
compressor_4_2 u2_935(.a(t_1777), .b(t_1774), .c(t_1782), .d(t_1779), .cin(t_2607), .o(t_2608), .co(t_2609), .cout(t_2610));
compressor_4_2 u2_936(.a(t_1783), .b(t_1780), .c(t_1788), .d(t_1785), .cin(t_2610), .o(t_2611), .co(t_2612), .cout(t_2613));
compressor_4_2 u2_937(.a(t_1786), .b(t_1794), .c(t_1791), .d(t_216), .cin(t_2613), .o(t_2614), .co(t_2615), .cout(t_2616));
compressor_4_2 u2_938(.a(t_1792), .b(t_1800), .c(t_1797), .d(t_228), .cin(t_2616), .o(t_2617), .co(t_2618), .cout(t_2619));
compressor_4_2 u2_939(.a(t_1798), .b(t_1809), .c(t_1806), .d(t_1803), .cin(t_2619), .o(t_2620), .co(t_2621), .cout(t_2622));
compressor_4_2 u2_940(.a(t_1804), .b(t_1817), .c(t_1814), .d(t_1811), .cin(t_2622), .o(t_2623), .co(t_2624), .cout(t_2625));
compressor_4_2 u2_941(.a(t_1812), .b(t_1825), .c(t_1822), .d(t_1819), .cin(t_2625), .o(t_2626), .co(t_2627), .cout(t_2628));
compressor_4_2 u2_942(.a(t_1833), .b(t_1830), .c(t_1827), .d(t_287), .cin(t_2628), .o(t_2629), .co(t_2630), .cout(t_2631));
half_adder u0_943(.a(t_1823), .b(t_1820), .o(t_2632), .cout(t_2633));
compressor_4_2 u2_944(.a(t_1841), .b(t_1838), .c(t_1835), .d(t_2631), .cin(t_2633), .o(t_2634), .co(t_2635), .cout(t_2636));
half_adder u0_945(.a(t_1831), .b(t_1828), .o(t_2637), .cout(t_2638));
compressor_4_2 u2_946(.a(t_1849), .b(t_1846), .c(t_1843), .d(t_2636), .cin(t_2638), .o(t_2639), .co(t_2640), .cout(t_2641));
half_adder u0_947(.a(t_1839), .b(t_1836), .o(t_2642), .cout(t_2643));
compressor_4_2 u2_948(.a(t_1854), .b(t_1851), .c(t_331), .d(t_2641), .cin(t_2643), .o(t_2644), .co(t_2645), .cout(t_2646));
compressor_3_2 u1_949(.a(t_1847), .b(t_1844), .cin(t_1857), .o(t_2647), .cout(t_2648));
compressor_4_2 u2_950(.a(t_1862), .b(t_1859), .c(t_346), .d(t_2646), .cin(t_2648), .o(t_2649), .co(t_2650), .cout(t_2651));
compressor_3_2 u1_951(.a(t_1855), .b(t_1852), .cin(t_1865), .o(t_2652), .cout(t_2653));
compressor_4_2 u2_952(.a(t_1873), .b(t_1870), .c(t_1867), .d(t_2651), .cin(t_2653), .o(t_2654), .co(t_2655), .cout(t_2656));
half_adder u0_953(.a(t_1863), .b(t_1860), .o(t_2657), .cout(t_2658));
compressor_4_2 u2_954(.a(t_1879), .b(t_1876), .c(t_380), .d(t_2656), .cin(t_2658), .o(t_2659), .co(t_2660), .cout(t_2661));
compressor_3_2 u1_955(.a(t_1871), .b(t_1868), .cin(t_1882), .o(t_2662), .cout(t_2663));
compressor_4_2 u2_956(.a(t_1887), .b(t_1884), .c(t_397), .d(t_2661), .cin(t_2663), .o(t_2664), .co(t_2665), .cout(t_2666));
compressor_3_2 u1_957(.a(t_1880), .b(t_1877), .cin(t_1890), .o(t_2667), .cout(t_2668));
compressor_4_2 u2_958(.a(t_1895), .b(t_1892), .c(t_417), .d(t_2666), .cin(t_2668), .o(t_2669), .co(t_2670), .cout(t_2671));
compressor_3_2 u1_959(.a(t_1888), .b(t_1885), .cin(t_1898), .o(t_2672), .cout(t_2673));
compressor_4_2 u2_960(.a(t_1907), .b(t_1904), .c(t_1901), .d(t_2671), .cin(t_2673), .o(t_2674), .co(t_2675), .cout(t_2676));
compressor_3_2 u1_961(.a(t_1899), .b(t_1896), .cin(t_1893), .o(t_2677), .cout(t_2678));
compressor_4_2 u2_962(.a(t_1916), .b(t_1913), .c(t_1910), .d(t_2676), .cin(t_2678), .o(t_2679), .co(t_2680), .cout(t_2681));
compressor_3_2 u1_963(.a(t_1908), .b(t_1905), .cin(t_1902), .o(t_2682), .cout(t_2683));
compressor_4_2 u2_964(.a(t_1922), .b(t_1919), .c(t_470), .d(t_2681), .cin(t_2683), .o(t_2684), .co(t_2685), .cout(t_2686));
compressor_3_2 u1_965(.a(t_1914), .b(t_1911), .cin(t_1925), .o(t_2687), .cout(t_2688));
compressor_4_2 u2_966(.a(t_1931), .b(t_1928), .c(t_488), .d(t_2686), .cin(t_2688), .o(t_2689), .co(t_2690), .cout(t_2691));
compressor_3_2 u1_967(.a(t_1923), .b(t_1920), .cin(t_1934), .o(t_2692), .cout(t_2693));
compressor_4_2 u2_968(.a(t_1943), .b(t_1940), .c(t_1937), .d(t_2691), .cin(t_2693), .o(t_2694), .co(t_2695), .cout(t_2696));
compressor_3_2 u1_969(.a(t_1932), .b(t_1929), .cin(t_1946), .o(t_2697), .cout(t_2698));
compressor_4_2 u2_970(.a(t_1954), .b(t_1951), .c(t_1948), .d(t_2696), .cin(t_2698), .o(t_2699), .co(t_2700), .cout(t_2701));
compressor_3_2 u1_971(.a(t_1941), .b(t_1938), .cin(t_1957), .o(t_2702), .cout(t_2703));
compressor_4_2 u2_972(.a(t_1965), .b(t_1962), .c(t_1959), .d(t_2701), .cin(t_2703), .o(t_2704), .co(t_2705), .cout(t_2706));
compressor_3_2 u1_973(.a(t_1952), .b(t_1949), .cin(t_1968), .o(t_2707), .cout(t_2708));
compressor_4_2 u2_974(.a(t_1973), .b(t_1970), .c(t_571), .d(t_2706), .cin(t_2708), .o(t_2709), .co(t_2710), .cout(t_2711));
compressor_4_2 u2_975(.a(t_1966), .b(t_1963), .c(t_1960), .d(t_1979), .cin(t_1976), .o(t_2712), .co(t_2713), .cout(t_2714));
compressor_4_2 u2_976(.a(t_1987), .b(t_1984), .c(t_1981), .d(t_2711), .cin(t_2714), .o(t_2715), .co(t_2716), .cout(t_2717));
compressor_3_2 u1_977(.a(t_1974), .b(t_1971), .cin(t_1990), .o(t_2718), .cout(t_2719));
compressor_4_2 u2_978(.a(t_1998), .b(t_1995), .c(t_1992), .d(t_2717), .cin(t_2719), .o(t_2720), .co(t_2721), .cout(t_2722));
compressor_3_2 u1_979(.a(t_1985), .b(t_1982), .cin(t_2001), .o(t_2723), .cout(t_2724));
compressor_4_2 u2_980(.a(t_2006), .b(t_2003), .c(t_633), .d(t_2722), .cin(t_2724), .o(t_2725), .co(t_2726), .cout(t_2727));
compressor_4_2 u2_981(.a(t_1999), .b(t_1996), .c(t_1993), .d(t_2012), .cin(t_2009), .o(t_2728), .co(t_2729), .cout(t_2730));
compressor_4_2 u2_982(.a(t_2017), .b(t_2014), .c(t_654), .d(t_2727), .cin(t_2730), .o(t_2731), .co(t_2732), .cout(t_2733));
compressor_4_2 u2_983(.a(t_2010), .b(t_2007), .c(t_2004), .d(t_2023), .cin(t_2020), .o(t_2734), .co(t_2735), .cout(t_2736));
compressor_4_2 u2_984(.a(t_2031), .b(t_2028), .c(t_2025), .d(t_2733), .cin(t_2736), .o(t_2737), .co(t_2738), .cout(t_2739));
compressor_3_2 u1_985(.a(t_2018), .b(t_2015), .cin(t_2034), .o(t_2740), .cout(t_2741));
compressor_4_2 u2_986(.a(t_2040), .b(t_2037), .c(t_700), .d(t_2739), .cin(t_2741), .o(t_2742), .co(t_2743), .cout(t_2744));
compressor_4_2 u2_987(.a(t_2032), .b(t_2029), .c(t_2026), .d(t_2046), .cin(t_2043), .o(t_2745), .co(t_2746), .cout(t_2747));
compressor_4_2 u2_988(.a(t_2051), .b(t_2048), .c(t_723), .d(t_2744), .cin(t_2747), .o(t_2748), .co(t_2749), .cout(t_2750));
compressor_4_2 u2_989(.a(t_2044), .b(t_2041), .c(t_2038), .d(t_2057), .cin(t_2054), .o(t_2751), .co(t_2752), .cout(t_2753));
compressor_4_2 u2_990(.a(t_2062), .b(t_2059), .c(t_749), .d(t_2750), .cin(t_2753), .o(t_2754), .co(t_2755), .cout(t_2756));
compressor_4_2 u2_991(.a(t_2055), .b(t_2052), .c(t_2049), .d(t_2068), .cin(t_2065), .o(t_2757), .co(t_2758), .cout(t_2759));
compressor_4_2 u2_992(.a(t_2077), .b(t_2074), .c(t_2071), .d(t_2756), .cin(t_2759), .o(t_2760), .co(t_2761), .cout(t_2762));
compressor_4_2 u2_993(.a(t_2069), .b(t_2066), .c(t_2063), .d(t_2060), .cin(t_2080), .o(t_2763), .co(t_2764), .cout(t_2765));
compressor_4_2 u2_994(.a(t_2089), .b(t_2086), .c(t_2083), .d(t_2762), .cin(t_2765), .o(t_2766), .co(t_2767), .cout(t_2768));
compressor_4_2 u2_995(.a(t_2081), .b(t_2078), .c(t_2075), .d(t_2072), .cin(t_2092), .o(t_2769), .co(t_2770), .cout(t_2771));
compressor_4_2 u2_996(.a(t_2098), .b(t_2095), .c(t_820), .d(t_2768), .cin(t_2771), .o(t_2772), .co(t_2773), .cout(t_2774));
compressor_4_2 u2_997(.a(t_2090), .b(t_2087), .c(t_2084), .d(t_2104), .cin(t_2101), .o(t_2775), .co(t_2776), .cout(t_2777));
compressor_4_2 u2_998(.a(t_2110), .b(t_2107), .c(t_844), .d(t_2774), .cin(t_2777), .o(t_2778), .co(t_2779), .cout(t_2780));
compressor_4_2 u2_999(.a(t_2102), .b(t_2099), .c(t_2096), .d(t_2116), .cin(t_2113), .o(t_2781), .co(t_2782), .cout(t_2783));
compressor_4_2 u2_1000(.a(t_2125), .b(t_2122), .c(t_2119), .d(t_2780), .cin(t_2783), .o(t_2784), .co(t_2785), .cout(t_2786));
compressor_4_2 u2_1001(.a(t_2117), .b(t_2114), .c(t_2111), .d(t_2108), .cin(t_2128), .o(t_2787), .co(t_2788), .cout(t_2789));
compressor_4_2 u2_1002(.a(t_2137), .b(t_2134), .c(t_2131), .d(t_2786), .cin(t_2789), .o(t_2790), .co(t_2791), .cout(t_2792));
compressor_4_2 u2_1003(.a(t_2129), .b(t_2126), .c(t_2123), .d(t_2120), .cin(t_2140), .o(t_2793), .co(t_2794), .cout(t_2795));
compressor_4_2 u2_1004(.a(t_2146), .b(t_2143), .c(t_916), .d(t_2792), .cin(t_2795), .o(t_2796), .co(t_2797), .cout(t_2798));
compressor_4_2 u2_1005(.a(t_2138), .b(t_2135), .c(t_2132), .d(t_2152), .cin(t_2149), .o(t_2799), .co(t_2800), .cout(t_2801));
compressor_4_2 u2_1006(.a(t_2161), .b(t_2158), .c(t_2155), .d(t_2798), .cin(t_2801), .o(t_2802), .co(t_2803), .cout(t_2804));
compressor_4_2 u2_1007(.a(t_2153), .b(t_2150), .c(t_2147), .d(t_2144), .cin(t_2164), .o(t_2805), .co(t_2806), .cout(t_2807));
compressor_4_2 u2_1008(.a(t_2170), .b(t_2167), .c(t_960), .d(t_2804), .cin(t_2807), .o(t_2808), .co(t_2809), .cout(t_2810));
compressor_4_2 u2_1009(.a(t_2162), .b(t_2159), .c(t_2156), .d(t_2176), .cin(t_2173), .o(t_2811), .co(t_2812), .cout(t_2813));
compressor_4_2 u2_1010(.a(t_2181), .b(t_2178), .c(t_983), .d(t_2810), .cin(t_2813), .o(t_2814), .co(t_2815), .cout(t_2816));
compressor_4_2 u2_1011(.a(t_2174), .b(t_2171), .c(t_2168), .d(t_2187), .cin(t_2184), .o(t_2817), .co(t_2818), .cout(t_2819));
compressor_4_2 u2_1012(.a(t_2192), .b(t_2189), .c(t_1006), .d(t_2816), .cin(t_2819), .o(t_2820), .co(t_2821), .cout(t_2822));
compressor_4_2 u2_1013(.a(t_2185), .b(t_2182), .c(t_2179), .d(t_2198), .cin(t_2195), .o(t_2823), .co(t_2824), .cout(t_2825));
compressor_4_2 u2_1014(.a(t_2203), .b(t_2200), .c(t_1029), .d(t_2822), .cin(t_2825), .o(t_2826), .co(t_2827), .cout(t_2828));
compressor_4_2 u2_1015(.a(t_2196), .b(t_2193), .c(t_2190), .d(t_2209), .cin(t_2206), .o(t_2829), .co(t_2830), .cout(t_2831));
compressor_4_2 u2_1016(.a(t_2214), .b(t_2211), .c(t_1052), .d(t_2828), .cin(t_2831), .o(t_2832), .co(t_2833), .cout(t_2834));
compressor_4_2 u2_1017(.a(t_2207), .b(t_2204), .c(t_2201), .d(t_2220), .cin(t_2217), .o(t_2835), .co(t_2836), .cout(t_2837));
compressor_4_2 u2_1018(.a(t_2228), .b(t_2225), .c(t_2222), .d(t_2834), .cin(t_2837), .o(t_2838), .co(t_2839), .cout(t_2840));
compressor_3_2 u1_1019(.a(t_2215), .b(t_2212), .cin(t_2231), .o(t_2841), .cout(t_2842));
compressor_4_2 u2_1020(.a(t_2236), .b(t_2233), .c(t_1096), .d(t_2840), .cin(t_2842), .o(t_2843), .co(t_2844), .cout(t_2845));
compressor_4_2 u2_1021(.a(t_2229), .b(t_2226), .c(t_2223), .d(t_2242), .cin(t_2239), .o(t_2846), .co(t_2847), .cout(t_2848));
compressor_4_2 u2_1022(.a(t_2250), .b(t_2247), .c(t_2244), .d(t_2845), .cin(t_2848), .o(t_2849), .co(t_2850), .cout(t_2851));
compressor_3_2 u1_1023(.a(t_2237), .b(t_2234), .cin(t_2253), .o(t_2852), .cout(t_2853));
compressor_4_2 u2_1024(.a(t_2261), .b(t_2258), .c(t_2255), .d(t_2851), .cin(t_2853), .o(t_2854), .co(t_2855), .cout(t_2856));
compressor_3_2 u1_1025(.a(t_2248), .b(t_2245), .cin(t_2264), .o(t_2857), .cout(t_2858));
compressor_4_2 u2_1026(.a(t_2272), .b(t_2269), .c(t_2266), .d(t_2856), .cin(t_2858), .o(t_2859), .co(t_2860), .cout(t_2861));
compressor_3_2 u1_1027(.a(t_2259), .b(t_2256), .cin(t_2275), .o(t_2862), .cout(t_2863));
compressor_4_2 u2_1028(.a(t_2283), .b(t_2280), .c(t_2277), .d(t_2861), .cin(t_2863), .o(t_2864), .co(t_2865), .cout(t_2866));
compressor_3_2 u1_1029(.a(t_2270), .b(t_2267), .cin(t_2286), .o(t_2867), .cout(t_2868));
compressor_4_2 u2_1030(.a(t_2294), .b(t_2291), .c(t_2288), .d(t_2866), .cin(t_2868), .o(t_2869), .co(t_2870), .cout(t_2871));
compressor_3_2 u1_1031(.a(t_2281), .b(t_2278), .cin(t_2297), .o(t_2872), .cout(t_2873));
compressor_4_2 u2_1032(.a(t_2305), .b(t_2302), .c(t_2299), .d(t_2871), .cin(t_2873), .o(t_2874), .co(t_2875), .cout(t_2876));
compressor_3_2 u1_1033(.a(t_2292), .b(t_2289), .cin(t_2308), .o(t_2877), .cout(t_2878));
compressor_4_2 u2_1034(.a(t_2313), .b(t_2310), .c(t_1234), .d(t_2876), .cin(t_2878), .o(t_2879), .co(t_2880), .cout(t_2881));
compressor_3_2 u1_1035(.a(t_2303), .b(t_2300), .cin(t_2316), .o(t_2882), .cout(t_2883));
compressor_4_2 u2_1036(.a(t_2322), .b(t_2319), .c(t_1252), .d(t_2881), .cin(t_2883), .o(t_2884), .co(t_2885), .cout(t_2886));
compressor_3_2 u1_1037(.a(t_2314), .b(t_2311), .cin(t_2325), .o(t_2887), .cout(t_2888));
compressor_4_2 u2_1038(.a(t_2334), .b(t_2331), .c(t_2328), .d(t_2886), .cin(t_2888), .o(t_2889), .co(t_2890), .cout(t_2891));
compressor_3_2 u1_1039(.a(t_2326), .b(t_2323), .cin(t_2320), .o(t_2892), .cout(t_2893));
compressor_4_2 u2_1040(.a(t_2340), .b(t_2337), .c(t_1284), .d(t_2891), .cin(t_2893), .o(t_2894), .co(t_2895), .cout(t_2896));
compressor_3_2 u1_1041(.a(t_2332), .b(t_2329), .cin(t_2343), .o(t_2897), .cout(t_2898));
compressor_4_2 u2_1042(.a(t_2348), .b(t_2345), .c(t_1301), .d(t_2896), .cin(t_2898), .o(t_2899), .co(t_2900), .cout(t_2901));
compressor_3_2 u1_1043(.a(t_2341), .b(t_2338), .cin(t_2351), .o(t_2902), .cout(t_2903));
compressor_4_2 u2_1044(.a(t_2356), .b(t_2353), .c(t_1318), .d(t_2901), .cin(t_2903), .o(t_2904), .co(t_2905), .cout(t_2906));
compressor_3_2 u1_1045(.a(t_2349), .b(t_2346), .cin(t_2359), .o(t_2907), .cout(t_2908));
compressor_4_2 u2_1046(.a(t_2364), .b(t_2361), .c(t_1335), .d(t_2906), .cin(t_2908), .o(t_2909), .co(t_2910), .cout(t_2911));
compressor_3_2 u1_1047(.a(t_2357), .b(t_2354), .cin(t_2367), .o(t_2912), .cout(t_2913));
compressor_4_2 u2_1048(.a(t_2372), .b(t_2369), .c(t_1352), .d(t_2911), .cin(t_2913), .o(t_2914), .co(t_2915), .cout(t_2916));
compressor_3_2 u1_1049(.a(t_2365), .b(t_2362), .cin(t_2375), .o(t_2917), .cout(t_2918));
compressor_4_2 u2_1050(.a(t_2383), .b(t_2380), .c(t_2377), .d(t_2916), .cin(t_2918), .o(t_2919), .co(t_2920), .cout(t_2921));
half_adder u0_1051(.a(t_2373), .b(t_2370), .o(t_2922), .cout(t_2923));
compressor_4_2 u2_1052(.a(t_2388), .b(t_2385), .c(t_1384), .d(t_2921), .cin(t_2923), .o(t_2924), .co(t_2925), .cout(t_2926));
compressor_3_2 u1_1053(.a(t_2381), .b(t_2378), .cin(t_2391), .o(t_2927), .cout(t_2928));
compressor_4_2 u2_1054(.a(t_2399), .b(t_2396), .c(t_2393), .d(t_2926), .cin(t_2928), .o(t_2929), .co(t_2930), .cout(t_2931));
half_adder u0_1055(.a(t_2389), .b(t_2386), .o(t_2932), .cout(t_2933));
compressor_4_2 u2_1056(.a(t_2407), .b(t_2404), .c(t_2401), .d(t_2931), .cin(t_2933), .o(t_2934), .co(t_2935), .cout(t_2936));
half_adder u0_1057(.a(t_2397), .b(t_2394), .o(t_2937), .cout(t_2938));
compressor_4_2 u2_1058(.a(t_2415), .b(t_2412), .c(t_2409), .d(t_2936), .cin(t_2938), .o(t_2939), .co(t_2940), .cout(t_2941));
half_adder u0_1059(.a(t_2405), .b(t_2402), .o(t_2942), .cout(t_2943));
compressor_4_2 u2_1060(.a(t_2423), .b(t_2420), .c(t_2417), .d(t_2941), .cin(t_2943), .o(t_2944), .co(t_2945), .cout(t_2946));
half_adder u0_1061(.a(t_2413), .b(t_2410), .o(t_2947), .cout(t_2948));
compressor_4_2 u2_1062(.a(t_2431), .b(t_2428), .c(t_2425), .d(t_2946), .cin(t_2948), .o(t_2949), .co(t_2950), .cout(t_2951));
half_adder u0_1063(.a(t_2421), .b(t_2418), .o(t_2952), .cout(t_2953));
compressor_4_2 u2_1064(.a(t_2439), .b(t_2436), .c(t_2433), .d(t_2951), .cin(t_2953), .o(t_2954), .co(t_2955), .cout(t_2956));
half_adder u0_1065(.a(t_2429), .b(t_2426), .o(t_2957), .cout(t_2958));
compressor_4_2 u2_1066(.a(t_2444), .b(t_2441), .c(t_1480), .d(t_2956), .cin(t_2958), .o(t_2959), .co(t_2960), .cout(t_2961));
half_adder u0_1067(.a(t_2437), .b(t_2434), .o(t_2962), .cout(t_2963));
compressor_4_2 u2_1068(.a(t_2450), .b(t_2447), .c(t_1492), .d(t_2961), .cin(t_2963), .o(t_2964), .co(t_2965), .cout(t_2966));
half_adder u0_1069(.a(t_2445), .b(t_2442), .o(t_2967), .cout(t_2968));
compressor_4_2 u2_1070(.a(t_2448), .b(t_2456), .c(t_2453), .d(t_2966), .cin(t_2968), .o(t_2969), .co(t_2970), .cout(t_2971));
compressor_4_2 u2_1071(.a(t_2454), .b(t_2462), .c(t_2459), .d(t_1512), .cin(t_2971), .o(t_2972), .co(t_2973), .cout(t_2974));
compressor_4_2 u2_1072(.a(t_2460), .b(t_2467), .c(t_2464), .d(t_1523), .cin(t_2974), .o(t_2975), .co(t_2976), .cout(t_2977));
compressor_4_2 u2_1073(.a(t_2465), .b(t_2472), .c(t_2469), .d(t_1534), .cin(t_2977), .o(t_2978), .co(t_2979), .cout(t_2980));
compressor_4_2 u2_1074(.a(t_2470), .b(t_2477), .c(t_2474), .d(t_1545), .cin(t_2980), .o(t_2981), .co(t_2982), .cout(t_2983));
compressor_4_2 u2_1075(.a(t_2475), .b(t_2482), .c(t_2479), .d(t_1556), .cin(t_2983), .o(t_2984), .co(t_2985), .cout(t_2986));
compressor_3_2 u1_1076(.a(t_2487), .b(t_2484), .cin(t_2986), .o(t_2987), .cout(t_2988));
compressor_3_2 u1_1077(.a(t_2492), .b(t_2489), .cin(t_1576), .o(t_2989), .cout(t_2990));
compressor_3_2 u1_1078(.a(t_2490), .b(t_2497), .cin(t_2494), .o(t_2991), .cout(t_2992));
compressor_3_2 u1_1079(.a(t_2495), .b(t_2502), .cin(t_2499), .o(t_2993), .cout(t_2994));
compressor_3_2 u1_1080(.a(t_2500), .b(t_2507), .cin(t_2504), .o(t_2995), .cout(t_2996));
compressor_3_2 u1_1081(.a(t_2505), .b(t_2512), .cin(t_2509), .o(t_2997), .cout(t_2998));
compressor_3_2 u1_1082(.a(t_2510), .b(t_2517), .cin(t_2514), .o(t_2999), .cout(t_3000));
compressor_3_2 u1_1083(.a(t_2515), .b(t_2522), .cin(t_2519), .o(t_3001), .cout(t_3002));
compressor_3_2 u1_1084(.a(t_2520), .b(t_2524), .cin(t_1630), .o(t_3003), .cout(t_3004));
compressor_3_2 u1_1085(.a(t_2525), .b(t_2527), .cin(t_1636), .o(t_3005), .cout(t_3006));
half_adder u0_1086(.a(t_2528), .b(t_2530), .o(t_3007), .cout(t_3008));
compressor_3_2 u1_1087(.a(t_2531), .b(t_2533), .cin(t_1644), .o(t_3009), .cout(t_3010));
half_adder u0_1088(.a(t_2534), .b(t_2535), .o(t_3011), .cout(t_3012));
half_adder u0_1089(.a(t_2536), .b(t_2537), .o(t_3013), .cout(t_3014));
half_adder u0_1090(.a(t_2538), .b(t_2539), .o(t_3015), .cout(t_3016));
half_adder u0_1091(.a(t_2540), .b(t_2541), .o(t_3017), .cout(t_3018));
half_adder u0_1092(.a(t_2542), .b(t_2543), .o(t_3019), .cout(t_3020));
half_adder u0_1093(.a(t_2544), .b(t_2545), .o(t_3021), .cout(t_3022));
half_adder u0_1094(.a(t_2546), .b(t_2547), .o(t_3023), .cout(t_3024));
half_adder u0_1095(.a(t_2548), .b(t_2549), .o(t_3025), .cout(t_3026));
half_adder u0_1096(.a(t_2550), .b(t_2551), .o(t_3027), .cout());

/* u0_1097 Output nets */
wire t_3028,   t_3029;
/* u0_1098 Output nets */
wire t_3030,   t_3031;
/* u0_1099 Output nets */
wire t_3032,   t_3033;
/* u0_1100 Output nets */
wire t_3034,   t_3035;
/* u0_1101 Output nets */
wire t_3036,   t_3037;
/* u0_1102 Output nets */
wire t_3038,   t_3039;
/* u0_1103 Output nets */
wire t_3040,   t_3041;
/* u0_1104 Output nets */
wire t_3042,   t_3043;
/* u0_1105 Output nets */
wire t_3044,   t_3045;
/* u0_1106 Output nets */
wire t_3046,   t_3047;
/* u0_1107 Output nets */
wire t_3048,   t_3049;
/* u0_1108 Output nets */
wire t_3050,   t_3051;
/* u0_1109 Output nets */
wire t_3052,   t_3053;
/* u0_1110 Output nets */
wire t_3054,   t_3055;
/* u0_1111 Output nets */
wire t_3056,   t_3057;
/* u1_1112 Output nets */
wire t_3058,   t_3059;
/* u0_1113 Output nets */
wire t_3060,   t_3061;
/* u0_1114 Output nets */
wire t_3062,   t_3063;
/* u1_1115 Output nets */
wire t_3064,   t_3065;
/* u0_1116 Output nets */
wire t_3066,   t_3067;
/* u0_1117 Output nets */
wire t_3068,   t_3069;
/* u0_1118 Output nets */
wire t_3070,   t_3071;
/* u0_1119 Output nets */
wire t_3072,   t_3073;
/* u0_1120 Output nets */
wire t_3074,   t_3075;
/* u1_1121 Output nets */
wire t_3076,   t_3077;
/* u1_1122 Output nets */
wire t_3078,   t_3079;
/* u1_1123 Output nets */
wire t_3080,   t_3081;
/* u1_1124 Output nets */
wire t_3082,   t_3083;
/* u1_1125 Output nets */
wire t_3084,   t_3085;
/* u1_1126 Output nets */
wire t_3086,   t_3087;
/* u1_1127 Output nets */
wire t_3088,   t_3089;
/* u1_1128 Output nets */
wire t_3090,   t_3091;
/* u1_1129 Output nets */
wire t_3092,   t_3093;
/* u1_1130 Output nets */
wire t_3094,   t_3095;
/* u1_1131 Output nets */
wire t_3096,   t_3097;
/* u2_1132 Output nets */
wire t_3098,   t_3099,   t_3100;
/* u1_1133 Output nets */
wire t_3101,   t_3102;
/* u1_1134 Output nets */
wire t_3103,   t_3104;
/* u1_1135 Output nets */
wire t_3105,   t_3106;
/* u1_1136 Output nets */
wire t_3107,   t_3108;
/* u2_1137 Output nets */
wire t_3109,   t_3110,   t_3111;
/* u2_1138 Output nets */
wire t_3112,   t_3113,   t_3114;
/* u2_1139 Output nets */
wire t_3115,   t_3116,   t_3117;
/* u2_1140 Output nets */
wire t_3118,   t_3119,   t_3120;
/* u2_1141 Output nets */
wire t_3121,   t_3122,   t_3123;
/* u1_1142 Output nets */
wire t_3124,   t_3125;
/* u2_1143 Output nets */
wire t_3126,   t_3127,   t_3128;
/* u2_1144 Output nets */
wire t_3129,   t_3130,   t_3131;
/* u1_1145 Output nets */
wire t_3132,   t_3133;
/* u1_1146 Output nets */
wire t_3134,   t_3135;
/* u2_1147 Output nets */
wire t_3136,   t_3137,   t_3138;
/* u2_1148 Output nets */
wire t_3139,   t_3140,   t_3141;
/* u2_1149 Output nets */
wire t_3142,   t_3143,   t_3144;
/* u2_1150 Output nets */
wire t_3145,   t_3146,   t_3147;
/* u2_1151 Output nets */
wire t_3148,   t_3149,   t_3150;
/* u2_1152 Output nets */
wire t_3151,   t_3152,   t_3153;
/* u2_1153 Output nets */
wire t_3154,   t_3155,   t_3156;
/* u2_1154 Output nets */
wire t_3157,   t_3158,   t_3159;
/* u2_1155 Output nets */
wire t_3160,   t_3161,   t_3162;
/* u2_1156 Output nets */
wire t_3163,   t_3164,   t_3165;
/* u2_1157 Output nets */
wire t_3166,   t_3167,   t_3168;
/* u2_1158 Output nets */
wire t_3169,   t_3170,   t_3171;
/* u2_1159 Output nets */
wire t_3172,   t_3173,   t_3174;
/* u2_1160 Output nets */
wire t_3175,   t_3176,   t_3177;
/* u2_1161 Output nets */
wire t_3178,   t_3179,   t_3180;
/* u2_1162 Output nets */
wire t_3181,   t_3182,   t_3183;
/* u2_1163 Output nets */
wire t_3184,   t_3185,   t_3186;
/* u2_1164 Output nets */
wire t_3187,   t_3188,   t_3189;
/* u1_1165 Output nets */
wire t_3190,   t_3191;
/* u2_1166 Output nets */
wire t_3192,   t_3193,   t_3194;
/* u2_1167 Output nets */
wire t_3195,   t_3196,   t_3197;
/* u2_1168 Output nets */
wire t_3198,   t_3199,   t_3200;
/* u2_1169 Output nets */
wire t_3201,   t_3202,   t_3203;
/* u2_1170 Output nets */
wire t_3204,   t_3205,   t_3206;
/* u2_1171 Output nets */
wire t_3207,   t_3208,   t_3209;
/* u2_1172 Output nets */
wire t_3210,   t_3211,   t_3212;
/* u2_1173 Output nets */
wire t_3213,   t_3214,   t_3215;
/* u1_1174 Output nets */
wire t_3216,   t_3217;
/* u1_1175 Output nets */
wire t_3218,   t_3219;
/* u1_1176 Output nets */
wire t_3220,   t_3221;
/* u1_1177 Output nets */
wire t_3222,   t_3223;
/* u1_1178 Output nets */
wire t_3224,   t_3225;
/* u1_1179 Output nets */
wire t_3226,   t_3227;
/* u1_1180 Output nets */
wire t_3228,   t_3229;
/* u1_1181 Output nets */
wire t_3230,   t_3231;
/* u1_1182 Output nets */
wire t_3232,   t_3233;
/* u1_1183 Output nets */
wire t_3234,   t_3235;
/* u1_1184 Output nets */
wire t_3236,   t_3237;
/* u1_1185 Output nets */
wire t_3238,   t_3239;
/* u1_1186 Output nets */
wire t_3240,   t_3241;
/* u1_1187 Output nets */
wire t_3242,   t_3243;
/* u1_1188 Output nets */
wire t_3244,   t_3245;
/* u1_1189 Output nets */
wire t_3246,   t_3247;
/* u1_1190 Output nets */
wire t_3248,   t_3249;
/* u1_1191 Output nets */
wire t_3250,   t_3251;
/* u0_1192 Output nets */
wire t_3252,   t_3253;
/* u0_1193 Output nets */
wire t_3254,   t_3255;
/* u0_1194 Output nets */
wire t_3256,   t_3257;
/* u0_1195 Output nets */
wire t_3258,   t_3259;
/* u1_1196 Output nets */
wire t_3260,   t_3261;
/* u1_1197 Output nets */
wire t_3262,   t_3263;
/* u0_1198 Output nets */
wire t_3264,   t_3265;
/* u0_1199 Output nets */
wire t_3266,   t_3267;
/* u0_1200 Output nets */
wire t_3268,   t_3269;
/* u0_1201 Output nets */
wire t_3270,   t_3271;
/* u0_1202 Output nets */
wire t_3272,   t_3273;
/* u0_1203 Output nets */
wire t_3274,   t_3275;
/* u0_1204 Output nets */
wire t_3276,   t_3277;
/* u0_1205 Output nets */
wire t_3278,   t_3279;
/* u0_1206 Output nets */
wire t_3280,   t_3281;
/* u0_1207 Output nets */
wire t_3282,   t_3283;
/* u0_1208 Output nets */
wire t_3284,   t_3285;
/* u0_1209 Output nets */
wire t_3286,   t_3287;
/* u0_1210 Output nets */
wire t_3288,   t_3289;
/* u0_1211 Output nets */
wire t_3290,   t_3291;
/* u0_1212 Output nets */
wire t_3292,   t_3293;
/* u0_1213 Output nets */
wire t_3294,   t_3295;
/* u0_1214 Output nets */
wire t_3296,   t_3297;
/* u0_1215 Output nets */
wire t_3298,   t_3299;
/* u0_1216 Output nets */
wire t_3300;

/* compress stage 4 */
half_adder u0_1097(.a(t_2553), .b(t_1683), .o(t_3028), .cout(t_3029));
half_adder u0_1098(.a(t_2555), .b(t_1685), .o(t_3030), .cout(t_3031));
half_adder u0_1099(.a(t_2557), .b(t_2558), .o(t_3032), .cout(t_3033));
half_adder u0_1100(.a(t_2559), .b(t_2560), .o(t_3034), .cout(t_3035));
half_adder u0_1101(.a(t_2561), .b(t_2562), .o(t_3036), .cout(t_3037));
half_adder u0_1102(.a(t_2563), .b(t_1695), .o(t_3038), .cout(t_3039));
half_adder u0_1103(.a(t_2565), .b(t_2566), .o(t_3040), .cout(t_3041));
half_adder u0_1104(.a(t_2567), .b(t_2568), .o(t_3042), .cout(t_3043));
half_adder u0_1105(.a(t_2569), .b(t_2570), .o(t_3044), .cout(t_3045));
half_adder u0_1106(.a(t_2571), .b(t_2572), .o(t_3046), .cout(t_3047));
half_adder u0_1107(.a(t_2573), .b(t_2574), .o(t_3048), .cout(t_3049));
half_adder u0_1108(.a(t_2575), .b(t_2576), .o(t_3050), .cout(t_3051));
half_adder u0_1109(.a(t_2577), .b(t_2578), .o(t_3052), .cout(t_3053));
half_adder u0_1110(.a(t_2579), .b(t_2580), .o(t_3054), .cout(t_3055));
half_adder u0_1111(.a(t_2581), .b(t_2582), .o(t_3056), .cout(t_3057));
compressor_3_2 u1_1112(.a(t_2585), .b(t_2587), .cin(t_1733), .o(t_3058), .cout(t_3059));
half_adder u0_1113(.a(t_2588), .b(t_2589), .o(t_3060), .cout(t_3061));
half_adder u0_1114(.a(t_2592), .b(t_2594), .o(t_3062), .cout(t_3063));
compressor_3_2 u1_1115(.a(t_2595), .b(t_2597), .cin(t_1753), .o(t_3064), .cout(t_3065));
half_adder u0_1116(.a(t_2598), .b(t_2599), .o(t_3066), .cout(t_3067));
half_adder u0_1117(.a(t_2600), .b(t_2602), .o(t_3068), .cout(t_3069));
half_adder u0_1118(.a(t_2603), .b(t_2605), .o(t_3070), .cout(t_3071));
half_adder u0_1119(.a(t_2606), .b(t_2608), .o(t_3072), .cout(t_3073));
half_adder u0_1120(.a(t_2609), .b(t_2611), .o(t_3074), .cout(t_3075));
compressor_3_2 u1_1121(.a(t_2612), .b(t_2614), .cin(t_1789), .o(t_3076), .cout(t_3077));
compressor_3_2 u1_1122(.a(t_2615), .b(t_2617), .cin(t_1795), .o(t_3078), .cout(t_3079));
compressor_3_2 u1_1123(.a(t_2618), .b(t_2620), .cin(t_1801), .o(t_3080), .cout(t_3081));
compressor_3_2 u1_1124(.a(t_2621), .b(t_2623), .cin(t_1807), .o(t_3082), .cout(t_3083));
compressor_3_2 u1_1125(.a(t_2624), .b(t_2626), .cin(t_1815), .o(t_3084), .cout(t_3085));
compressor_3_2 u1_1126(.a(t_2627), .b(t_2632), .cin(t_2629), .o(t_3086), .cout(t_3087));
compressor_3_2 u1_1127(.a(t_2630), .b(t_2637), .cin(t_2634), .o(t_3088), .cout(t_3089));
compressor_3_2 u1_1128(.a(t_2635), .b(t_2642), .cin(t_2639), .o(t_3090), .cout(t_3091));
compressor_3_2 u1_1129(.a(t_2640), .b(t_2647), .cin(t_2644), .o(t_3092), .cout(t_3093));
compressor_3_2 u1_1130(.a(t_2645), .b(t_2652), .cin(t_2649), .o(t_3094), .cout(t_3095));
compressor_3_2 u1_1131(.a(t_2650), .b(t_2657), .cin(t_2654), .o(t_3096), .cout(t_3097));
compressor_4_2 u2_1132(.a(t_2655), .b(t_2662), .c(t_2659), .d(t_1874), .cin(t_3097), .o(t_3098), .co(t_3099), .cout(t_3100));
compressor_3_2 u1_1133(.a(t_2667), .b(t_2664), .cin(t_3100), .o(t_3101), .cout(t_3102));
compressor_3_2 u1_1134(.a(t_2665), .b(t_2672), .cin(t_2669), .o(t_3103), .cout(t_3104));
compressor_3_2 u1_1135(.a(t_2670), .b(t_2677), .cin(t_2674), .o(t_3105), .cout(t_3106));
compressor_3_2 u1_1136(.a(t_2675), .b(t_2682), .cin(t_2679), .o(t_3107), .cout(t_3108));
compressor_4_2 u2_1137(.a(t_2680), .b(t_2687), .c(t_2684), .d(t_1917), .cin(t_3108), .o(t_3109), .co(t_3110), .cout(t_3111));
compressor_4_2 u2_1138(.a(t_2685), .b(t_2692), .c(t_2689), .d(t_1926), .cin(t_3111), .o(t_3112), .co(t_3113), .cout(t_3114));
compressor_4_2 u2_1139(.a(t_2690), .b(t_2697), .c(t_2694), .d(t_1935), .cin(t_3114), .o(t_3115), .co(t_3116), .cout(t_3117));
compressor_4_2 u2_1140(.a(t_2695), .b(t_2702), .c(t_2699), .d(t_1944), .cin(t_3117), .o(t_3118), .co(t_3119), .cout(t_3120));
compressor_4_2 u2_1141(.a(t_2700), .b(t_2707), .c(t_2704), .d(t_1955), .cin(t_3120), .o(t_3121), .co(t_3122), .cout(t_3123));
compressor_3_2 u1_1142(.a(t_2712), .b(t_2709), .cin(t_3123), .o(t_3124), .cout(t_3125));
compressor_4_2 u2_1143(.a(t_2713), .b(t_2710), .c(t_2718), .d(t_2715), .cin(t_1977), .o(t_3126), .co(t_3127), .cout(t_3128));
compressor_4_2 u2_1144(.a(t_2716), .b(t_2723), .c(t_2720), .d(t_1988), .cin(t_3128), .o(t_3129), .co(t_3130), .cout(t_3131));
compressor_3_2 u1_1145(.a(t_2728), .b(t_2725), .cin(t_3131), .o(t_3132), .cout(t_3133));
compressor_3_2 u1_1146(.a(t_2726), .b(t_2734), .cin(t_2731), .o(t_3134), .cout(t_3135));
compressor_4_2 u2_1147(.a(t_2732), .b(t_2740), .c(t_2737), .d(t_2021), .cin(t_3135), .o(t_3136), .co(t_3137), .cout(t_3138));
compressor_4_2 u2_1148(.a(t_2738), .b(t_2745), .c(t_2742), .d(t_2035), .cin(t_3138), .o(t_3139), .co(t_3140), .cout(t_3141));
compressor_4_2 u2_1149(.a(t_2746), .b(t_2743), .c(t_2751), .d(t_2748), .cin(t_3141), .o(t_3142), .co(t_3143), .cout(t_3144));
compressor_4_2 u2_1150(.a(t_2752), .b(t_2749), .c(t_2757), .d(t_2754), .cin(t_3144), .o(t_3145), .co(t_3146), .cout(t_3147));
compressor_4_2 u2_1151(.a(t_2758), .b(t_2755), .c(t_2763), .d(t_2760), .cin(t_3147), .o(t_3148), .co(t_3149), .cout(t_3150));
compressor_4_2 u2_1152(.a(t_2764), .b(t_2761), .c(t_2769), .d(t_2766), .cin(t_3150), .o(t_3151), .co(t_3152), .cout(t_3153));
compressor_4_2 u2_1153(.a(t_2767), .b(t_2775), .c(t_2772), .d(t_2093), .cin(t_3153), .o(t_3154), .co(t_3155), .cout(t_3156));
compressor_4_2 u2_1154(.a(t_2773), .b(t_2781), .c(t_2778), .d(t_2105), .cin(t_3156), .o(t_3157), .co(t_3158), .cout(t_3159));
compressor_4_2 u2_1155(.a(t_2782), .b(t_2779), .c(t_2787), .d(t_2784), .cin(t_3159), .o(t_3160), .co(t_3161), .cout(t_3162));
compressor_4_2 u2_1156(.a(t_2788), .b(t_2785), .c(t_2793), .d(t_2790), .cin(t_3162), .o(t_3163), .co(t_3164), .cout(t_3165));
compressor_4_2 u2_1157(.a(t_2791), .b(t_2799), .c(t_2796), .d(t_2141), .cin(t_3165), .o(t_3166), .co(t_3167), .cout(t_3168));
compressor_4_2 u2_1158(.a(t_2800), .b(t_2797), .c(t_2805), .d(t_2802), .cin(t_3168), .o(t_3169), .co(t_3170), .cout(t_3171));
compressor_4_2 u2_1159(.a(t_2803), .b(t_2811), .c(t_2808), .d(t_2165), .cin(t_3171), .o(t_3172), .co(t_3173), .cout(t_3174));
compressor_4_2 u2_1160(.a(t_2812), .b(t_2809), .c(t_2817), .d(t_2814), .cin(t_3174), .o(t_3175), .co(t_3176), .cout(t_3177));
compressor_4_2 u2_1161(.a(t_2818), .b(t_2815), .c(t_2823), .d(t_2820), .cin(t_3177), .o(t_3178), .co(t_3179), .cout(t_3180));
compressor_4_2 u2_1162(.a(t_2824), .b(t_2821), .c(t_2829), .d(t_2826), .cin(t_3180), .o(t_3181), .co(t_3182), .cout(t_3183));
compressor_4_2 u2_1163(.a(t_2830), .b(t_2827), .c(t_2835), .d(t_2832), .cin(t_3183), .o(t_3184), .co(t_3185), .cout(t_3186));
compressor_4_2 u2_1164(.a(t_2833), .b(t_2841), .c(t_2838), .d(t_2218), .cin(t_3186), .o(t_3187), .co(t_3188), .cout(t_3189));
compressor_3_2 u1_1165(.a(t_2846), .b(t_2843), .cin(t_3189), .o(t_3190), .cout(t_3191));
compressor_4_2 u2_1166(.a(t_2847), .b(t_2844), .c(t_2852), .d(t_2849), .cin(t_2240), .o(t_3192), .co(t_3193), .cout(t_3194));
compressor_4_2 u2_1167(.a(t_2850), .b(t_2857), .c(t_2854), .d(t_2251), .cin(t_3194), .o(t_3195), .co(t_3196), .cout(t_3197));
compressor_4_2 u2_1168(.a(t_2855), .b(t_2862), .c(t_2859), .d(t_2262), .cin(t_3197), .o(t_3198), .co(t_3199), .cout(t_3200));
compressor_4_2 u2_1169(.a(t_2860), .b(t_2867), .c(t_2864), .d(t_2273), .cin(t_3200), .o(t_3201), .co(t_3202), .cout(t_3203));
compressor_4_2 u2_1170(.a(t_2865), .b(t_2872), .c(t_2869), .d(t_2284), .cin(t_3203), .o(t_3204), .co(t_3205), .cout(t_3206));
compressor_4_2 u2_1171(.a(t_2870), .b(t_2877), .c(t_2874), .d(t_2295), .cin(t_3206), .o(t_3207), .co(t_3208), .cout(t_3209));
compressor_4_2 u2_1172(.a(t_2875), .b(t_2882), .c(t_2879), .d(t_2306), .cin(t_3209), .o(t_3210), .co(t_3211), .cout(t_3212));
compressor_4_2 u2_1173(.a(t_2880), .b(t_2887), .c(t_2884), .d(t_2317), .cin(t_3212), .o(t_3213), .co(t_3214), .cout(t_3215));
compressor_3_2 u1_1174(.a(t_2892), .b(t_2889), .cin(t_3215), .o(t_3216), .cout(t_3217));
compressor_3_2 u1_1175(.a(t_2897), .b(t_2894), .cin(t_2335), .o(t_3218), .cout(t_3219));
compressor_3_2 u1_1176(.a(t_2895), .b(t_2902), .cin(t_2899), .o(t_3220), .cout(t_3221));
compressor_3_2 u1_1177(.a(t_2900), .b(t_2907), .cin(t_2904), .o(t_3222), .cout(t_3223));
compressor_3_2 u1_1178(.a(t_2905), .b(t_2912), .cin(t_2909), .o(t_3224), .cout(t_3225));
compressor_3_2 u1_1179(.a(t_2910), .b(t_2917), .cin(t_2914), .o(t_3226), .cout(t_3227));
compressor_3_2 u1_1180(.a(t_2915), .b(t_2922), .cin(t_2919), .o(t_3228), .cout(t_3229));
compressor_3_2 u1_1181(.a(t_2920), .b(t_2927), .cin(t_2924), .o(t_3230), .cout(t_3231));
compressor_3_2 u1_1182(.a(t_2925), .b(t_2932), .cin(t_2929), .o(t_3232), .cout(t_3233));
compressor_3_2 u1_1183(.a(t_2930), .b(t_2937), .cin(t_2934), .o(t_3234), .cout(t_3235));
compressor_3_2 u1_1184(.a(t_2935), .b(t_2942), .cin(t_2939), .o(t_3236), .cout(t_3237));
compressor_3_2 u1_1185(.a(t_2940), .b(t_2947), .cin(t_2944), .o(t_3238), .cout(t_3239));
compressor_3_2 u1_1186(.a(t_2945), .b(t_2952), .cin(t_2949), .o(t_3240), .cout(t_3241));
compressor_3_2 u1_1187(.a(t_2950), .b(t_2957), .cin(t_2954), .o(t_3242), .cout(t_3243));
compressor_3_2 u1_1188(.a(t_2955), .b(t_2962), .cin(t_2959), .o(t_3244), .cout(t_3245));
compressor_3_2 u1_1189(.a(t_2960), .b(t_2967), .cin(t_2964), .o(t_3246), .cout(t_3247));
compressor_3_2 u1_1190(.a(t_2965), .b(t_2969), .cin(t_2451), .o(t_3248), .cout(t_3249));
compressor_3_2 u1_1191(.a(t_2970), .b(t_2972), .cin(t_2457), .o(t_3250), .cout(t_3251));
half_adder u0_1192(.a(t_2973), .b(t_2975), .o(t_3252), .cout(t_3253));
half_adder u0_1193(.a(t_2976), .b(t_2978), .o(t_3254), .cout(t_3255));
half_adder u0_1194(.a(t_2979), .b(t_2981), .o(t_3256), .cout(t_3257));
half_adder u0_1195(.a(t_2982), .b(t_2984), .o(t_3258), .cout(t_3259));
compressor_3_2 u1_1196(.a(t_2985), .b(t_2987), .cin(t_2480), .o(t_3260), .cout(t_3261));
compressor_3_2 u1_1197(.a(t_2988), .b(t_2989), .cin(t_2485), .o(t_3262), .cout(t_3263));
half_adder u0_1198(.a(t_2990), .b(t_2991), .o(t_3264), .cout(t_3265));
half_adder u0_1199(.a(t_2992), .b(t_2993), .o(t_3266), .cout(t_3267));
half_adder u0_1200(.a(t_2994), .b(t_2995), .o(t_3268), .cout(t_3269));
half_adder u0_1201(.a(t_2996), .b(t_2997), .o(t_3270), .cout(t_3271));
half_adder u0_1202(.a(t_2998), .b(t_2999), .o(t_3272), .cout(t_3273));
half_adder u0_1203(.a(t_3000), .b(t_3001), .o(t_3274), .cout(t_3275));
half_adder u0_1204(.a(t_3002), .b(t_3003), .o(t_3276), .cout(t_3277));
half_adder u0_1205(.a(t_3004), .b(t_3005), .o(t_3278), .cout(t_3279));
half_adder u0_1206(.a(t_3006), .b(t_3007), .o(t_3280), .cout(t_3281));
half_adder u0_1207(.a(t_3008), .b(t_3009), .o(t_3282), .cout(t_3283));
half_adder u0_1208(.a(t_3010), .b(t_3011), .o(t_3284), .cout(t_3285));
half_adder u0_1209(.a(t_3012), .b(t_3013), .o(t_3286), .cout(t_3287));
half_adder u0_1210(.a(t_3014), .b(t_3015), .o(t_3288), .cout(t_3289));
half_adder u0_1211(.a(t_3016), .b(t_3017), .o(t_3290), .cout(t_3291));
half_adder u0_1212(.a(t_3018), .b(t_3019), .o(t_3292), .cout(t_3293));
half_adder u0_1213(.a(t_3020), .b(t_3021), .o(t_3294), .cout(t_3295));
half_adder u0_1214(.a(t_3022), .b(t_3023), .o(t_3296), .cout(t_3297));
half_adder u0_1215(.a(t_3024), .b(t_3025), .o(t_3298), .cout(t_3299));
half_adder u0_1216(.a(t_3026), .b(t_3027), .o(t_3300), .cout());

/* u0_1217 Output nets */
wire t_3301,   t_3302;
/* u0_1218 Output nets */
wire t_3303,   t_3304;
/* u0_1219 Output nets */
wire t_3305,   t_3306;
/* u0_1220 Output nets */
wire t_3307,   t_3308;
/* u0_1221 Output nets */
wire t_3309,   t_3310;
/* u0_1222 Output nets */
wire t_3311,   t_3312;
/* u0_1223 Output nets */
wire t_3313,   t_3314;
/* u0_1224 Output nets */
wire t_3315,   t_3316;
/* u0_1225 Output nets */
wire t_3317,   t_3318;
/* u0_1226 Output nets */
wire t_3319,   t_3320;
/* u0_1227 Output nets */
wire t_3321,   t_3322;
/* u0_1228 Output nets */
wire t_3323,   t_3324;
/* u0_1229 Output nets */
wire t_3325,   t_3326;
/* u0_1230 Output nets */
wire t_3327,   t_3328;
/* u0_1231 Output nets */
wire t_3329,   t_3330;
/* u0_1232 Output nets */
wire t_3331,   t_3332;
/* u0_1233 Output nets */
wire t_3333,   t_3334;
/* u0_1234 Output nets */
wire t_3335,   t_3336;
/* u0_1235 Output nets */
wire t_3337,   t_3338;
/* u0_1236 Output nets */
wire t_3339,   t_3340;
/* u0_1237 Output nets */
wire t_3341,   t_3342;
/* u0_1238 Output nets */
wire t_3343,   t_3344;
/* u0_1239 Output nets */
wire t_3345,   t_3346;
/* u0_1240 Output nets */
wire t_3347,   t_3348;
/* u0_1241 Output nets */
wire t_3349,   t_3350;
/* u0_1242 Output nets */
wire t_3351,   t_3352;
/* u0_1243 Output nets */
wire t_3353,   t_3354;
/* u0_1244 Output nets */
wire t_3355,   t_3356;
/* u0_1245 Output nets */
wire t_3357,   t_3358;
/* u0_1246 Output nets */
wire t_3359,   t_3360;
/* u0_1247 Output nets */
wire t_3361,   t_3362;
/* u0_1248 Output nets */
wire t_3363,   t_3364;
/* u0_1249 Output nets */
wire t_3365,   t_3366;
/* u0_1250 Output nets */
wire t_3367,   t_3368;
/* u1_1251 Output nets */
wire t_3369,   t_3370;
/* u0_1252 Output nets */
wire t_3371,   t_3372;
/* u0_1253 Output nets */
wire t_3373,   t_3374;
/* u0_1254 Output nets */
wire t_3375,   t_3376;
/* u0_1255 Output nets */
wire t_3377,   t_3378;
/* u0_1256 Output nets */
wire t_3379,   t_3380;
/* u0_1257 Output nets */
wire t_3381,   t_3382;
/* u0_1258 Output nets */
wire t_3383,   t_3384;
/* u1_1259 Output nets */
wire t_3385,   t_3386;
/* u0_1260 Output nets */
wire t_3387,   t_3388;
/* u0_1261 Output nets */
wire t_3389,   t_3390;
/* u1_1262 Output nets */
wire t_3391,   t_3392;
/* u1_1263 Output nets */
wire t_3393,   t_3394;
/* u0_1264 Output nets */
wire t_3395,   t_3396;
/* u0_1265 Output nets */
wire t_3397,   t_3398;
/* u0_1266 Output nets */
wire t_3399,   t_3400;
/* u0_1267 Output nets */
wire t_3401,   t_3402;
/* u0_1268 Output nets */
wire t_3403,   t_3404;
/* u0_1269 Output nets */
wire t_3405,   t_3406;
/* u1_1270 Output nets */
wire t_3407,   t_3408;
/* u1_1271 Output nets */
wire t_3409,   t_3410;
/* u0_1272 Output nets */
wire t_3411,   t_3412;
/* u0_1273 Output nets */
wire t_3413,   t_3414;
/* u1_1274 Output nets */
wire t_3415,   t_3416;
/* u0_1275 Output nets */
wire t_3417,   t_3418;
/* u1_1276 Output nets */
wire t_3419,   t_3420;
/* u0_1277 Output nets */
wire t_3421,   t_3422;
/* u0_1278 Output nets */
wire t_3423,   t_3424;
/* u0_1279 Output nets */
wire t_3425,   t_3426;
/* u0_1280 Output nets */
wire t_3427,   t_3428;
/* u1_1281 Output nets */
wire t_3429,   t_3430;
/* u1_1282 Output nets */
wire t_3431,   t_3432;
/* u0_1283 Output nets */
wire t_3433,   t_3434;
/* u0_1284 Output nets */
wire t_3435,   t_3436;
/* u0_1285 Output nets */
wire t_3437,   t_3438;
/* u0_1286 Output nets */
wire t_3439,   t_3440;
/* u0_1287 Output nets */
wire t_3441,   t_3442;
/* u0_1288 Output nets */
wire t_3443,   t_3444;
/* u0_1289 Output nets */
wire t_3445,   t_3446;
/* u0_1290 Output nets */
wire t_3447,   t_3448;
/* u1_1291 Output nets */
wire t_3449,   t_3450;
/* u1_1292 Output nets */
wire t_3451,   t_3452;
/* u0_1293 Output nets */
wire t_3453,   t_3454;
/* u0_1294 Output nets */
wire t_3455,   t_3456;
/* u0_1295 Output nets */
wire t_3457,   t_3458;
/* u0_1296 Output nets */
wire t_3459,   t_3460;
/* u0_1297 Output nets */
wire t_3461,   t_3462;
/* u0_1298 Output nets */
wire t_3463,   t_3464;
/* u0_1299 Output nets */
wire t_3465,   t_3466;
/* u0_1300 Output nets */
wire t_3467,   t_3468;
/* u0_1301 Output nets */
wire t_3469,   t_3470;
/* u0_1302 Output nets */
wire t_3471,   t_3472;
/* u0_1303 Output nets */
wire t_3473,   t_3474;
/* u0_1304 Output nets */
wire t_3475,   t_3476;
/* u0_1305 Output nets */
wire t_3477,   t_3478;
/* u0_1306 Output nets */
wire t_3479,   t_3480;
/* u0_1307 Output nets */
wire t_3481,   t_3482;
/* u0_1308 Output nets */
wire t_3483,   t_3484;
/* u0_1309 Output nets */
wire t_3485,   t_3486;
/* u0_1310 Output nets */
wire t_3487,   t_3488;
/* u0_1311 Output nets */
wire t_3489,   t_3490;
/* u0_1312 Output nets */
wire t_3491,   t_3492;
/* u0_1313 Output nets */
wire t_3493,   t_3494;
/* u0_1314 Output nets */
wire t_3495,   t_3496;
/* u0_1315 Output nets */
wire t_3497,   t_3498;
/* u0_1316 Output nets */
wire t_3499,   t_3500;
/* u0_1317 Output nets */
wire t_3501,   t_3502;
/* u0_1318 Output nets */
wire t_3503,   t_3504;
/* u0_1319 Output nets */
wire t_3505,   t_3506;
/* u0_1320 Output nets */
wire t_3507,   t_3508;
/* u0_1321 Output nets */
wire t_3509,   t_3510;
/* u0_1322 Output nets */
wire t_3511,   t_3512;
/* u0_1323 Output nets */
wire t_3513,   t_3514;
/* u0_1324 Output nets */
wire t_3515,   t_3516;
/* u0_1325 Output nets */
wire t_3517,   t_3518;
/* u0_1326 Output nets */
wire t_3519,   t_3520;
/* u0_1327 Output nets */
wire t_3521,   t_3522;
/* u0_1328 Output nets */
wire t_3523,   t_3524;
/* u0_1329 Output nets */
wire t_3525,   t_3526;
/* u0_1330 Output nets */
wire t_3527,   t_3528;
/* u0_1331 Output nets */
wire t_3529,   t_3530;
/* u0_1332 Output nets */
wire t_3531,   t_3532;
/* u0_1333 Output nets */
wire t_3533;

/* compress stage 5 */
half_adder u0_1217(.a(t_3029), .b(t_2554), .o(t_3301), .cout(t_3302));
half_adder u0_1218(.a(t_3031), .b(t_2556), .o(t_3303), .cout(t_3304));
half_adder u0_1219(.a(t_3033), .b(t_3034), .o(t_3305), .cout(t_3306));
half_adder u0_1220(.a(t_3035), .b(t_3036), .o(t_3307), .cout(t_3308));
half_adder u0_1221(.a(t_3037), .b(t_3038), .o(t_3309), .cout(t_3310));
half_adder u0_1222(.a(t_3039), .b(t_2564), .o(t_3311), .cout(t_3312));
half_adder u0_1223(.a(t_3041), .b(t_3042), .o(t_3313), .cout(t_3314));
half_adder u0_1224(.a(t_3043), .b(t_3044), .o(t_3315), .cout(t_3316));
half_adder u0_1225(.a(t_3045), .b(t_3046), .o(t_3317), .cout(t_3318));
half_adder u0_1226(.a(t_3047), .b(t_3048), .o(t_3319), .cout(t_3320));
half_adder u0_1227(.a(t_3049), .b(t_3050), .o(t_3321), .cout(t_3322));
half_adder u0_1228(.a(t_3051), .b(t_3052), .o(t_3323), .cout(t_3324));
half_adder u0_1229(.a(t_3053), .b(t_3054), .o(t_3325), .cout(t_3326));
half_adder u0_1230(.a(t_3055), .b(t_3056), .o(t_3327), .cout(t_3328));
half_adder u0_1231(.a(t_3057), .b(t_2584), .o(t_3329), .cout(t_3330));
half_adder u0_1232(.a(t_3059), .b(t_3060), .o(t_3331), .cout(t_3332));
half_adder u0_1233(.a(t_3061), .b(t_2591), .o(t_3333), .cout(t_3334));
half_adder u0_1234(.a(t_3063), .b(t_3064), .o(t_3335), .cout(t_3336));
half_adder u0_1235(.a(t_3065), .b(t_3066), .o(t_3337), .cout(t_3338));
half_adder u0_1236(.a(t_3067), .b(t_3068), .o(t_3339), .cout(t_3340));
half_adder u0_1237(.a(t_3069), .b(t_3070), .o(t_3341), .cout(t_3342));
half_adder u0_1238(.a(t_3071), .b(t_3072), .o(t_3343), .cout(t_3344));
half_adder u0_1239(.a(t_3073), .b(t_3074), .o(t_3345), .cout(t_3346));
half_adder u0_1240(.a(t_3075), .b(t_3076), .o(t_3347), .cout(t_3348));
half_adder u0_1241(.a(t_3077), .b(t_3078), .o(t_3349), .cout(t_3350));
half_adder u0_1242(.a(t_3079), .b(t_3080), .o(t_3351), .cout(t_3352));
half_adder u0_1243(.a(t_3081), .b(t_3082), .o(t_3353), .cout(t_3354));
half_adder u0_1244(.a(t_3083), .b(t_3084), .o(t_3355), .cout(t_3356));
half_adder u0_1245(.a(t_3085), .b(t_3086), .o(t_3357), .cout(t_3358));
half_adder u0_1246(.a(t_3087), .b(t_3088), .o(t_3359), .cout(t_3360));
half_adder u0_1247(.a(t_3089), .b(t_3090), .o(t_3361), .cout(t_3362));
half_adder u0_1248(.a(t_3091), .b(t_3092), .o(t_3363), .cout(t_3364));
half_adder u0_1249(.a(t_3093), .b(t_3094), .o(t_3365), .cout(t_3366));
half_adder u0_1250(.a(t_3095), .b(t_3096), .o(t_3367), .cout(t_3368));
compressor_3_2 u1_1251(.a(t_3099), .b(t_3101), .cin(t_2660), .o(t_3369), .cout(t_3370));
half_adder u0_1252(.a(t_3102), .b(t_3103), .o(t_3371), .cout(t_3372));
half_adder u0_1253(.a(t_3104), .b(t_3105), .o(t_3373), .cout(t_3374));
half_adder u0_1254(.a(t_3106), .b(t_3107), .o(t_3375), .cout(t_3376));
half_adder u0_1255(.a(t_3110), .b(t_3112), .o(t_3377), .cout(t_3378));
half_adder u0_1256(.a(t_3113), .b(t_3115), .o(t_3379), .cout(t_3380));
half_adder u0_1257(.a(t_3116), .b(t_3118), .o(t_3381), .cout(t_3382));
half_adder u0_1258(.a(t_3119), .b(t_3121), .o(t_3383), .cout(t_3384));
compressor_3_2 u1_1259(.a(t_3122), .b(t_3124), .cin(t_2705), .o(t_3385), .cout(t_3386));
half_adder u0_1260(.a(t_3125), .b(t_3126), .o(t_3387), .cout(t_3388));
half_adder u0_1261(.a(t_3127), .b(t_3129), .o(t_3389), .cout(t_3390));
compressor_3_2 u1_1262(.a(t_3130), .b(t_3132), .cin(t_2721), .o(t_3391), .cout(t_3392));
compressor_3_2 u1_1263(.a(t_3133), .b(t_3134), .cin(t_2729), .o(t_3393), .cout(t_3394));
half_adder u0_1264(.a(t_3136), .b(t_2735), .o(t_3395), .cout(t_3396));
half_adder u0_1265(.a(t_3137), .b(t_3139), .o(t_3397), .cout(t_3398));
half_adder u0_1266(.a(t_3140), .b(t_3142), .o(t_3399), .cout(t_3400));
half_adder u0_1267(.a(t_3143), .b(t_3145), .o(t_3401), .cout(t_3402));
half_adder u0_1268(.a(t_3146), .b(t_3148), .o(t_3403), .cout(t_3404));
half_adder u0_1269(.a(t_3149), .b(t_3151), .o(t_3405), .cout(t_3406));
compressor_3_2 u1_1270(.a(t_3152), .b(t_3154), .cin(t_2770), .o(t_3407), .cout(t_3408));
compressor_3_2 u1_1271(.a(t_3155), .b(t_3157), .cin(t_2776), .o(t_3409), .cout(t_3410));
half_adder u0_1272(.a(t_3158), .b(t_3160), .o(t_3411), .cout(t_3412));
half_adder u0_1273(.a(t_3161), .b(t_3163), .o(t_3413), .cout(t_3414));
compressor_3_2 u1_1274(.a(t_3164), .b(t_3166), .cin(t_2794), .o(t_3415), .cout(t_3416));
half_adder u0_1275(.a(t_3167), .b(t_3169), .o(t_3417), .cout(t_3418));
compressor_3_2 u1_1276(.a(t_3170), .b(t_3172), .cin(t_2806), .o(t_3419), .cout(t_3420));
half_adder u0_1277(.a(t_3173), .b(t_3175), .o(t_3421), .cout(t_3422));
half_adder u0_1278(.a(t_3176), .b(t_3178), .o(t_3423), .cout(t_3424));
half_adder u0_1279(.a(t_3179), .b(t_3181), .o(t_3425), .cout(t_3426));
half_adder u0_1280(.a(t_3182), .b(t_3184), .o(t_3427), .cout(t_3428));
compressor_3_2 u1_1281(.a(t_3185), .b(t_3187), .cin(t_2836), .o(t_3429), .cout(t_3430));
compressor_3_2 u1_1282(.a(t_3188), .b(t_3190), .cin(t_2839), .o(t_3431), .cout(t_3432));
half_adder u0_1283(.a(t_3191), .b(t_3192), .o(t_3433), .cout(t_3434));
half_adder u0_1284(.a(t_3193), .b(t_3195), .o(t_3435), .cout(t_3436));
half_adder u0_1285(.a(t_3196), .b(t_3198), .o(t_3437), .cout(t_3438));
half_adder u0_1286(.a(t_3199), .b(t_3201), .o(t_3439), .cout(t_3440));
half_adder u0_1287(.a(t_3202), .b(t_3204), .o(t_3441), .cout(t_3442));
half_adder u0_1288(.a(t_3205), .b(t_3207), .o(t_3443), .cout(t_3444));
half_adder u0_1289(.a(t_3208), .b(t_3210), .o(t_3445), .cout(t_3446));
half_adder u0_1290(.a(t_3211), .b(t_3213), .o(t_3447), .cout(t_3448));
compressor_3_2 u1_1291(.a(t_3214), .b(t_3216), .cin(t_2885), .o(t_3449), .cout(t_3450));
compressor_3_2 u1_1292(.a(t_3217), .b(t_3218), .cin(t_2890), .o(t_3451), .cout(t_3452));
half_adder u0_1293(.a(t_3219), .b(t_3220), .o(t_3453), .cout(t_3454));
half_adder u0_1294(.a(t_3221), .b(t_3222), .o(t_3455), .cout(t_3456));
half_adder u0_1295(.a(t_3223), .b(t_3224), .o(t_3457), .cout(t_3458));
half_adder u0_1296(.a(t_3225), .b(t_3226), .o(t_3459), .cout(t_3460));
half_adder u0_1297(.a(t_3227), .b(t_3228), .o(t_3461), .cout(t_3462));
half_adder u0_1298(.a(t_3229), .b(t_3230), .o(t_3463), .cout(t_3464));
half_adder u0_1299(.a(t_3231), .b(t_3232), .o(t_3465), .cout(t_3466));
half_adder u0_1300(.a(t_3233), .b(t_3234), .o(t_3467), .cout(t_3468));
half_adder u0_1301(.a(t_3235), .b(t_3236), .o(t_3469), .cout(t_3470));
half_adder u0_1302(.a(t_3237), .b(t_3238), .o(t_3471), .cout(t_3472));
half_adder u0_1303(.a(t_3239), .b(t_3240), .o(t_3473), .cout(t_3474));
half_adder u0_1304(.a(t_3241), .b(t_3242), .o(t_3475), .cout(t_3476));
half_adder u0_1305(.a(t_3243), .b(t_3244), .o(t_3477), .cout(t_3478));
half_adder u0_1306(.a(t_3245), .b(t_3246), .o(t_3479), .cout(t_3480));
half_adder u0_1307(.a(t_3247), .b(t_3248), .o(t_3481), .cout(t_3482));
half_adder u0_1308(.a(t_3249), .b(t_3250), .o(t_3483), .cout(t_3484));
half_adder u0_1309(.a(t_3251), .b(t_3252), .o(t_3485), .cout(t_3486));
half_adder u0_1310(.a(t_3253), .b(t_3254), .o(t_3487), .cout(t_3488));
half_adder u0_1311(.a(t_3255), .b(t_3256), .o(t_3489), .cout(t_3490));
half_adder u0_1312(.a(t_3257), .b(t_3258), .o(t_3491), .cout(t_3492));
half_adder u0_1313(.a(t_3259), .b(t_3260), .o(t_3493), .cout(t_3494));
half_adder u0_1314(.a(t_3261), .b(t_3262), .o(t_3495), .cout(t_3496));
half_adder u0_1315(.a(t_3263), .b(t_3264), .o(t_3497), .cout(t_3498));
half_adder u0_1316(.a(t_3265), .b(t_3266), .o(t_3499), .cout(t_3500));
half_adder u0_1317(.a(t_3267), .b(t_3268), .o(t_3501), .cout(t_3502));
half_adder u0_1318(.a(t_3269), .b(t_3270), .o(t_3503), .cout(t_3504));
half_adder u0_1319(.a(t_3271), .b(t_3272), .o(t_3505), .cout(t_3506));
half_adder u0_1320(.a(t_3273), .b(t_3274), .o(t_3507), .cout(t_3508));
half_adder u0_1321(.a(t_3275), .b(t_3276), .o(t_3509), .cout(t_3510));
half_adder u0_1322(.a(t_3277), .b(t_3278), .o(t_3511), .cout(t_3512));
half_adder u0_1323(.a(t_3279), .b(t_3280), .o(t_3513), .cout(t_3514));
half_adder u0_1324(.a(t_3281), .b(t_3282), .o(t_3515), .cout(t_3516));
half_adder u0_1325(.a(t_3283), .b(t_3284), .o(t_3517), .cout(t_3518));
half_adder u0_1326(.a(t_3285), .b(t_3286), .o(t_3519), .cout(t_3520));
half_adder u0_1327(.a(t_3287), .b(t_3288), .o(t_3521), .cout(t_3522));
half_adder u0_1328(.a(t_3289), .b(t_3290), .o(t_3523), .cout(t_3524));
half_adder u0_1329(.a(t_3291), .b(t_3292), .o(t_3525), .cout(t_3526));
half_adder u0_1330(.a(t_3293), .b(t_3294), .o(t_3527), .cout(t_3528));
half_adder u0_1331(.a(t_3295), .b(t_3296), .o(t_3529), .cout(t_3530));
half_adder u0_1332(.a(t_3297), .b(t_3298), .o(t_3531), .cout(t_3532));
half_adder u0_1333(.a(t_3299), .b(t_3300), .o(t_3533), .cout());

/* Output nets Compression result */
assign compress_a = {
  t_3533,  t_3531,  t_3529,  t_3527,
  t_3525,  t_3523,  t_3521,  t_3519,
  t_3517,  t_3515,  t_3513,  t_3511,
  t_3509,  t_3507,  t_3505,  t_3503,
  t_3501,  t_3499,  t_3497,  t_3495,
  t_3493,  t_3491,  t_3489,  t_3487,
  t_3485,  t_3483,  t_3481,  t_3479,
  t_3477,  t_3475,  t_3473,  t_3471,
  t_3469,  t_3467,  t_3465,  t_3463,
  t_3461,  t_3459,  t_3457,  t_3455,
  t_3453,  t_3451,  t_3449,  t_3447,
  t_3445,  t_3443,  t_3441,  t_3439,
  t_3437,  t_3435,  t_3433,  t_3431,
  t_3429,  t_3427,  t_3425,  t_3423,
  t_3421,  t_3419,  t_3417,  t_3415,
  t_3413,  t_3411,  t_3409,  t_3407,
  t_3405,  t_3403,  t_3401,  t_3399,
  t_3397,  t_3395,  t_3393,  t_3391,
  t_3389,  t_3387,  t_3385,  t_3383,
  t_3381,  t_3379,  t_3377,  t_3109,
  t_3375,  t_3373,  t_3371,  t_3369,
  t_3098,  t_3367,  t_3365,  t_3363,
  t_3361,  t_3359,  t_3357,  t_3355,
  t_3353,  t_3351,  t_3349,  t_3347,
  t_3345,  t_3343,  t_3341,  t_3339,
  t_3337,  t_3335,  t_3062,  t_3333,
  t_3331,  t_3058,  t_3329,  t_3327,
  t_3325,  t_3323,  t_3321,  t_3319,
  t_3317,  t_3315,  t_3313,  t_3040,
  t_3311,  t_3309,  t_3307,  t_3305,
  t_3032,  t_3303,  t_3030,  t_3301,
  t_3028,  t_2552,  t_1681,     t_0
};
assign compress_b = {
  t_3532,  t_3530,  t_3528,  t_3526,
  t_3524,  t_3522,  t_3520,  t_3518,
  t_3516,  t_3514,  t_3512,  t_3510,
  t_3508,  t_3506,  t_3504,  t_3502,
  t_3500,  t_3498,  t_3496,  t_3494,
  t_3492,  t_3490,  t_3488,  t_3486,
  t_3484,  t_3482,  t_3480,  t_3478,
  t_3476,  t_3474,  t_3472,  t_3470,
  t_3468,  t_3466,  t_3464,  t_3462,
  t_3460,  t_3458,  t_3456,  t_3454,
  t_3452,  t_3450,  t_3448,  t_3446,
  t_3444,  t_3442,  t_3440,  t_3438,
  t_3436,  t_3434,  t_3432,  t_3430,
  t_3428,  t_3426,  t_3424,  t_3422,
  t_3420,  t_3418,  t_3416,  t_3414,
  t_3412,  t_3410,  t_3408,  t_3406,
  t_3404,  t_3402,  t_3400,  t_3398,
  t_3396,  t_3394,  t_3392,  t_3390,
  t_3388,  t_3386,  t_3384,  t_3382,
  t_3380,  t_3378,    1'b0,  t_3376,
  t_3374,  t_3372,  t_3370,    1'b0,
  t_3368,  t_3366,  t_3364,  t_3362,
  t_3360,  t_3358,  t_3356,  t_3354,
  t_3352,  t_3350,  t_3348,  t_3346,
  t_3344,  t_3342,  t_3340,  t_3338,
  t_3336,    1'b0,  t_3334,  t_3332,
    1'b0,  t_3330,  t_3328,  t_3326,
  t_3324,  t_3322,  t_3320,  t_3318,
  t_3316,  t_3314,    1'b0,  t_3312,
  t_3310,  t_3308,  t_3306,    1'b0,
  t_3304,    1'b0,  t_3302,    1'b0,
    1'b0,    1'b0,    1'b0,    1'b0
};

endmodule

/********************************************************************************/

module _128_wallace_tree(
//inputs
	partial_products,
	carry,
//outputs
	compress_a,
	compress_b
);

localparam width = 128;

input wire [(width+2)*(width/2+1)-1:0] partial_products;
input wire [width/2-1:0] carry;
output wire [2*width-1:0] compress_a;
output wire [2*width-1:0] compress_b;

/* Input nets */
wire    s_0_0,    s_0_1,    s_1_0,    s_2_0,    s_2_1,    s_2_2;
wire    s_3_0,    s_3_1,    s_4_0,    s_4_1,    s_4_2,    s_4_3;
wire    s_5_0,    s_5_1,    s_5_2,    s_6_0,    s_6_1,    s_6_2;
wire    s_6_3,    s_6_4,    s_7_0,    s_7_1,    s_7_2,    s_7_3;
wire    s_8_0,    s_8_1,    s_8_2,    s_8_3,    s_8_4,    s_8_5;
wire    s_9_0,    s_9_1,    s_9_2,    s_9_3,    s_9_4,   s_10_0;
wire   s_10_1,   s_10_2,   s_10_3,   s_10_4,   s_10_5,   s_10_6;
wire   s_11_0,   s_11_1,   s_11_2,   s_11_3,   s_11_4,   s_11_5;
wire   s_12_0,   s_12_1,   s_12_2,   s_12_3,   s_12_4,   s_12_5;
wire   s_12_6,   s_12_7,   s_13_0,   s_13_1,   s_13_2,   s_13_3;
wire   s_13_4,   s_13_5,   s_13_6,   s_14_0,   s_14_1,   s_14_2;
wire   s_14_3,   s_14_4,   s_14_5,   s_14_6,   s_14_7,   s_14_8;
wire   s_15_0,   s_15_1,   s_15_2,   s_15_3,   s_15_4,   s_15_5;
wire   s_15_6,   s_15_7,   s_16_0,   s_16_1,   s_16_2,   s_16_3;
wire   s_16_4,   s_16_5,   s_16_6,   s_16_7,   s_16_8,   s_16_9;
wire   s_17_0,   s_17_1,   s_17_2,   s_17_3,   s_17_4,   s_17_5;
wire   s_17_6,   s_17_7,   s_17_8,   s_18_0,   s_18_1,   s_18_2;
wire   s_18_3,   s_18_4,   s_18_5,   s_18_6,   s_18_7,   s_18_8;
wire   s_18_9,  s_18_10,   s_19_0,   s_19_1,   s_19_2,   s_19_3;
wire   s_19_4,   s_19_5,   s_19_6,   s_19_7,   s_19_8,   s_19_9;
wire   s_20_0,   s_20_1,   s_20_2,   s_20_3,   s_20_4,   s_20_5;
wire   s_20_6,   s_20_7,   s_20_8,   s_20_9,  s_20_10,  s_20_11;
wire   s_21_0,   s_21_1,   s_21_2,   s_21_3,   s_21_4,   s_21_5;
wire   s_21_6,   s_21_7,   s_21_8,   s_21_9,  s_21_10,   s_22_0;
wire   s_22_1,   s_22_2,   s_22_3,   s_22_4,   s_22_5,   s_22_6;
wire   s_22_7,   s_22_8,   s_22_9,  s_22_10,  s_22_11,  s_22_12;
wire   s_23_0,   s_23_1,   s_23_2,   s_23_3,   s_23_4,   s_23_5;
wire   s_23_6,   s_23_7,   s_23_8,   s_23_9,  s_23_10,  s_23_11;
wire   s_24_0,   s_24_1,   s_24_2,   s_24_3,   s_24_4,   s_24_5;
wire   s_24_6,   s_24_7,   s_24_8,   s_24_9,  s_24_10,  s_24_11;
wire  s_24_12,  s_24_13,   s_25_0,   s_25_1,   s_25_2,   s_25_3;
wire   s_25_4,   s_25_5,   s_25_6,   s_25_7,   s_25_8,   s_25_9;
wire  s_25_10,  s_25_11,  s_25_12,   s_26_0,   s_26_1,   s_26_2;
wire   s_26_3,   s_26_4,   s_26_5,   s_26_6,   s_26_7,   s_26_8;
wire   s_26_9,  s_26_10,  s_26_11,  s_26_12,  s_26_13,  s_26_14;
wire   s_27_0,   s_27_1,   s_27_2,   s_27_3,   s_27_4,   s_27_5;
wire   s_27_6,   s_27_7,   s_27_8,   s_27_9,  s_27_10,  s_27_11;
wire  s_27_12,  s_27_13,   s_28_0,   s_28_1,   s_28_2,   s_28_3;
wire   s_28_4,   s_28_5,   s_28_6,   s_28_7,   s_28_8,   s_28_9;
wire  s_28_10,  s_28_11,  s_28_12,  s_28_13,  s_28_14,  s_28_15;
wire   s_29_0,   s_29_1,   s_29_2,   s_29_3,   s_29_4,   s_29_5;
wire   s_29_6,   s_29_7,   s_29_8,   s_29_9,  s_29_10,  s_29_11;
wire  s_29_12,  s_29_13,  s_29_14,   s_30_0,   s_30_1,   s_30_2;
wire   s_30_3,   s_30_4,   s_30_5,   s_30_6,   s_30_7,   s_30_8;
wire   s_30_9,  s_30_10,  s_30_11,  s_30_12,  s_30_13,  s_30_14;
wire  s_30_15,  s_30_16,   s_31_0,   s_31_1,   s_31_2,   s_31_3;
wire   s_31_4,   s_31_5,   s_31_6,   s_31_7,   s_31_8,   s_31_9;
wire  s_31_10,  s_31_11,  s_31_12,  s_31_13,  s_31_14,  s_31_15;
wire   s_32_0,   s_32_1,   s_32_2,   s_32_3,   s_32_4,   s_32_5;
wire   s_32_6,   s_32_7,   s_32_8,   s_32_9,  s_32_10,  s_32_11;
wire  s_32_12,  s_32_13,  s_32_14,  s_32_15,  s_32_16,  s_32_17;
wire   s_33_0,   s_33_1,   s_33_2,   s_33_3,   s_33_4,   s_33_5;
wire   s_33_6,   s_33_7,   s_33_8,   s_33_9,  s_33_10,  s_33_11;
wire  s_33_12,  s_33_13,  s_33_14,  s_33_15,  s_33_16,   s_34_0;
wire   s_34_1,   s_34_2,   s_34_3,   s_34_4,   s_34_5,   s_34_6;
wire   s_34_7,   s_34_8,   s_34_9,  s_34_10,  s_34_11,  s_34_12;
wire  s_34_13,  s_34_14,  s_34_15,  s_34_16,  s_34_17,  s_34_18;
wire   s_35_0,   s_35_1,   s_35_2,   s_35_3,   s_35_4,   s_35_5;
wire   s_35_6,   s_35_7,   s_35_8,   s_35_9,  s_35_10,  s_35_11;
wire  s_35_12,  s_35_13,  s_35_14,  s_35_15,  s_35_16,  s_35_17;
wire   s_36_0,   s_36_1,   s_36_2,   s_36_3,   s_36_4,   s_36_5;
wire   s_36_6,   s_36_7,   s_36_8,   s_36_9,  s_36_10,  s_36_11;
wire  s_36_12,  s_36_13,  s_36_14,  s_36_15,  s_36_16,  s_36_17;
wire  s_36_18,  s_36_19,   s_37_0,   s_37_1,   s_37_2,   s_37_3;
wire   s_37_4,   s_37_5,   s_37_6,   s_37_7,   s_37_8,   s_37_9;
wire  s_37_10,  s_37_11,  s_37_12,  s_37_13,  s_37_14,  s_37_15;
wire  s_37_16,  s_37_17,  s_37_18,   s_38_0,   s_38_1,   s_38_2;
wire   s_38_3,   s_38_4,   s_38_5,   s_38_6,   s_38_7,   s_38_8;
wire   s_38_9,  s_38_10,  s_38_11,  s_38_12,  s_38_13,  s_38_14;
wire  s_38_15,  s_38_16,  s_38_17,  s_38_18,  s_38_19,  s_38_20;
wire   s_39_0,   s_39_1,   s_39_2,   s_39_3,   s_39_4,   s_39_5;
wire   s_39_6,   s_39_7,   s_39_8,   s_39_9,  s_39_10,  s_39_11;
wire  s_39_12,  s_39_13,  s_39_14,  s_39_15,  s_39_16,  s_39_17;
wire  s_39_18,  s_39_19,   s_40_0,   s_40_1,   s_40_2,   s_40_3;
wire   s_40_4,   s_40_5,   s_40_6,   s_40_7,   s_40_8,   s_40_9;
wire  s_40_10,  s_40_11,  s_40_12,  s_40_13,  s_40_14,  s_40_15;
wire  s_40_16,  s_40_17,  s_40_18,  s_40_19,  s_40_20,  s_40_21;
wire   s_41_0,   s_41_1,   s_41_2,   s_41_3,   s_41_4,   s_41_5;
wire   s_41_6,   s_41_7,   s_41_8,   s_41_9,  s_41_10,  s_41_11;
wire  s_41_12,  s_41_13,  s_41_14,  s_41_15,  s_41_16,  s_41_17;
wire  s_41_18,  s_41_19,  s_41_20,   s_42_0,   s_42_1,   s_42_2;
wire   s_42_3,   s_42_4,   s_42_5,   s_42_6,   s_42_7,   s_42_8;
wire   s_42_9,  s_42_10,  s_42_11,  s_42_12,  s_42_13,  s_42_14;
wire  s_42_15,  s_42_16,  s_42_17,  s_42_18,  s_42_19,  s_42_20;
wire  s_42_21,  s_42_22,   s_43_0,   s_43_1,   s_43_2,   s_43_3;
wire   s_43_4,   s_43_5,   s_43_6,   s_43_7,   s_43_8,   s_43_9;
wire  s_43_10,  s_43_11,  s_43_12,  s_43_13,  s_43_14,  s_43_15;
wire  s_43_16,  s_43_17,  s_43_18,  s_43_19,  s_43_20,  s_43_21;
wire   s_44_0,   s_44_1,   s_44_2,   s_44_3,   s_44_4,   s_44_5;
wire   s_44_6,   s_44_7,   s_44_8,   s_44_9,  s_44_10,  s_44_11;
wire  s_44_12,  s_44_13,  s_44_14,  s_44_15,  s_44_16,  s_44_17;
wire  s_44_18,  s_44_19,  s_44_20,  s_44_21,  s_44_22,  s_44_23;
wire   s_45_0,   s_45_1,   s_45_2,   s_45_3,   s_45_4,   s_45_5;
wire   s_45_6,   s_45_7,   s_45_8,   s_45_9,  s_45_10,  s_45_11;
wire  s_45_12,  s_45_13,  s_45_14,  s_45_15,  s_45_16,  s_45_17;
wire  s_45_18,  s_45_19,  s_45_20,  s_45_21,  s_45_22,   s_46_0;
wire   s_46_1,   s_46_2,   s_46_3,   s_46_4,   s_46_5,   s_46_6;
wire   s_46_7,   s_46_8,   s_46_9,  s_46_10,  s_46_11,  s_46_12;
wire  s_46_13,  s_46_14,  s_46_15,  s_46_16,  s_46_17,  s_46_18;
wire  s_46_19,  s_46_20,  s_46_21,  s_46_22,  s_46_23,  s_46_24;
wire   s_47_0,   s_47_1,   s_47_2,   s_47_3,   s_47_4,   s_47_5;
wire   s_47_6,   s_47_7,   s_47_8,   s_47_9,  s_47_10,  s_47_11;
wire  s_47_12,  s_47_13,  s_47_14,  s_47_15,  s_47_16,  s_47_17;
wire  s_47_18,  s_47_19,  s_47_20,  s_47_21,  s_47_22,  s_47_23;
wire   s_48_0,   s_48_1,   s_48_2,   s_48_3,   s_48_4,   s_48_5;
wire   s_48_6,   s_48_7,   s_48_8,   s_48_9,  s_48_10,  s_48_11;
wire  s_48_12,  s_48_13,  s_48_14,  s_48_15,  s_48_16,  s_48_17;
wire  s_48_18,  s_48_19,  s_48_20,  s_48_21,  s_48_22,  s_48_23;
wire  s_48_24,  s_48_25,   s_49_0,   s_49_1,   s_49_2,   s_49_3;
wire   s_49_4,   s_49_5,   s_49_6,   s_49_7,   s_49_8,   s_49_9;
wire  s_49_10,  s_49_11,  s_49_12,  s_49_13,  s_49_14,  s_49_15;
wire  s_49_16,  s_49_17,  s_49_18,  s_49_19,  s_49_20,  s_49_21;
wire  s_49_22,  s_49_23,  s_49_24,   s_50_0,   s_50_1,   s_50_2;
wire   s_50_3,   s_50_4,   s_50_5,   s_50_6,   s_50_7,   s_50_8;
wire   s_50_9,  s_50_10,  s_50_11,  s_50_12,  s_50_13,  s_50_14;
wire  s_50_15,  s_50_16,  s_50_17,  s_50_18,  s_50_19,  s_50_20;
wire  s_50_21,  s_50_22,  s_50_23,  s_50_24,  s_50_25,  s_50_26;
wire   s_51_0,   s_51_1,   s_51_2,   s_51_3,   s_51_4,   s_51_5;
wire   s_51_6,   s_51_7,   s_51_8,   s_51_9,  s_51_10,  s_51_11;
wire  s_51_12,  s_51_13,  s_51_14,  s_51_15,  s_51_16,  s_51_17;
wire  s_51_18,  s_51_19,  s_51_20,  s_51_21,  s_51_22,  s_51_23;
wire  s_51_24,  s_51_25,   s_52_0,   s_52_1,   s_52_2,   s_52_3;
wire   s_52_4,   s_52_5,   s_52_6,   s_52_7,   s_52_8,   s_52_9;
wire  s_52_10,  s_52_11,  s_52_12,  s_52_13,  s_52_14,  s_52_15;
wire  s_52_16,  s_52_17,  s_52_18,  s_52_19,  s_52_20,  s_52_21;
wire  s_52_22,  s_52_23,  s_52_24,  s_52_25,  s_52_26,  s_52_27;
wire   s_53_0,   s_53_1,   s_53_2,   s_53_3,   s_53_4,   s_53_5;
wire   s_53_6,   s_53_7,   s_53_8,   s_53_9,  s_53_10,  s_53_11;
wire  s_53_12,  s_53_13,  s_53_14,  s_53_15,  s_53_16,  s_53_17;
wire  s_53_18,  s_53_19,  s_53_20,  s_53_21,  s_53_22,  s_53_23;
wire  s_53_24,  s_53_25,  s_53_26,   s_54_0,   s_54_1,   s_54_2;
wire   s_54_3,   s_54_4,   s_54_5,   s_54_6,   s_54_7,   s_54_8;
wire   s_54_9,  s_54_10,  s_54_11,  s_54_12,  s_54_13,  s_54_14;
wire  s_54_15,  s_54_16,  s_54_17,  s_54_18,  s_54_19,  s_54_20;
wire  s_54_21,  s_54_22,  s_54_23,  s_54_24,  s_54_25,  s_54_26;
wire  s_54_27,  s_54_28,   s_55_0,   s_55_1,   s_55_2,   s_55_3;
wire   s_55_4,   s_55_5,   s_55_6,   s_55_7,   s_55_8,   s_55_9;
wire  s_55_10,  s_55_11,  s_55_12,  s_55_13,  s_55_14,  s_55_15;
wire  s_55_16,  s_55_17,  s_55_18,  s_55_19,  s_55_20,  s_55_21;
wire  s_55_22,  s_55_23,  s_55_24,  s_55_25,  s_55_26,  s_55_27;
wire   s_56_0,   s_56_1,   s_56_2,   s_56_3,   s_56_4,   s_56_5;
wire   s_56_6,   s_56_7,   s_56_8,   s_56_9,  s_56_10,  s_56_11;
wire  s_56_12,  s_56_13,  s_56_14,  s_56_15,  s_56_16,  s_56_17;
wire  s_56_18,  s_56_19,  s_56_20,  s_56_21,  s_56_22,  s_56_23;
wire  s_56_24,  s_56_25,  s_56_26,  s_56_27,  s_56_28,  s_56_29;
wire   s_57_0,   s_57_1,   s_57_2,   s_57_3,   s_57_4,   s_57_5;
wire   s_57_6,   s_57_7,   s_57_8,   s_57_9,  s_57_10,  s_57_11;
wire  s_57_12,  s_57_13,  s_57_14,  s_57_15,  s_57_16,  s_57_17;
wire  s_57_18,  s_57_19,  s_57_20,  s_57_21,  s_57_22,  s_57_23;
wire  s_57_24,  s_57_25,  s_57_26,  s_57_27,  s_57_28,   s_58_0;
wire   s_58_1,   s_58_2,   s_58_3,   s_58_4,   s_58_5,   s_58_6;
wire   s_58_7,   s_58_8,   s_58_9,  s_58_10,  s_58_11,  s_58_12;
wire  s_58_13,  s_58_14,  s_58_15,  s_58_16,  s_58_17,  s_58_18;
wire  s_58_19,  s_58_20,  s_58_21,  s_58_22,  s_58_23,  s_58_24;
wire  s_58_25,  s_58_26,  s_58_27,  s_58_28,  s_58_29,  s_58_30;
wire   s_59_0,   s_59_1,   s_59_2,   s_59_3,   s_59_4,   s_59_5;
wire   s_59_6,   s_59_7,   s_59_8,   s_59_9,  s_59_10,  s_59_11;
wire  s_59_12,  s_59_13,  s_59_14,  s_59_15,  s_59_16,  s_59_17;
wire  s_59_18,  s_59_19,  s_59_20,  s_59_21,  s_59_22,  s_59_23;
wire  s_59_24,  s_59_25,  s_59_26,  s_59_27,  s_59_28,  s_59_29;
wire   s_60_0,   s_60_1,   s_60_2,   s_60_3,   s_60_4,   s_60_5;
wire   s_60_6,   s_60_7,   s_60_8,   s_60_9,  s_60_10,  s_60_11;
wire  s_60_12,  s_60_13,  s_60_14,  s_60_15,  s_60_16,  s_60_17;
wire  s_60_18,  s_60_19,  s_60_20,  s_60_21,  s_60_22,  s_60_23;
wire  s_60_24,  s_60_25,  s_60_26,  s_60_27,  s_60_28,  s_60_29;
wire  s_60_30,  s_60_31,   s_61_0,   s_61_1,   s_61_2,   s_61_3;
wire   s_61_4,   s_61_5,   s_61_6,   s_61_7,   s_61_8,   s_61_9;
wire  s_61_10,  s_61_11,  s_61_12,  s_61_13,  s_61_14,  s_61_15;
wire  s_61_16,  s_61_17,  s_61_18,  s_61_19,  s_61_20,  s_61_21;
wire  s_61_22,  s_61_23,  s_61_24,  s_61_25,  s_61_26,  s_61_27;
wire  s_61_28,  s_61_29,  s_61_30,   s_62_0,   s_62_1,   s_62_2;
wire   s_62_3,   s_62_4,   s_62_5,   s_62_6,   s_62_7,   s_62_8;
wire   s_62_9,  s_62_10,  s_62_11,  s_62_12,  s_62_13,  s_62_14;
wire  s_62_15,  s_62_16,  s_62_17,  s_62_18,  s_62_19,  s_62_20;
wire  s_62_21,  s_62_22,  s_62_23,  s_62_24,  s_62_25,  s_62_26;
wire  s_62_27,  s_62_28,  s_62_29,  s_62_30,  s_62_31,  s_62_32;
wire   s_63_0,   s_63_1,   s_63_2,   s_63_3,   s_63_4,   s_63_5;
wire   s_63_6,   s_63_7,   s_63_8,   s_63_9,  s_63_10,  s_63_11;
wire  s_63_12,  s_63_13,  s_63_14,  s_63_15,  s_63_16,  s_63_17;
wire  s_63_18,  s_63_19,  s_63_20,  s_63_21,  s_63_22,  s_63_23;
wire  s_63_24,  s_63_25,  s_63_26,  s_63_27,  s_63_28,  s_63_29;
wire  s_63_30,  s_63_31,   s_64_0,   s_64_1,   s_64_2,   s_64_3;
wire   s_64_4,   s_64_5,   s_64_6,   s_64_7,   s_64_8,   s_64_9;
wire  s_64_10,  s_64_11,  s_64_12,  s_64_13,  s_64_14,  s_64_15;
wire  s_64_16,  s_64_17,  s_64_18,  s_64_19,  s_64_20,  s_64_21;
wire  s_64_22,  s_64_23,  s_64_24,  s_64_25,  s_64_26,  s_64_27;
wire  s_64_28,  s_64_29,  s_64_30,  s_64_31,  s_64_32,  s_64_33;
wire   s_65_0,   s_65_1,   s_65_2,   s_65_3,   s_65_4,   s_65_5;
wire   s_65_6,   s_65_7,   s_65_8,   s_65_9,  s_65_10,  s_65_11;
wire  s_65_12,  s_65_13,  s_65_14,  s_65_15,  s_65_16,  s_65_17;
wire  s_65_18,  s_65_19,  s_65_20,  s_65_21,  s_65_22,  s_65_23;
wire  s_65_24,  s_65_25,  s_65_26,  s_65_27,  s_65_28,  s_65_29;
wire  s_65_30,  s_65_31,  s_65_32,   s_66_0,   s_66_1,   s_66_2;
wire   s_66_3,   s_66_4,   s_66_5,   s_66_6,   s_66_7,   s_66_8;
wire   s_66_9,  s_66_10,  s_66_11,  s_66_12,  s_66_13,  s_66_14;
wire  s_66_15,  s_66_16,  s_66_17,  s_66_18,  s_66_19,  s_66_20;
wire  s_66_21,  s_66_22,  s_66_23,  s_66_24,  s_66_25,  s_66_26;
wire  s_66_27,  s_66_28,  s_66_29,  s_66_30,  s_66_31,  s_66_32;
wire  s_66_33,  s_66_34,   s_67_0,   s_67_1,   s_67_2,   s_67_3;
wire   s_67_4,   s_67_5,   s_67_6,   s_67_7,   s_67_8,   s_67_9;
wire  s_67_10,  s_67_11,  s_67_12,  s_67_13,  s_67_14,  s_67_15;
wire  s_67_16,  s_67_17,  s_67_18,  s_67_19,  s_67_20,  s_67_21;
wire  s_67_22,  s_67_23,  s_67_24,  s_67_25,  s_67_26,  s_67_27;
wire  s_67_28,  s_67_29,  s_67_30,  s_67_31,  s_67_32,  s_67_33;
wire   s_68_0,   s_68_1,   s_68_2,   s_68_3,   s_68_4,   s_68_5;
wire   s_68_6,   s_68_7,   s_68_8,   s_68_9,  s_68_10,  s_68_11;
wire  s_68_12,  s_68_13,  s_68_14,  s_68_15,  s_68_16,  s_68_17;
wire  s_68_18,  s_68_19,  s_68_20,  s_68_21,  s_68_22,  s_68_23;
wire  s_68_24,  s_68_25,  s_68_26,  s_68_27,  s_68_28,  s_68_29;
wire  s_68_30,  s_68_31,  s_68_32,  s_68_33,  s_68_34,  s_68_35;
wire   s_69_0,   s_69_1,   s_69_2,   s_69_3,   s_69_4,   s_69_5;
wire   s_69_6,   s_69_7,   s_69_8,   s_69_9,  s_69_10,  s_69_11;
wire  s_69_12,  s_69_13,  s_69_14,  s_69_15,  s_69_16,  s_69_17;
wire  s_69_18,  s_69_19,  s_69_20,  s_69_21,  s_69_22,  s_69_23;
wire  s_69_24,  s_69_25,  s_69_26,  s_69_27,  s_69_28,  s_69_29;
wire  s_69_30,  s_69_31,  s_69_32,  s_69_33,  s_69_34,   s_70_0;
wire   s_70_1,   s_70_2,   s_70_3,   s_70_4,   s_70_5,   s_70_6;
wire   s_70_7,   s_70_8,   s_70_9,  s_70_10,  s_70_11,  s_70_12;
wire  s_70_13,  s_70_14,  s_70_15,  s_70_16,  s_70_17,  s_70_18;
wire  s_70_19,  s_70_20,  s_70_21,  s_70_22,  s_70_23,  s_70_24;
wire  s_70_25,  s_70_26,  s_70_27,  s_70_28,  s_70_29,  s_70_30;
wire  s_70_31,  s_70_32,  s_70_33,  s_70_34,  s_70_35,  s_70_36;
wire   s_71_0,   s_71_1,   s_71_2,   s_71_3,   s_71_4,   s_71_5;
wire   s_71_6,   s_71_7,   s_71_8,   s_71_9,  s_71_10,  s_71_11;
wire  s_71_12,  s_71_13,  s_71_14,  s_71_15,  s_71_16,  s_71_17;
wire  s_71_18,  s_71_19,  s_71_20,  s_71_21,  s_71_22,  s_71_23;
wire  s_71_24,  s_71_25,  s_71_26,  s_71_27,  s_71_28,  s_71_29;
wire  s_71_30,  s_71_31,  s_71_32,  s_71_33,  s_71_34,  s_71_35;
wire   s_72_0,   s_72_1,   s_72_2,   s_72_3,   s_72_4,   s_72_5;
wire   s_72_6,   s_72_7,   s_72_8,   s_72_9,  s_72_10,  s_72_11;
wire  s_72_12,  s_72_13,  s_72_14,  s_72_15,  s_72_16,  s_72_17;
wire  s_72_18,  s_72_19,  s_72_20,  s_72_21,  s_72_22,  s_72_23;
wire  s_72_24,  s_72_25,  s_72_26,  s_72_27,  s_72_28,  s_72_29;
wire  s_72_30,  s_72_31,  s_72_32,  s_72_33,  s_72_34,  s_72_35;
wire  s_72_36,  s_72_37,   s_73_0,   s_73_1,   s_73_2,   s_73_3;
wire   s_73_4,   s_73_5,   s_73_6,   s_73_7,   s_73_8,   s_73_9;
wire  s_73_10,  s_73_11,  s_73_12,  s_73_13,  s_73_14,  s_73_15;
wire  s_73_16,  s_73_17,  s_73_18,  s_73_19,  s_73_20,  s_73_21;
wire  s_73_22,  s_73_23,  s_73_24,  s_73_25,  s_73_26,  s_73_27;
wire  s_73_28,  s_73_29,  s_73_30,  s_73_31,  s_73_32,  s_73_33;
wire  s_73_34,  s_73_35,  s_73_36,   s_74_0,   s_74_1,   s_74_2;
wire   s_74_3,   s_74_4,   s_74_5,   s_74_6,   s_74_7,   s_74_8;
wire   s_74_9,  s_74_10,  s_74_11,  s_74_12,  s_74_13,  s_74_14;
wire  s_74_15,  s_74_16,  s_74_17,  s_74_18,  s_74_19,  s_74_20;
wire  s_74_21,  s_74_22,  s_74_23,  s_74_24,  s_74_25,  s_74_26;
wire  s_74_27,  s_74_28,  s_74_29,  s_74_30,  s_74_31,  s_74_32;
wire  s_74_33,  s_74_34,  s_74_35,  s_74_36,  s_74_37,  s_74_38;
wire   s_75_0,   s_75_1,   s_75_2,   s_75_3,   s_75_4,   s_75_5;
wire   s_75_6,   s_75_7,   s_75_8,   s_75_9,  s_75_10,  s_75_11;
wire  s_75_12,  s_75_13,  s_75_14,  s_75_15,  s_75_16,  s_75_17;
wire  s_75_18,  s_75_19,  s_75_20,  s_75_21,  s_75_22,  s_75_23;
wire  s_75_24,  s_75_25,  s_75_26,  s_75_27,  s_75_28,  s_75_29;
wire  s_75_30,  s_75_31,  s_75_32,  s_75_33,  s_75_34,  s_75_35;
wire  s_75_36,  s_75_37,   s_76_0,   s_76_1,   s_76_2,   s_76_3;
wire   s_76_4,   s_76_5,   s_76_6,   s_76_7,   s_76_8,   s_76_9;
wire  s_76_10,  s_76_11,  s_76_12,  s_76_13,  s_76_14,  s_76_15;
wire  s_76_16,  s_76_17,  s_76_18,  s_76_19,  s_76_20,  s_76_21;
wire  s_76_22,  s_76_23,  s_76_24,  s_76_25,  s_76_26,  s_76_27;
wire  s_76_28,  s_76_29,  s_76_30,  s_76_31,  s_76_32,  s_76_33;
wire  s_76_34,  s_76_35,  s_76_36,  s_76_37,  s_76_38,  s_76_39;
wire   s_77_0,   s_77_1,   s_77_2,   s_77_3,   s_77_4,   s_77_5;
wire   s_77_6,   s_77_7,   s_77_8,   s_77_9,  s_77_10,  s_77_11;
wire  s_77_12,  s_77_13,  s_77_14,  s_77_15,  s_77_16,  s_77_17;
wire  s_77_18,  s_77_19,  s_77_20,  s_77_21,  s_77_22,  s_77_23;
wire  s_77_24,  s_77_25,  s_77_26,  s_77_27,  s_77_28,  s_77_29;
wire  s_77_30,  s_77_31,  s_77_32,  s_77_33,  s_77_34,  s_77_35;
wire  s_77_36,  s_77_37,  s_77_38,   s_78_0,   s_78_1,   s_78_2;
wire   s_78_3,   s_78_4,   s_78_5,   s_78_6,   s_78_7,   s_78_8;
wire   s_78_9,  s_78_10,  s_78_11,  s_78_12,  s_78_13,  s_78_14;
wire  s_78_15,  s_78_16,  s_78_17,  s_78_18,  s_78_19,  s_78_20;
wire  s_78_21,  s_78_22,  s_78_23,  s_78_24,  s_78_25,  s_78_26;
wire  s_78_27,  s_78_28,  s_78_29,  s_78_30,  s_78_31,  s_78_32;
wire  s_78_33,  s_78_34,  s_78_35,  s_78_36,  s_78_37,  s_78_38;
wire  s_78_39,  s_78_40,   s_79_0,   s_79_1,   s_79_2,   s_79_3;
wire   s_79_4,   s_79_5,   s_79_6,   s_79_7,   s_79_8,   s_79_9;
wire  s_79_10,  s_79_11,  s_79_12,  s_79_13,  s_79_14,  s_79_15;
wire  s_79_16,  s_79_17,  s_79_18,  s_79_19,  s_79_20,  s_79_21;
wire  s_79_22,  s_79_23,  s_79_24,  s_79_25,  s_79_26,  s_79_27;
wire  s_79_28,  s_79_29,  s_79_30,  s_79_31,  s_79_32,  s_79_33;
wire  s_79_34,  s_79_35,  s_79_36,  s_79_37,  s_79_38,  s_79_39;
wire   s_80_0,   s_80_1,   s_80_2,   s_80_3,   s_80_4,   s_80_5;
wire   s_80_6,   s_80_7,   s_80_8,   s_80_9,  s_80_10,  s_80_11;
wire  s_80_12,  s_80_13,  s_80_14,  s_80_15,  s_80_16,  s_80_17;
wire  s_80_18,  s_80_19,  s_80_20,  s_80_21,  s_80_22,  s_80_23;
wire  s_80_24,  s_80_25,  s_80_26,  s_80_27,  s_80_28,  s_80_29;
wire  s_80_30,  s_80_31,  s_80_32,  s_80_33,  s_80_34,  s_80_35;
wire  s_80_36,  s_80_37,  s_80_38,  s_80_39,  s_80_40,  s_80_41;
wire   s_81_0,   s_81_1,   s_81_2,   s_81_3,   s_81_4,   s_81_5;
wire   s_81_6,   s_81_7,   s_81_8,   s_81_9,  s_81_10,  s_81_11;
wire  s_81_12,  s_81_13,  s_81_14,  s_81_15,  s_81_16,  s_81_17;
wire  s_81_18,  s_81_19,  s_81_20,  s_81_21,  s_81_22,  s_81_23;
wire  s_81_24,  s_81_25,  s_81_26,  s_81_27,  s_81_28,  s_81_29;
wire  s_81_30,  s_81_31,  s_81_32,  s_81_33,  s_81_34,  s_81_35;
wire  s_81_36,  s_81_37,  s_81_38,  s_81_39,  s_81_40,   s_82_0;
wire   s_82_1,   s_82_2,   s_82_3,   s_82_4,   s_82_5,   s_82_6;
wire   s_82_7,   s_82_8,   s_82_9,  s_82_10,  s_82_11,  s_82_12;
wire  s_82_13,  s_82_14,  s_82_15,  s_82_16,  s_82_17,  s_82_18;
wire  s_82_19,  s_82_20,  s_82_21,  s_82_22,  s_82_23,  s_82_24;
wire  s_82_25,  s_82_26,  s_82_27,  s_82_28,  s_82_29,  s_82_30;
wire  s_82_31,  s_82_32,  s_82_33,  s_82_34,  s_82_35,  s_82_36;
wire  s_82_37,  s_82_38,  s_82_39,  s_82_40,  s_82_41,  s_82_42;
wire   s_83_0,   s_83_1,   s_83_2,   s_83_3,   s_83_4,   s_83_5;
wire   s_83_6,   s_83_7,   s_83_8,   s_83_9,  s_83_10,  s_83_11;
wire  s_83_12,  s_83_13,  s_83_14,  s_83_15,  s_83_16,  s_83_17;
wire  s_83_18,  s_83_19,  s_83_20,  s_83_21,  s_83_22,  s_83_23;
wire  s_83_24,  s_83_25,  s_83_26,  s_83_27,  s_83_28,  s_83_29;
wire  s_83_30,  s_83_31,  s_83_32,  s_83_33,  s_83_34,  s_83_35;
wire  s_83_36,  s_83_37,  s_83_38,  s_83_39,  s_83_40,  s_83_41;
wire   s_84_0,   s_84_1,   s_84_2,   s_84_3,   s_84_4,   s_84_5;
wire   s_84_6,   s_84_7,   s_84_8,   s_84_9,  s_84_10,  s_84_11;
wire  s_84_12,  s_84_13,  s_84_14,  s_84_15,  s_84_16,  s_84_17;
wire  s_84_18,  s_84_19,  s_84_20,  s_84_21,  s_84_22,  s_84_23;
wire  s_84_24,  s_84_25,  s_84_26,  s_84_27,  s_84_28,  s_84_29;
wire  s_84_30,  s_84_31,  s_84_32,  s_84_33,  s_84_34,  s_84_35;
wire  s_84_36,  s_84_37,  s_84_38,  s_84_39,  s_84_40,  s_84_41;
wire  s_84_42,  s_84_43,   s_85_0,   s_85_1,   s_85_2,   s_85_3;
wire   s_85_4,   s_85_5,   s_85_6,   s_85_7,   s_85_8,   s_85_9;
wire  s_85_10,  s_85_11,  s_85_12,  s_85_13,  s_85_14,  s_85_15;
wire  s_85_16,  s_85_17,  s_85_18,  s_85_19,  s_85_20,  s_85_21;
wire  s_85_22,  s_85_23,  s_85_24,  s_85_25,  s_85_26,  s_85_27;
wire  s_85_28,  s_85_29,  s_85_30,  s_85_31,  s_85_32,  s_85_33;
wire  s_85_34,  s_85_35,  s_85_36,  s_85_37,  s_85_38,  s_85_39;
wire  s_85_40,  s_85_41,  s_85_42,   s_86_0,   s_86_1,   s_86_2;
wire   s_86_3,   s_86_4,   s_86_5,   s_86_6,   s_86_7,   s_86_8;
wire   s_86_9,  s_86_10,  s_86_11,  s_86_12,  s_86_13,  s_86_14;
wire  s_86_15,  s_86_16,  s_86_17,  s_86_18,  s_86_19,  s_86_20;
wire  s_86_21,  s_86_22,  s_86_23,  s_86_24,  s_86_25,  s_86_26;
wire  s_86_27,  s_86_28,  s_86_29,  s_86_30,  s_86_31,  s_86_32;
wire  s_86_33,  s_86_34,  s_86_35,  s_86_36,  s_86_37,  s_86_38;
wire  s_86_39,  s_86_40,  s_86_41,  s_86_42,  s_86_43,  s_86_44;
wire   s_87_0,   s_87_1,   s_87_2,   s_87_3,   s_87_4,   s_87_5;
wire   s_87_6,   s_87_7,   s_87_8,   s_87_9,  s_87_10,  s_87_11;
wire  s_87_12,  s_87_13,  s_87_14,  s_87_15,  s_87_16,  s_87_17;
wire  s_87_18,  s_87_19,  s_87_20,  s_87_21,  s_87_22,  s_87_23;
wire  s_87_24,  s_87_25,  s_87_26,  s_87_27,  s_87_28,  s_87_29;
wire  s_87_30,  s_87_31,  s_87_32,  s_87_33,  s_87_34,  s_87_35;
wire  s_87_36,  s_87_37,  s_87_38,  s_87_39,  s_87_40,  s_87_41;
wire  s_87_42,  s_87_43,   s_88_0,   s_88_1,   s_88_2,   s_88_3;
wire   s_88_4,   s_88_5,   s_88_6,   s_88_7,   s_88_8,   s_88_9;
wire  s_88_10,  s_88_11,  s_88_12,  s_88_13,  s_88_14,  s_88_15;
wire  s_88_16,  s_88_17,  s_88_18,  s_88_19,  s_88_20,  s_88_21;
wire  s_88_22,  s_88_23,  s_88_24,  s_88_25,  s_88_26,  s_88_27;
wire  s_88_28,  s_88_29,  s_88_30,  s_88_31,  s_88_32,  s_88_33;
wire  s_88_34,  s_88_35,  s_88_36,  s_88_37,  s_88_38,  s_88_39;
wire  s_88_40,  s_88_41,  s_88_42,  s_88_43,  s_88_44,  s_88_45;
wire   s_89_0,   s_89_1,   s_89_2,   s_89_3,   s_89_4,   s_89_5;
wire   s_89_6,   s_89_7,   s_89_8,   s_89_9,  s_89_10,  s_89_11;
wire  s_89_12,  s_89_13,  s_89_14,  s_89_15,  s_89_16,  s_89_17;
wire  s_89_18,  s_89_19,  s_89_20,  s_89_21,  s_89_22,  s_89_23;
wire  s_89_24,  s_89_25,  s_89_26,  s_89_27,  s_89_28,  s_89_29;
wire  s_89_30,  s_89_31,  s_89_32,  s_89_33,  s_89_34,  s_89_35;
wire  s_89_36,  s_89_37,  s_89_38,  s_89_39,  s_89_40,  s_89_41;
wire  s_89_42,  s_89_43,  s_89_44,   s_90_0,   s_90_1,   s_90_2;
wire   s_90_3,   s_90_4,   s_90_5,   s_90_6,   s_90_7,   s_90_8;
wire   s_90_9,  s_90_10,  s_90_11,  s_90_12,  s_90_13,  s_90_14;
wire  s_90_15,  s_90_16,  s_90_17,  s_90_18,  s_90_19,  s_90_20;
wire  s_90_21,  s_90_22,  s_90_23,  s_90_24,  s_90_25,  s_90_26;
wire  s_90_27,  s_90_28,  s_90_29,  s_90_30,  s_90_31,  s_90_32;
wire  s_90_33,  s_90_34,  s_90_35,  s_90_36,  s_90_37,  s_90_38;
wire  s_90_39,  s_90_40,  s_90_41,  s_90_42,  s_90_43,  s_90_44;
wire  s_90_45,  s_90_46,   s_91_0,   s_91_1,   s_91_2,   s_91_3;
wire   s_91_4,   s_91_5,   s_91_6,   s_91_7,   s_91_8,   s_91_9;
wire  s_91_10,  s_91_11,  s_91_12,  s_91_13,  s_91_14,  s_91_15;
wire  s_91_16,  s_91_17,  s_91_18,  s_91_19,  s_91_20,  s_91_21;
wire  s_91_22,  s_91_23,  s_91_24,  s_91_25,  s_91_26,  s_91_27;
wire  s_91_28,  s_91_29,  s_91_30,  s_91_31,  s_91_32,  s_91_33;
wire  s_91_34,  s_91_35,  s_91_36,  s_91_37,  s_91_38,  s_91_39;
wire  s_91_40,  s_91_41,  s_91_42,  s_91_43,  s_91_44,  s_91_45;
wire   s_92_0,   s_92_1,   s_92_2,   s_92_3,   s_92_4,   s_92_5;
wire   s_92_6,   s_92_7,   s_92_8,   s_92_9,  s_92_10,  s_92_11;
wire  s_92_12,  s_92_13,  s_92_14,  s_92_15,  s_92_16,  s_92_17;
wire  s_92_18,  s_92_19,  s_92_20,  s_92_21,  s_92_22,  s_92_23;
wire  s_92_24,  s_92_25,  s_92_26,  s_92_27,  s_92_28,  s_92_29;
wire  s_92_30,  s_92_31,  s_92_32,  s_92_33,  s_92_34,  s_92_35;
wire  s_92_36,  s_92_37,  s_92_38,  s_92_39,  s_92_40,  s_92_41;
wire  s_92_42,  s_92_43,  s_92_44,  s_92_45,  s_92_46,  s_92_47;
wire   s_93_0,   s_93_1,   s_93_2,   s_93_3,   s_93_4,   s_93_5;
wire   s_93_6,   s_93_7,   s_93_8,   s_93_9,  s_93_10,  s_93_11;
wire  s_93_12,  s_93_13,  s_93_14,  s_93_15,  s_93_16,  s_93_17;
wire  s_93_18,  s_93_19,  s_93_20,  s_93_21,  s_93_22,  s_93_23;
wire  s_93_24,  s_93_25,  s_93_26,  s_93_27,  s_93_28,  s_93_29;
wire  s_93_30,  s_93_31,  s_93_32,  s_93_33,  s_93_34,  s_93_35;
wire  s_93_36,  s_93_37,  s_93_38,  s_93_39,  s_93_40,  s_93_41;
wire  s_93_42,  s_93_43,  s_93_44,  s_93_45,  s_93_46,   s_94_0;
wire   s_94_1,   s_94_2,   s_94_3,   s_94_4,   s_94_5,   s_94_6;
wire   s_94_7,   s_94_8,   s_94_9,  s_94_10,  s_94_11,  s_94_12;
wire  s_94_13,  s_94_14,  s_94_15,  s_94_16,  s_94_17,  s_94_18;
wire  s_94_19,  s_94_20,  s_94_21,  s_94_22,  s_94_23,  s_94_24;
wire  s_94_25,  s_94_26,  s_94_27,  s_94_28,  s_94_29,  s_94_30;
wire  s_94_31,  s_94_32,  s_94_33,  s_94_34,  s_94_35,  s_94_36;
wire  s_94_37,  s_94_38,  s_94_39,  s_94_40,  s_94_41,  s_94_42;
wire  s_94_43,  s_94_44,  s_94_45,  s_94_46,  s_94_47,  s_94_48;
wire   s_95_0,   s_95_1,   s_95_2,   s_95_3,   s_95_4,   s_95_5;
wire   s_95_6,   s_95_7,   s_95_8,   s_95_9,  s_95_10,  s_95_11;
wire  s_95_12,  s_95_13,  s_95_14,  s_95_15,  s_95_16,  s_95_17;
wire  s_95_18,  s_95_19,  s_95_20,  s_95_21,  s_95_22,  s_95_23;
wire  s_95_24,  s_95_25,  s_95_26,  s_95_27,  s_95_28,  s_95_29;
wire  s_95_30,  s_95_31,  s_95_32,  s_95_33,  s_95_34,  s_95_35;
wire  s_95_36,  s_95_37,  s_95_38,  s_95_39,  s_95_40,  s_95_41;
wire  s_95_42,  s_95_43,  s_95_44,  s_95_45,  s_95_46,  s_95_47;
wire   s_96_0,   s_96_1,   s_96_2,   s_96_3,   s_96_4,   s_96_5;
wire   s_96_6,   s_96_7,   s_96_8,   s_96_9,  s_96_10,  s_96_11;
wire  s_96_12,  s_96_13,  s_96_14,  s_96_15,  s_96_16,  s_96_17;
wire  s_96_18,  s_96_19,  s_96_20,  s_96_21,  s_96_22,  s_96_23;
wire  s_96_24,  s_96_25,  s_96_26,  s_96_27,  s_96_28,  s_96_29;
wire  s_96_30,  s_96_31,  s_96_32,  s_96_33,  s_96_34,  s_96_35;
wire  s_96_36,  s_96_37,  s_96_38,  s_96_39,  s_96_40,  s_96_41;
wire  s_96_42,  s_96_43,  s_96_44,  s_96_45,  s_96_46,  s_96_47;
wire  s_96_48,  s_96_49,   s_97_0,   s_97_1,   s_97_2,   s_97_3;
wire   s_97_4,   s_97_5,   s_97_6,   s_97_7,   s_97_8,   s_97_9;
wire  s_97_10,  s_97_11,  s_97_12,  s_97_13,  s_97_14,  s_97_15;
wire  s_97_16,  s_97_17,  s_97_18,  s_97_19,  s_97_20,  s_97_21;
wire  s_97_22,  s_97_23,  s_97_24,  s_97_25,  s_97_26,  s_97_27;
wire  s_97_28,  s_97_29,  s_97_30,  s_97_31,  s_97_32,  s_97_33;
wire  s_97_34,  s_97_35,  s_97_36,  s_97_37,  s_97_38,  s_97_39;
wire  s_97_40,  s_97_41,  s_97_42,  s_97_43,  s_97_44,  s_97_45;
wire  s_97_46,  s_97_47,  s_97_48,   s_98_0,   s_98_1,   s_98_2;
wire   s_98_3,   s_98_4,   s_98_5,   s_98_6,   s_98_7,   s_98_8;
wire   s_98_9,  s_98_10,  s_98_11,  s_98_12,  s_98_13,  s_98_14;
wire  s_98_15,  s_98_16,  s_98_17,  s_98_18,  s_98_19,  s_98_20;
wire  s_98_21,  s_98_22,  s_98_23,  s_98_24,  s_98_25,  s_98_26;
wire  s_98_27,  s_98_28,  s_98_29,  s_98_30,  s_98_31,  s_98_32;
wire  s_98_33,  s_98_34,  s_98_35,  s_98_36,  s_98_37,  s_98_38;
wire  s_98_39,  s_98_40,  s_98_41,  s_98_42,  s_98_43,  s_98_44;
wire  s_98_45,  s_98_46,  s_98_47,  s_98_48,  s_98_49,  s_98_50;
wire   s_99_0,   s_99_1,   s_99_2,   s_99_3,   s_99_4,   s_99_5;
wire   s_99_6,   s_99_7,   s_99_8,   s_99_9,  s_99_10,  s_99_11;
wire  s_99_12,  s_99_13,  s_99_14,  s_99_15,  s_99_16,  s_99_17;
wire  s_99_18,  s_99_19,  s_99_20,  s_99_21,  s_99_22,  s_99_23;
wire  s_99_24,  s_99_25,  s_99_26,  s_99_27,  s_99_28,  s_99_29;
wire  s_99_30,  s_99_31,  s_99_32,  s_99_33,  s_99_34,  s_99_35;
wire  s_99_36,  s_99_37,  s_99_38,  s_99_39,  s_99_40,  s_99_41;
wire  s_99_42,  s_99_43,  s_99_44,  s_99_45,  s_99_46,  s_99_47;
wire  s_99_48,  s_99_49,  s_100_0,  s_100_1,  s_100_2,  s_100_3;
wire  s_100_4,  s_100_5,  s_100_6,  s_100_7,  s_100_8,  s_100_9;
wire s_100_10, s_100_11, s_100_12, s_100_13, s_100_14, s_100_15;
wire s_100_16, s_100_17, s_100_18, s_100_19, s_100_20, s_100_21;
wire s_100_22, s_100_23, s_100_24, s_100_25, s_100_26, s_100_27;
wire s_100_28, s_100_29, s_100_30, s_100_31, s_100_32, s_100_33;
wire s_100_34, s_100_35, s_100_36, s_100_37, s_100_38, s_100_39;
wire s_100_40, s_100_41, s_100_42, s_100_43, s_100_44, s_100_45;
wire s_100_46, s_100_47, s_100_48, s_100_49, s_100_50, s_100_51;
wire  s_101_0,  s_101_1,  s_101_2,  s_101_3,  s_101_4,  s_101_5;
wire  s_101_6,  s_101_7,  s_101_8,  s_101_9, s_101_10, s_101_11;
wire s_101_12, s_101_13, s_101_14, s_101_15, s_101_16, s_101_17;
wire s_101_18, s_101_19, s_101_20, s_101_21, s_101_22, s_101_23;
wire s_101_24, s_101_25, s_101_26, s_101_27, s_101_28, s_101_29;
wire s_101_30, s_101_31, s_101_32, s_101_33, s_101_34, s_101_35;
wire s_101_36, s_101_37, s_101_38, s_101_39, s_101_40, s_101_41;
wire s_101_42, s_101_43, s_101_44, s_101_45, s_101_46, s_101_47;
wire s_101_48, s_101_49, s_101_50,  s_102_0,  s_102_1,  s_102_2;
wire  s_102_3,  s_102_4,  s_102_5,  s_102_6,  s_102_7,  s_102_8;
wire  s_102_9, s_102_10, s_102_11, s_102_12, s_102_13, s_102_14;
wire s_102_15, s_102_16, s_102_17, s_102_18, s_102_19, s_102_20;
wire s_102_21, s_102_22, s_102_23, s_102_24, s_102_25, s_102_26;
wire s_102_27, s_102_28, s_102_29, s_102_30, s_102_31, s_102_32;
wire s_102_33, s_102_34, s_102_35, s_102_36, s_102_37, s_102_38;
wire s_102_39, s_102_40, s_102_41, s_102_42, s_102_43, s_102_44;
wire s_102_45, s_102_46, s_102_47, s_102_48, s_102_49, s_102_50;
wire s_102_51, s_102_52,  s_103_0,  s_103_1,  s_103_2,  s_103_3;
wire  s_103_4,  s_103_5,  s_103_6,  s_103_7,  s_103_8,  s_103_9;
wire s_103_10, s_103_11, s_103_12, s_103_13, s_103_14, s_103_15;
wire s_103_16, s_103_17, s_103_18, s_103_19, s_103_20, s_103_21;
wire s_103_22, s_103_23, s_103_24, s_103_25, s_103_26, s_103_27;
wire s_103_28, s_103_29, s_103_30, s_103_31, s_103_32, s_103_33;
wire s_103_34, s_103_35, s_103_36, s_103_37, s_103_38, s_103_39;
wire s_103_40, s_103_41, s_103_42, s_103_43, s_103_44, s_103_45;
wire s_103_46, s_103_47, s_103_48, s_103_49, s_103_50, s_103_51;
wire  s_104_0,  s_104_1,  s_104_2,  s_104_3,  s_104_4,  s_104_5;
wire  s_104_6,  s_104_7,  s_104_8,  s_104_9, s_104_10, s_104_11;
wire s_104_12, s_104_13, s_104_14, s_104_15, s_104_16, s_104_17;
wire s_104_18, s_104_19, s_104_20, s_104_21, s_104_22, s_104_23;
wire s_104_24, s_104_25, s_104_26, s_104_27, s_104_28, s_104_29;
wire s_104_30, s_104_31, s_104_32, s_104_33, s_104_34, s_104_35;
wire s_104_36, s_104_37, s_104_38, s_104_39, s_104_40, s_104_41;
wire s_104_42, s_104_43, s_104_44, s_104_45, s_104_46, s_104_47;
wire s_104_48, s_104_49, s_104_50, s_104_51, s_104_52, s_104_53;
wire  s_105_0,  s_105_1,  s_105_2,  s_105_3,  s_105_4,  s_105_5;
wire  s_105_6,  s_105_7,  s_105_8,  s_105_9, s_105_10, s_105_11;
wire s_105_12, s_105_13, s_105_14, s_105_15, s_105_16, s_105_17;
wire s_105_18, s_105_19, s_105_20, s_105_21, s_105_22, s_105_23;
wire s_105_24, s_105_25, s_105_26, s_105_27, s_105_28, s_105_29;
wire s_105_30, s_105_31, s_105_32, s_105_33, s_105_34, s_105_35;
wire s_105_36, s_105_37, s_105_38, s_105_39, s_105_40, s_105_41;
wire s_105_42, s_105_43, s_105_44, s_105_45, s_105_46, s_105_47;
wire s_105_48, s_105_49, s_105_50, s_105_51, s_105_52,  s_106_0;
wire  s_106_1,  s_106_2,  s_106_3,  s_106_4,  s_106_5,  s_106_6;
wire  s_106_7,  s_106_8,  s_106_9, s_106_10, s_106_11, s_106_12;
wire s_106_13, s_106_14, s_106_15, s_106_16, s_106_17, s_106_18;
wire s_106_19, s_106_20, s_106_21, s_106_22, s_106_23, s_106_24;
wire s_106_25, s_106_26, s_106_27, s_106_28, s_106_29, s_106_30;
wire s_106_31, s_106_32, s_106_33, s_106_34, s_106_35, s_106_36;
wire s_106_37, s_106_38, s_106_39, s_106_40, s_106_41, s_106_42;
wire s_106_43, s_106_44, s_106_45, s_106_46, s_106_47, s_106_48;
wire s_106_49, s_106_50, s_106_51, s_106_52, s_106_53, s_106_54;
wire  s_107_0,  s_107_1,  s_107_2,  s_107_3,  s_107_4,  s_107_5;
wire  s_107_6,  s_107_7,  s_107_8,  s_107_9, s_107_10, s_107_11;
wire s_107_12, s_107_13, s_107_14, s_107_15, s_107_16, s_107_17;
wire s_107_18, s_107_19, s_107_20, s_107_21, s_107_22, s_107_23;
wire s_107_24, s_107_25, s_107_26, s_107_27, s_107_28, s_107_29;
wire s_107_30, s_107_31, s_107_32, s_107_33, s_107_34, s_107_35;
wire s_107_36, s_107_37, s_107_38, s_107_39, s_107_40, s_107_41;
wire s_107_42, s_107_43, s_107_44, s_107_45, s_107_46, s_107_47;
wire s_107_48, s_107_49, s_107_50, s_107_51, s_107_52, s_107_53;
wire  s_108_0,  s_108_1,  s_108_2,  s_108_3,  s_108_4,  s_108_5;
wire  s_108_6,  s_108_7,  s_108_8,  s_108_9, s_108_10, s_108_11;
wire s_108_12, s_108_13, s_108_14, s_108_15, s_108_16, s_108_17;
wire s_108_18, s_108_19, s_108_20, s_108_21, s_108_22, s_108_23;
wire s_108_24, s_108_25, s_108_26, s_108_27, s_108_28, s_108_29;
wire s_108_30, s_108_31, s_108_32, s_108_33, s_108_34, s_108_35;
wire s_108_36, s_108_37, s_108_38, s_108_39, s_108_40, s_108_41;
wire s_108_42, s_108_43, s_108_44, s_108_45, s_108_46, s_108_47;
wire s_108_48, s_108_49, s_108_50, s_108_51, s_108_52, s_108_53;
wire s_108_54, s_108_55,  s_109_0,  s_109_1,  s_109_2,  s_109_3;
wire  s_109_4,  s_109_5,  s_109_6,  s_109_7,  s_109_8,  s_109_9;
wire s_109_10, s_109_11, s_109_12, s_109_13, s_109_14, s_109_15;
wire s_109_16, s_109_17, s_109_18, s_109_19, s_109_20, s_109_21;
wire s_109_22, s_109_23, s_109_24, s_109_25, s_109_26, s_109_27;
wire s_109_28, s_109_29, s_109_30, s_109_31, s_109_32, s_109_33;
wire s_109_34, s_109_35, s_109_36, s_109_37, s_109_38, s_109_39;
wire s_109_40, s_109_41, s_109_42, s_109_43, s_109_44, s_109_45;
wire s_109_46, s_109_47, s_109_48, s_109_49, s_109_50, s_109_51;
wire s_109_52, s_109_53, s_109_54,  s_110_0,  s_110_1,  s_110_2;
wire  s_110_3,  s_110_4,  s_110_5,  s_110_6,  s_110_7,  s_110_8;
wire  s_110_9, s_110_10, s_110_11, s_110_12, s_110_13, s_110_14;
wire s_110_15, s_110_16, s_110_17, s_110_18, s_110_19, s_110_20;
wire s_110_21, s_110_22, s_110_23, s_110_24, s_110_25, s_110_26;
wire s_110_27, s_110_28, s_110_29, s_110_30, s_110_31, s_110_32;
wire s_110_33, s_110_34, s_110_35, s_110_36, s_110_37, s_110_38;
wire s_110_39, s_110_40, s_110_41, s_110_42, s_110_43, s_110_44;
wire s_110_45, s_110_46, s_110_47, s_110_48, s_110_49, s_110_50;
wire s_110_51, s_110_52, s_110_53, s_110_54, s_110_55, s_110_56;
wire  s_111_0,  s_111_1,  s_111_2,  s_111_3,  s_111_4,  s_111_5;
wire  s_111_6,  s_111_7,  s_111_8,  s_111_9, s_111_10, s_111_11;
wire s_111_12, s_111_13, s_111_14, s_111_15, s_111_16, s_111_17;
wire s_111_18, s_111_19, s_111_20, s_111_21, s_111_22, s_111_23;
wire s_111_24, s_111_25, s_111_26, s_111_27, s_111_28, s_111_29;
wire s_111_30, s_111_31, s_111_32, s_111_33, s_111_34, s_111_35;
wire s_111_36, s_111_37, s_111_38, s_111_39, s_111_40, s_111_41;
wire s_111_42, s_111_43, s_111_44, s_111_45, s_111_46, s_111_47;
wire s_111_48, s_111_49, s_111_50, s_111_51, s_111_52, s_111_53;
wire s_111_54, s_111_55,  s_112_0,  s_112_1,  s_112_2,  s_112_3;
wire  s_112_4,  s_112_5,  s_112_6,  s_112_7,  s_112_8,  s_112_9;
wire s_112_10, s_112_11, s_112_12, s_112_13, s_112_14, s_112_15;
wire s_112_16, s_112_17, s_112_18, s_112_19, s_112_20, s_112_21;
wire s_112_22, s_112_23, s_112_24, s_112_25, s_112_26, s_112_27;
wire s_112_28, s_112_29, s_112_30, s_112_31, s_112_32, s_112_33;
wire s_112_34, s_112_35, s_112_36, s_112_37, s_112_38, s_112_39;
wire s_112_40, s_112_41, s_112_42, s_112_43, s_112_44, s_112_45;
wire s_112_46, s_112_47, s_112_48, s_112_49, s_112_50, s_112_51;
wire s_112_52, s_112_53, s_112_54, s_112_55, s_112_56, s_112_57;
wire  s_113_0,  s_113_1,  s_113_2,  s_113_3,  s_113_4,  s_113_5;
wire  s_113_6,  s_113_7,  s_113_8,  s_113_9, s_113_10, s_113_11;
wire s_113_12, s_113_13, s_113_14, s_113_15, s_113_16, s_113_17;
wire s_113_18, s_113_19, s_113_20, s_113_21, s_113_22, s_113_23;
wire s_113_24, s_113_25, s_113_26, s_113_27, s_113_28, s_113_29;
wire s_113_30, s_113_31, s_113_32, s_113_33, s_113_34, s_113_35;
wire s_113_36, s_113_37, s_113_38, s_113_39, s_113_40, s_113_41;
wire s_113_42, s_113_43, s_113_44, s_113_45, s_113_46, s_113_47;
wire s_113_48, s_113_49, s_113_50, s_113_51, s_113_52, s_113_53;
wire s_113_54, s_113_55, s_113_56,  s_114_0,  s_114_1,  s_114_2;
wire  s_114_3,  s_114_4,  s_114_5,  s_114_6,  s_114_7,  s_114_8;
wire  s_114_9, s_114_10, s_114_11, s_114_12, s_114_13, s_114_14;
wire s_114_15, s_114_16, s_114_17, s_114_18, s_114_19, s_114_20;
wire s_114_21, s_114_22, s_114_23, s_114_24, s_114_25, s_114_26;
wire s_114_27, s_114_28, s_114_29, s_114_30, s_114_31, s_114_32;
wire s_114_33, s_114_34, s_114_35, s_114_36, s_114_37, s_114_38;
wire s_114_39, s_114_40, s_114_41, s_114_42, s_114_43, s_114_44;
wire s_114_45, s_114_46, s_114_47, s_114_48, s_114_49, s_114_50;
wire s_114_51, s_114_52, s_114_53, s_114_54, s_114_55, s_114_56;
wire s_114_57, s_114_58,  s_115_0,  s_115_1,  s_115_2,  s_115_3;
wire  s_115_4,  s_115_5,  s_115_6,  s_115_7,  s_115_8,  s_115_9;
wire s_115_10, s_115_11, s_115_12, s_115_13, s_115_14, s_115_15;
wire s_115_16, s_115_17, s_115_18, s_115_19, s_115_20, s_115_21;
wire s_115_22, s_115_23, s_115_24, s_115_25, s_115_26, s_115_27;
wire s_115_28, s_115_29, s_115_30, s_115_31, s_115_32, s_115_33;
wire s_115_34, s_115_35, s_115_36, s_115_37, s_115_38, s_115_39;
wire s_115_40, s_115_41, s_115_42, s_115_43, s_115_44, s_115_45;
wire s_115_46, s_115_47, s_115_48, s_115_49, s_115_50, s_115_51;
wire s_115_52, s_115_53, s_115_54, s_115_55, s_115_56, s_115_57;
wire  s_116_0,  s_116_1,  s_116_2,  s_116_3,  s_116_4,  s_116_5;
wire  s_116_6,  s_116_7,  s_116_8,  s_116_9, s_116_10, s_116_11;
wire s_116_12, s_116_13, s_116_14, s_116_15, s_116_16, s_116_17;
wire s_116_18, s_116_19, s_116_20, s_116_21, s_116_22, s_116_23;
wire s_116_24, s_116_25, s_116_26, s_116_27, s_116_28, s_116_29;
wire s_116_30, s_116_31, s_116_32, s_116_33, s_116_34, s_116_35;
wire s_116_36, s_116_37, s_116_38, s_116_39, s_116_40, s_116_41;
wire s_116_42, s_116_43, s_116_44, s_116_45, s_116_46, s_116_47;
wire s_116_48, s_116_49, s_116_50, s_116_51, s_116_52, s_116_53;
wire s_116_54, s_116_55, s_116_56, s_116_57, s_116_58, s_116_59;
wire  s_117_0,  s_117_1,  s_117_2,  s_117_3,  s_117_4,  s_117_5;
wire  s_117_6,  s_117_7,  s_117_8,  s_117_9, s_117_10, s_117_11;
wire s_117_12, s_117_13, s_117_14, s_117_15, s_117_16, s_117_17;
wire s_117_18, s_117_19, s_117_20, s_117_21, s_117_22, s_117_23;
wire s_117_24, s_117_25, s_117_26, s_117_27, s_117_28, s_117_29;
wire s_117_30, s_117_31, s_117_32, s_117_33, s_117_34, s_117_35;
wire s_117_36, s_117_37, s_117_38, s_117_39, s_117_40, s_117_41;
wire s_117_42, s_117_43, s_117_44, s_117_45, s_117_46, s_117_47;
wire s_117_48, s_117_49, s_117_50, s_117_51, s_117_52, s_117_53;
wire s_117_54, s_117_55, s_117_56, s_117_57, s_117_58,  s_118_0;
wire  s_118_1,  s_118_2,  s_118_3,  s_118_4,  s_118_5,  s_118_6;
wire  s_118_7,  s_118_8,  s_118_9, s_118_10, s_118_11, s_118_12;
wire s_118_13, s_118_14, s_118_15, s_118_16, s_118_17, s_118_18;
wire s_118_19, s_118_20, s_118_21, s_118_22, s_118_23, s_118_24;
wire s_118_25, s_118_26, s_118_27, s_118_28, s_118_29, s_118_30;
wire s_118_31, s_118_32, s_118_33, s_118_34, s_118_35, s_118_36;
wire s_118_37, s_118_38, s_118_39, s_118_40, s_118_41, s_118_42;
wire s_118_43, s_118_44, s_118_45, s_118_46, s_118_47, s_118_48;
wire s_118_49, s_118_50, s_118_51, s_118_52, s_118_53, s_118_54;
wire s_118_55, s_118_56, s_118_57, s_118_58, s_118_59, s_118_60;
wire  s_119_0,  s_119_1,  s_119_2,  s_119_3,  s_119_4,  s_119_5;
wire  s_119_6,  s_119_7,  s_119_8,  s_119_9, s_119_10, s_119_11;
wire s_119_12, s_119_13, s_119_14, s_119_15, s_119_16, s_119_17;
wire s_119_18, s_119_19, s_119_20, s_119_21, s_119_22, s_119_23;
wire s_119_24, s_119_25, s_119_26, s_119_27, s_119_28, s_119_29;
wire s_119_30, s_119_31, s_119_32, s_119_33, s_119_34, s_119_35;
wire s_119_36, s_119_37, s_119_38, s_119_39, s_119_40, s_119_41;
wire s_119_42, s_119_43, s_119_44, s_119_45, s_119_46, s_119_47;
wire s_119_48, s_119_49, s_119_50, s_119_51, s_119_52, s_119_53;
wire s_119_54, s_119_55, s_119_56, s_119_57, s_119_58, s_119_59;
wire  s_120_0,  s_120_1,  s_120_2,  s_120_3,  s_120_4,  s_120_5;
wire  s_120_6,  s_120_7,  s_120_8,  s_120_9, s_120_10, s_120_11;
wire s_120_12, s_120_13, s_120_14, s_120_15, s_120_16, s_120_17;
wire s_120_18, s_120_19, s_120_20, s_120_21, s_120_22, s_120_23;
wire s_120_24, s_120_25, s_120_26, s_120_27, s_120_28, s_120_29;
wire s_120_30, s_120_31, s_120_32, s_120_33, s_120_34, s_120_35;
wire s_120_36, s_120_37, s_120_38, s_120_39, s_120_40, s_120_41;
wire s_120_42, s_120_43, s_120_44, s_120_45, s_120_46, s_120_47;
wire s_120_48, s_120_49, s_120_50, s_120_51, s_120_52, s_120_53;
wire s_120_54, s_120_55, s_120_56, s_120_57, s_120_58, s_120_59;
wire s_120_60, s_120_61,  s_121_0,  s_121_1,  s_121_2,  s_121_3;
wire  s_121_4,  s_121_5,  s_121_6,  s_121_7,  s_121_8,  s_121_9;
wire s_121_10, s_121_11, s_121_12, s_121_13, s_121_14, s_121_15;
wire s_121_16, s_121_17, s_121_18, s_121_19, s_121_20, s_121_21;
wire s_121_22, s_121_23, s_121_24, s_121_25, s_121_26, s_121_27;
wire s_121_28, s_121_29, s_121_30, s_121_31, s_121_32, s_121_33;
wire s_121_34, s_121_35, s_121_36, s_121_37, s_121_38, s_121_39;
wire s_121_40, s_121_41, s_121_42, s_121_43, s_121_44, s_121_45;
wire s_121_46, s_121_47, s_121_48, s_121_49, s_121_50, s_121_51;
wire s_121_52, s_121_53, s_121_54, s_121_55, s_121_56, s_121_57;
wire s_121_58, s_121_59, s_121_60,  s_122_0,  s_122_1,  s_122_2;
wire  s_122_3,  s_122_4,  s_122_5,  s_122_6,  s_122_7,  s_122_8;
wire  s_122_9, s_122_10, s_122_11, s_122_12, s_122_13, s_122_14;
wire s_122_15, s_122_16, s_122_17, s_122_18, s_122_19, s_122_20;
wire s_122_21, s_122_22, s_122_23, s_122_24, s_122_25, s_122_26;
wire s_122_27, s_122_28, s_122_29, s_122_30, s_122_31, s_122_32;
wire s_122_33, s_122_34, s_122_35, s_122_36, s_122_37, s_122_38;
wire s_122_39, s_122_40, s_122_41, s_122_42, s_122_43, s_122_44;
wire s_122_45, s_122_46, s_122_47, s_122_48, s_122_49, s_122_50;
wire s_122_51, s_122_52, s_122_53, s_122_54, s_122_55, s_122_56;
wire s_122_57, s_122_58, s_122_59, s_122_60, s_122_61, s_122_62;
wire  s_123_0,  s_123_1,  s_123_2,  s_123_3,  s_123_4,  s_123_5;
wire  s_123_6,  s_123_7,  s_123_8,  s_123_9, s_123_10, s_123_11;
wire s_123_12, s_123_13, s_123_14, s_123_15, s_123_16, s_123_17;
wire s_123_18, s_123_19, s_123_20, s_123_21, s_123_22, s_123_23;
wire s_123_24, s_123_25, s_123_26, s_123_27, s_123_28, s_123_29;
wire s_123_30, s_123_31, s_123_32, s_123_33, s_123_34, s_123_35;
wire s_123_36, s_123_37, s_123_38, s_123_39, s_123_40, s_123_41;
wire s_123_42, s_123_43, s_123_44, s_123_45, s_123_46, s_123_47;
wire s_123_48, s_123_49, s_123_50, s_123_51, s_123_52, s_123_53;
wire s_123_54, s_123_55, s_123_56, s_123_57, s_123_58, s_123_59;
wire s_123_60, s_123_61,  s_124_0,  s_124_1,  s_124_2,  s_124_3;
wire  s_124_4,  s_124_5,  s_124_6,  s_124_7,  s_124_8,  s_124_9;
wire s_124_10, s_124_11, s_124_12, s_124_13, s_124_14, s_124_15;
wire s_124_16, s_124_17, s_124_18, s_124_19, s_124_20, s_124_21;
wire s_124_22, s_124_23, s_124_24, s_124_25, s_124_26, s_124_27;
wire s_124_28, s_124_29, s_124_30, s_124_31, s_124_32, s_124_33;
wire s_124_34, s_124_35, s_124_36, s_124_37, s_124_38, s_124_39;
wire s_124_40, s_124_41, s_124_42, s_124_43, s_124_44, s_124_45;
wire s_124_46, s_124_47, s_124_48, s_124_49, s_124_50, s_124_51;
wire s_124_52, s_124_53, s_124_54, s_124_55, s_124_56, s_124_57;
wire s_124_58, s_124_59, s_124_60, s_124_61, s_124_62, s_124_63;
wire  s_125_0,  s_125_1,  s_125_2,  s_125_3,  s_125_4,  s_125_5;
wire  s_125_6,  s_125_7,  s_125_8,  s_125_9, s_125_10, s_125_11;
wire s_125_12, s_125_13, s_125_14, s_125_15, s_125_16, s_125_17;
wire s_125_18, s_125_19, s_125_20, s_125_21, s_125_22, s_125_23;
wire s_125_24, s_125_25, s_125_26, s_125_27, s_125_28, s_125_29;
wire s_125_30, s_125_31, s_125_32, s_125_33, s_125_34, s_125_35;
wire s_125_36, s_125_37, s_125_38, s_125_39, s_125_40, s_125_41;
wire s_125_42, s_125_43, s_125_44, s_125_45, s_125_46, s_125_47;
wire s_125_48, s_125_49, s_125_50, s_125_51, s_125_52, s_125_53;
wire s_125_54, s_125_55, s_125_56, s_125_57, s_125_58, s_125_59;
wire s_125_60, s_125_61, s_125_62,  s_126_0,  s_126_1,  s_126_2;
wire  s_126_3,  s_126_4,  s_126_5,  s_126_6,  s_126_7,  s_126_8;
wire  s_126_9, s_126_10, s_126_11, s_126_12, s_126_13, s_126_14;
wire s_126_15, s_126_16, s_126_17, s_126_18, s_126_19, s_126_20;
wire s_126_21, s_126_22, s_126_23, s_126_24, s_126_25, s_126_26;
wire s_126_27, s_126_28, s_126_29, s_126_30, s_126_31, s_126_32;
wire s_126_33, s_126_34, s_126_35, s_126_36, s_126_37, s_126_38;
wire s_126_39, s_126_40, s_126_41, s_126_42, s_126_43, s_126_44;
wire s_126_45, s_126_46, s_126_47, s_126_48, s_126_49, s_126_50;
wire s_126_51, s_126_52, s_126_53, s_126_54, s_126_55, s_126_56;
wire s_126_57, s_126_58, s_126_59, s_126_60, s_126_61, s_126_62;
wire s_126_63, s_126_64,  s_127_0,  s_127_1,  s_127_2,  s_127_3;
wire  s_127_4,  s_127_5,  s_127_6,  s_127_7,  s_127_8,  s_127_9;
wire s_127_10, s_127_11, s_127_12, s_127_13, s_127_14, s_127_15;
wire s_127_16, s_127_17, s_127_18, s_127_19, s_127_20, s_127_21;
wire s_127_22, s_127_23, s_127_24, s_127_25, s_127_26, s_127_27;
wire s_127_28, s_127_29, s_127_30, s_127_31, s_127_32, s_127_33;
wire s_127_34, s_127_35, s_127_36, s_127_37, s_127_38, s_127_39;
wire s_127_40, s_127_41, s_127_42, s_127_43, s_127_44, s_127_45;
wire s_127_46, s_127_47, s_127_48, s_127_49, s_127_50, s_127_51;
wire s_127_52, s_127_53, s_127_54, s_127_55, s_127_56, s_127_57;
wire s_127_58, s_127_59, s_127_60, s_127_61, s_127_62, s_127_63;
wire  s_128_0,  s_128_1,  s_128_2,  s_128_3,  s_128_4,  s_128_5;
wire  s_128_6,  s_128_7,  s_128_8,  s_128_9, s_128_10, s_128_11;
wire s_128_12, s_128_13, s_128_14, s_128_15, s_128_16, s_128_17;
wire s_128_18, s_128_19, s_128_20, s_128_21, s_128_22, s_128_23;
wire s_128_24, s_128_25, s_128_26, s_128_27, s_128_28, s_128_29;
wire s_128_30, s_128_31, s_128_32, s_128_33, s_128_34, s_128_35;
wire s_128_36, s_128_37, s_128_38, s_128_39, s_128_40, s_128_41;
wire s_128_42, s_128_43, s_128_44, s_128_45, s_128_46, s_128_47;
wire s_128_48, s_128_49, s_128_50, s_128_51, s_128_52, s_128_53;
wire s_128_54, s_128_55, s_128_56, s_128_57, s_128_58, s_128_59;
wire s_128_60, s_128_61, s_128_62, s_128_63, s_128_64,  s_129_0;
wire  s_129_1,  s_129_2,  s_129_3,  s_129_4,  s_129_5,  s_129_6;
wire  s_129_7,  s_129_8,  s_129_9, s_129_10, s_129_11, s_129_12;
wire s_129_13, s_129_14, s_129_15, s_129_16, s_129_17, s_129_18;
wire s_129_19, s_129_20, s_129_21, s_129_22, s_129_23, s_129_24;
wire s_129_25, s_129_26, s_129_27, s_129_28, s_129_29, s_129_30;
wire s_129_31, s_129_32, s_129_33, s_129_34, s_129_35, s_129_36;
wire s_129_37, s_129_38, s_129_39, s_129_40, s_129_41, s_129_42;
wire s_129_43, s_129_44, s_129_45, s_129_46, s_129_47, s_129_48;
wire s_129_49, s_129_50, s_129_51, s_129_52, s_129_53, s_129_54;
wire s_129_55, s_129_56, s_129_57, s_129_58, s_129_59, s_129_60;
wire s_129_61, s_129_62, s_129_63, s_129_64,  s_130_0,  s_130_1;
wire  s_130_2,  s_130_3,  s_130_4,  s_130_5,  s_130_6,  s_130_7;
wire  s_130_8,  s_130_9, s_130_10, s_130_11, s_130_12, s_130_13;
wire s_130_14, s_130_15, s_130_16, s_130_17, s_130_18, s_130_19;
wire s_130_20, s_130_21, s_130_22, s_130_23, s_130_24, s_130_25;
wire s_130_26, s_130_27, s_130_28, s_130_29, s_130_30, s_130_31;
wire s_130_32, s_130_33, s_130_34, s_130_35, s_130_36, s_130_37;
wire s_130_38, s_130_39, s_130_40, s_130_41, s_130_42, s_130_43;
wire s_130_44, s_130_45, s_130_46, s_130_47, s_130_48, s_130_49;
wire s_130_50, s_130_51, s_130_52, s_130_53, s_130_54, s_130_55;
wire s_130_56, s_130_57, s_130_58, s_130_59, s_130_60, s_130_61;
wire s_130_62, s_130_63,  s_131_0,  s_131_1,  s_131_2,  s_131_3;
wire  s_131_4,  s_131_5,  s_131_6,  s_131_7,  s_131_8,  s_131_9;
wire s_131_10, s_131_11, s_131_12, s_131_13, s_131_14, s_131_15;
wire s_131_16, s_131_17, s_131_18, s_131_19, s_131_20, s_131_21;
wire s_131_22, s_131_23, s_131_24, s_131_25, s_131_26, s_131_27;
wire s_131_28, s_131_29, s_131_30, s_131_31, s_131_32, s_131_33;
wire s_131_34, s_131_35, s_131_36, s_131_37, s_131_38, s_131_39;
wire s_131_40, s_131_41, s_131_42, s_131_43, s_131_44, s_131_45;
wire s_131_46, s_131_47, s_131_48, s_131_49, s_131_50, s_131_51;
wire s_131_52, s_131_53, s_131_54, s_131_55, s_131_56, s_131_57;
wire s_131_58, s_131_59, s_131_60, s_131_61, s_131_62, s_131_63;
wire  s_132_0,  s_132_1,  s_132_2,  s_132_3,  s_132_4,  s_132_5;
wire  s_132_6,  s_132_7,  s_132_8,  s_132_9, s_132_10, s_132_11;
wire s_132_12, s_132_13, s_132_14, s_132_15, s_132_16, s_132_17;
wire s_132_18, s_132_19, s_132_20, s_132_21, s_132_22, s_132_23;
wire s_132_24, s_132_25, s_132_26, s_132_27, s_132_28, s_132_29;
wire s_132_30, s_132_31, s_132_32, s_132_33, s_132_34, s_132_35;
wire s_132_36, s_132_37, s_132_38, s_132_39, s_132_40, s_132_41;
wire s_132_42, s_132_43, s_132_44, s_132_45, s_132_46, s_132_47;
wire s_132_48, s_132_49, s_132_50, s_132_51, s_132_52, s_132_53;
wire s_132_54, s_132_55, s_132_56, s_132_57, s_132_58, s_132_59;
wire s_132_60, s_132_61, s_132_62,  s_133_0,  s_133_1,  s_133_2;
wire  s_133_3,  s_133_4,  s_133_5,  s_133_6,  s_133_7,  s_133_8;
wire  s_133_9, s_133_10, s_133_11, s_133_12, s_133_13, s_133_14;
wire s_133_15, s_133_16, s_133_17, s_133_18, s_133_19, s_133_20;
wire s_133_21, s_133_22, s_133_23, s_133_24, s_133_25, s_133_26;
wire s_133_27, s_133_28, s_133_29, s_133_30, s_133_31, s_133_32;
wire s_133_33, s_133_34, s_133_35, s_133_36, s_133_37, s_133_38;
wire s_133_39, s_133_40, s_133_41, s_133_42, s_133_43, s_133_44;
wire s_133_45, s_133_46, s_133_47, s_133_48, s_133_49, s_133_50;
wire s_133_51, s_133_52, s_133_53, s_133_54, s_133_55, s_133_56;
wire s_133_57, s_133_58, s_133_59, s_133_60, s_133_61, s_133_62;
wire  s_134_0,  s_134_1,  s_134_2,  s_134_3,  s_134_4,  s_134_5;
wire  s_134_6,  s_134_7,  s_134_8,  s_134_9, s_134_10, s_134_11;
wire s_134_12, s_134_13, s_134_14, s_134_15, s_134_16, s_134_17;
wire s_134_18, s_134_19, s_134_20, s_134_21, s_134_22, s_134_23;
wire s_134_24, s_134_25, s_134_26, s_134_27, s_134_28, s_134_29;
wire s_134_30, s_134_31, s_134_32, s_134_33, s_134_34, s_134_35;
wire s_134_36, s_134_37, s_134_38, s_134_39, s_134_40, s_134_41;
wire s_134_42, s_134_43, s_134_44, s_134_45, s_134_46, s_134_47;
wire s_134_48, s_134_49, s_134_50, s_134_51, s_134_52, s_134_53;
wire s_134_54, s_134_55, s_134_56, s_134_57, s_134_58, s_134_59;
wire s_134_60, s_134_61,  s_135_0,  s_135_1,  s_135_2,  s_135_3;
wire  s_135_4,  s_135_5,  s_135_6,  s_135_7,  s_135_8,  s_135_9;
wire s_135_10, s_135_11, s_135_12, s_135_13, s_135_14, s_135_15;
wire s_135_16, s_135_17, s_135_18, s_135_19, s_135_20, s_135_21;
wire s_135_22, s_135_23, s_135_24, s_135_25, s_135_26, s_135_27;
wire s_135_28, s_135_29, s_135_30, s_135_31, s_135_32, s_135_33;
wire s_135_34, s_135_35, s_135_36, s_135_37, s_135_38, s_135_39;
wire s_135_40, s_135_41, s_135_42, s_135_43, s_135_44, s_135_45;
wire s_135_46, s_135_47, s_135_48, s_135_49, s_135_50, s_135_51;
wire s_135_52, s_135_53, s_135_54, s_135_55, s_135_56, s_135_57;
wire s_135_58, s_135_59, s_135_60, s_135_61,  s_136_0,  s_136_1;
wire  s_136_2,  s_136_3,  s_136_4,  s_136_5,  s_136_6,  s_136_7;
wire  s_136_8,  s_136_9, s_136_10, s_136_11, s_136_12, s_136_13;
wire s_136_14, s_136_15, s_136_16, s_136_17, s_136_18, s_136_19;
wire s_136_20, s_136_21, s_136_22, s_136_23, s_136_24, s_136_25;
wire s_136_26, s_136_27, s_136_28, s_136_29, s_136_30, s_136_31;
wire s_136_32, s_136_33, s_136_34, s_136_35, s_136_36, s_136_37;
wire s_136_38, s_136_39, s_136_40, s_136_41, s_136_42, s_136_43;
wire s_136_44, s_136_45, s_136_46, s_136_47, s_136_48, s_136_49;
wire s_136_50, s_136_51, s_136_52, s_136_53, s_136_54, s_136_55;
wire s_136_56, s_136_57, s_136_58, s_136_59, s_136_60,  s_137_0;
wire  s_137_1,  s_137_2,  s_137_3,  s_137_4,  s_137_5,  s_137_6;
wire  s_137_7,  s_137_8,  s_137_9, s_137_10, s_137_11, s_137_12;
wire s_137_13, s_137_14, s_137_15, s_137_16, s_137_17, s_137_18;
wire s_137_19, s_137_20, s_137_21, s_137_22, s_137_23, s_137_24;
wire s_137_25, s_137_26, s_137_27, s_137_28, s_137_29, s_137_30;
wire s_137_31, s_137_32, s_137_33, s_137_34, s_137_35, s_137_36;
wire s_137_37, s_137_38, s_137_39, s_137_40, s_137_41, s_137_42;
wire s_137_43, s_137_44, s_137_45, s_137_46, s_137_47, s_137_48;
wire s_137_49, s_137_50, s_137_51, s_137_52, s_137_53, s_137_54;
wire s_137_55, s_137_56, s_137_57, s_137_58, s_137_59, s_137_60;
wire  s_138_0,  s_138_1,  s_138_2,  s_138_3,  s_138_4,  s_138_5;
wire  s_138_6,  s_138_7,  s_138_8,  s_138_9, s_138_10, s_138_11;
wire s_138_12, s_138_13, s_138_14, s_138_15, s_138_16, s_138_17;
wire s_138_18, s_138_19, s_138_20, s_138_21, s_138_22, s_138_23;
wire s_138_24, s_138_25, s_138_26, s_138_27, s_138_28, s_138_29;
wire s_138_30, s_138_31, s_138_32, s_138_33, s_138_34, s_138_35;
wire s_138_36, s_138_37, s_138_38, s_138_39, s_138_40, s_138_41;
wire s_138_42, s_138_43, s_138_44, s_138_45, s_138_46, s_138_47;
wire s_138_48, s_138_49, s_138_50, s_138_51, s_138_52, s_138_53;
wire s_138_54, s_138_55, s_138_56, s_138_57, s_138_58, s_138_59;
wire  s_139_0,  s_139_1,  s_139_2,  s_139_3,  s_139_4,  s_139_5;
wire  s_139_6,  s_139_7,  s_139_8,  s_139_9, s_139_10, s_139_11;
wire s_139_12, s_139_13, s_139_14, s_139_15, s_139_16, s_139_17;
wire s_139_18, s_139_19, s_139_20, s_139_21, s_139_22, s_139_23;
wire s_139_24, s_139_25, s_139_26, s_139_27, s_139_28, s_139_29;
wire s_139_30, s_139_31, s_139_32, s_139_33, s_139_34, s_139_35;
wire s_139_36, s_139_37, s_139_38, s_139_39, s_139_40, s_139_41;
wire s_139_42, s_139_43, s_139_44, s_139_45, s_139_46, s_139_47;
wire s_139_48, s_139_49, s_139_50, s_139_51, s_139_52, s_139_53;
wire s_139_54, s_139_55, s_139_56, s_139_57, s_139_58, s_139_59;
wire  s_140_0,  s_140_1,  s_140_2,  s_140_3,  s_140_4,  s_140_5;
wire  s_140_6,  s_140_7,  s_140_8,  s_140_9, s_140_10, s_140_11;
wire s_140_12, s_140_13, s_140_14, s_140_15, s_140_16, s_140_17;
wire s_140_18, s_140_19, s_140_20, s_140_21, s_140_22, s_140_23;
wire s_140_24, s_140_25, s_140_26, s_140_27, s_140_28, s_140_29;
wire s_140_30, s_140_31, s_140_32, s_140_33, s_140_34, s_140_35;
wire s_140_36, s_140_37, s_140_38, s_140_39, s_140_40, s_140_41;
wire s_140_42, s_140_43, s_140_44, s_140_45, s_140_46, s_140_47;
wire s_140_48, s_140_49, s_140_50, s_140_51, s_140_52, s_140_53;
wire s_140_54, s_140_55, s_140_56, s_140_57, s_140_58,  s_141_0;
wire  s_141_1,  s_141_2,  s_141_3,  s_141_4,  s_141_5,  s_141_6;
wire  s_141_7,  s_141_8,  s_141_9, s_141_10, s_141_11, s_141_12;
wire s_141_13, s_141_14, s_141_15, s_141_16, s_141_17, s_141_18;
wire s_141_19, s_141_20, s_141_21, s_141_22, s_141_23, s_141_24;
wire s_141_25, s_141_26, s_141_27, s_141_28, s_141_29, s_141_30;
wire s_141_31, s_141_32, s_141_33, s_141_34, s_141_35, s_141_36;
wire s_141_37, s_141_38, s_141_39, s_141_40, s_141_41, s_141_42;
wire s_141_43, s_141_44, s_141_45, s_141_46, s_141_47, s_141_48;
wire s_141_49, s_141_50, s_141_51, s_141_52, s_141_53, s_141_54;
wire s_141_55, s_141_56, s_141_57, s_141_58,  s_142_0,  s_142_1;
wire  s_142_2,  s_142_3,  s_142_4,  s_142_5,  s_142_6,  s_142_7;
wire  s_142_8,  s_142_9, s_142_10, s_142_11, s_142_12, s_142_13;
wire s_142_14, s_142_15, s_142_16, s_142_17, s_142_18, s_142_19;
wire s_142_20, s_142_21, s_142_22, s_142_23, s_142_24, s_142_25;
wire s_142_26, s_142_27, s_142_28, s_142_29, s_142_30, s_142_31;
wire s_142_32, s_142_33, s_142_34, s_142_35, s_142_36, s_142_37;
wire s_142_38, s_142_39, s_142_40, s_142_41, s_142_42, s_142_43;
wire s_142_44, s_142_45, s_142_46, s_142_47, s_142_48, s_142_49;
wire s_142_50, s_142_51, s_142_52, s_142_53, s_142_54, s_142_55;
wire s_142_56, s_142_57,  s_143_0,  s_143_1,  s_143_2,  s_143_3;
wire  s_143_4,  s_143_5,  s_143_6,  s_143_7,  s_143_8,  s_143_9;
wire s_143_10, s_143_11, s_143_12, s_143_13, s_143_14, s_143_15;
wire s_143_16, s_143_17, s_143_18, s_143_19, s_143_20, s_143_21;
wire s_143_22, s_143_23, s_143_24, s_143_25, s_143_26, s_143_27;
wire s_143_28, s_143_29, s_143_30, s_143_31, s_143_32, s_143_33;
wire s_143_34, s_143_35, s_143_36, s_143_37, s_143_38, s_143_39;
wire s_143_40, s_143_41, s_143_42, s_143_43, s_143_44, s_143_45;
wire s_143_46, s_143_47, s_143_48, s_143_49, s_143_50, s_143_51;
wire s_143_52, s_143_53, s_143_54, s_143_55, s_143_56, s_143_57;
wire  s_144_0,  s_144_1,  s_144_2,  s_144_3,  s_144_4,  s_144_5;
wire  s_144_6,  s_144_7,  s_144_8,  s_144_9, s_144_10, s_144_11;
wire s_144_12, s_144_13, s_144_14, s_144_15, s_144_16, s_144_17;
wire s_144_18, s_144_19, s_144_20, s_144_21, s_144_22, s_144_23;
wire s_144_24, s_144_25, s_144_26, s_144_27, s_144_28, s_144_29;
wire s_144_30, s_144_31, s_144_32, s_144_33, s_144_34, s_144_35;
wire s_144_36, s_144_37, s_144_38, s_144_39, s_144_40, s_144_41;
wire s_144_42, s_144_43, s_144_44, s_144_45, s_144_46, s_144_47;
wire s_144_48, s_144_49, s_144_50, s_144_51, s_144_52, s_144_53;
wire s_144_54, s_144_55, s_144_56,  s_145_0,  s_145_1,  s_145_2;
wire  s_145_3,  s_145_4,  s_145_5,  s_145_6,  s_145_7,  s_145_8;
wire  s_145_9, s_145_10, s_145_11, s_145_12, s_145_13, s_145_14;
wire s_145_15, s_145_16, s_145_17, s_145_18, s_145_19, s_145_20;
wire s_145_21, s_145_22, s_145_23, s_145_24, s_145_25, s_145_26;
wire s_145_27, s_145_28, s_145_29, s_145_30, s_145_31, s_145_32;
wire s_145_33, s_145_34, s_145_35, s_145_36, s_145_37, s_145_38;
wire s_145_39, s_145_40, s_145_41, s_145_42, s_145_43, s_145_44;
wire s_145_45, s_145_46, s_145_47, s_145_48, s_145_49, s_145_50;
wire s_145_51, s_145_52, s_145_53, s_145_54, s_145_55, s_145_56;
wire  s_146_0,  s_146_1,  s_146_2,  s_146_3,  s_146_4,  s_146_5;
wire  s_146_6,  s_146_7,  s_146_8,  s_146_9, s_146_10, s_146_11;
wire s_146_12, s_146_13, s_146_14, s_146_15, s_146_16, s_146_17;
wire s_146_18, s_146_19, s_146_20, s_146_21, s_146_22, s_146_23;
wire s_146_24, s_146_25, s_146_26, s_146_27, s_146_28, s_146_29;
wire s_146_30, s_146_31, s_146_32, s_146_33, s_146_34, s_146_35;
wire s_146_36, s_146_37, s_146_38, s_146_39, s_146_40, s_146_41;
wire s_146_42, s_146_43, s_146_44, s_146_45, s_146_46, s_146_47;
wire s_146_48, s_146_49, s_146_50, s_146_51, s_146_52, s_146_53;
wire s_146_54, s_146_55,  s_147_0,  s_147_1,  s_147_2,  s_147_3;
wire  s_147_4,  s_147_5,  s_147_6,  s_147_7,  s_147_8,  s_147_9;
wire s_147_10, s_147_11, s_147_12, s_147_13, s_147_14, s_147_15;
wire s_147_16, s_147_17, s_147_18, s_147_19, s_147_20, s_147_21;
wire s_147_22, s_147_23, s_147_24, s_147_25, s_147_26, s_147_27;
wire s_147_28, s_147_29, s_147_30, s_147_31, s_147_32, s_147_33;
wire s_147_34, s_147_35, s_147_36, s_147_37, s_147_38, s_147_39;
wire s_147_40, s_147_41, s_147_42, s_147_43, s_147_44, s_147_45;
wire s_147_46, s_147_47, s_147_48, s_147_49, s_147_50, s_147_51;
wire s_147_52, s_147_53, s_147_54, s_147_55,  s_148_0,  s_148_1;
wire  s_148_2,  s_148_3,  s_148_4,  s_148_5,  s_148_6,  s_148_7;
wire  s_148_8,  s_148_9, s_148_10, s_148_11, s_148_12, s_148_13;
wire s_148_14, s_148_15, s_148_16, s_148_17, s_148_18, s_148_19;
wire s_148_20, s_148_21, s_148_22, s_148_23, s_148_24, s_148_25;
wire s_148_26, s_148_27, s_148_28, s_148_29, s_148_30, s_148_31;
wire s_148_32, s_148_33, s_148_34, s_148_35, s_148_36, s_148_37;
wire s_148_38, s_148_39, s_148_40, s_148_41, s_148_42, s_148_43;
wire s_148_44, s_148_45, s_148_46, s_148_47, s_148_48, s_148_49;
wire s_148_50, s_148_51, s_148_52, s_148_53, s_148_54,  s_149_0;
wire  s_149_1,  s_149_2,  s_149_3,  s_149_4,  s_149_5,  s_149_6;
wire  s_149_7,  s_149_8,  s_149_9, s_149_10, s_149_11, s_149_12;
wire s_149_13, s_149_14, s_149_15, s_149_16, s_149_17, s_149_18;
wire s_149_19, s_149_20, s_149_21, s_149_22, s_149_23, s_149_24;
wire s_149_25, s_149_26, s_149_27, s_149_28, s_149_29, s_149_30;
wire s_149_31, s_149_32, s_149_33, s_149_34, s_149_35, s_149_36;
wire s_149_37, s_149_38, s_149_39, s_149_40, s_149_41, s_149_42;
wire s_149_43, s_149_44, s_149_45, s_149_46, s_149_47, s_149_48;
wire s_149_49, s_149_50, s_149_51, s_149_52, s_149_53, s_149_54;
wire  s_150_0,  s_150_1,  s_150_2,  s_150_3,  s_150_4,  s_150_5;
wire  s_150_6,  s_150_7,  s_150_8,  s_150_9, s_150_10, s_150_11;
wire s_150_12, s_150_13, s_150_14, s_150_15, s_150_16, s_150_17;
wire s_150_18, s_150_19, s_150_20, s_150_21, s_150_22, s_150_23;
wire s_150_24, s_150_25, s_150_26, s_150_27, s_150_28, s_150_29;
wire s_150_30, s_150_31, s_150_32, s_150_33, s_150_34, s_150_35;
wire s_150_36, s_150_37, s_150_38, s_150_39, s_150_40, s_150_41;
wire s_150_42, s_150_43, s_150_44, s_150_45, s_150_46, s_150_47;
wire s_150_48, s_150_49, s_150_50, s_150_51, s_150_52, s_150_53;
wire  s_151_0,  s_151_1,  s_151_2,  s_151_3,  s_151_4,  s_151_5;
wire  s_151_6,  s_151_7,  s_151_8,  s_151_9, s_151_10, s_151_11;
wire s_151_12, s_151_13, s_151_14, s_151_15, s_151_16, s_151_17;
wire s_151_18, s_151_19, s_151_20, s_151_21, s_151_22, s_151_23;
wire s_151_24, s_151_25, s_151_26, s_151_27, s_151_28, s_151_29;
wire s_151_30, s_151_31, s_151_32, s_151_33, s_151_34, s_151_35;
wire s_151_36, s_151_37, s_151_38, s_151_39, s_151_40, s_151_41;
wire s_151_42, s_151_43, s_151_44, s_151_45, s_151_46, s_151_47;
wire s_151_48, s_151_49, s_151_50, s_151_51, s_151_52, s_151_53;
wire  s_152_0,  s_152_1,  s_152_2,  s_152_3,  s_152_4,  s_152_5;
wire  s_152_6,  s_152_7,  s_152_8,  s_152_9, s_152_10, s_152_11;
wire s_152_12, s_152_13, s_152_14, s_152_15, s_152_16, s_152_17;
wire s_152_18, s_152_19, s_152_20, s_152_21, s_152_22, s_152_23;
wire s_152_24, s_152_25, s_152_26, s_152_27, s_152_28, s_152_29;
wire s_152_30, s_152_31, s_152_32, s_152_33, s_152_34, s_152_35;
wire s_152_36, s_152_37, s_152_38, s_152_39, s_152_40, s_152_41;
wire s_152_42, s_152_43, s_152_44, s_152_45, s_152_46, s_152_47;
wire s_152_48, s_152_49, s_152_50, s_152_51, s_152_52,  s_153_0;
wire  s_153_1,  s_153_2,  s_153_3,  s_153_4,  s_153_5,  s_153_6;
wire  s_153_7,  s_153_8,  s_153_9, s_153_10, s_153_11, s_153_12;
wire s_153_13, s_153_14, s_153_15, s_153_16, s_153_17, s_153_18;
wire s_153_19, s_153_20, s_153_21, s_153_22, s_153_23, s_153_24;
wire s_153_25, s_153_26, s_153_27, s_153_28, s_153_29, s_153_30;
wire s_153_31, s_153_32, s_153_33, s_153_34, s_153_35, s_153_36;
wire s_153_37, s_153_38, s_153_39, s_153_40, s_153_41, s_153_42;
wire s_153_43, s_153_44, s_153_45, s_153_46, s_153_47, s_153_48;
wire s_153_49, s_153_50, s_153_51, s_153_52,  s_154_0,  s_154_1;
wire  s_154_2,  s_154_3,  s_154_4,  s_154_5,  s_154_6,  s_154_7;
wire  s_154_8,  s_154_9, s_154_10, s_154_11, s_154_12, s_154_13;
wire s_154_14, s_154_15, s_154_16, s_154_17, s_154_18, s_154_19;
wire s_154_20, s_154_21, s_154_22, s_154_23, s_154_24, s_154_25;
wire s_154_26, s_154_27, s_154_28, s_154_29, s_154_30, s_154_31;
wire s_154_32, s_154_33, s_154_34, s_154_35, s_154_36, s_154_37;
wire s_154_38, s_154_39, s_154_40, s_154_41, s_154_42, s_154_43;
wire s_154_44, s_154_45, s_154_46, s_154_47, s_154_48, s_154_49;
wire s_154_50, s_154_51,  s_155_0,  s_155_1,  s_155_2,  s_155_3;
wire  s_155_4,  s_155_5,  s_155_6,  s_155_7,  s_155_8,  s_155_9;
wire s_155_10, s_155_11, s_155_12, s_155_13, s_155_14, s_155_15;
wire s_155_16, s_155_17, s_155_18, s_155_19, s_155_20, s_155_21;
wire s_155_22, s_155_23, s_155_24, s_155_25, s_155_26, s_155_27;
wire s_155_28, s_155_29, s_155_30, s_155_31, s_155_32, s_155_33;
wire s_155_34, s_155_35, s_155_36, s_155_37, s_155_38, s_155_39;
wire s_155_40, s_155_41, s_155_42, s_155_43, s_155_44, s_155_45;
wire s_155_46, s_155_47, s_155_48, s_155_49, s_155_50, s_155_51;
wire  s_156_0,  s_156_1,  s_156_2,  s_156_3,  s_156_4,  s_156_5;
wire  s_156_6,  s_156_7,  s_156_8,  s_156_9, s_156_10, s_156_11;
wire s_156_12, s_156_13, s_156_14, s_156_15, s_156_16, s_156_17;
wire s_156_18, s_156_19, s_156_20, s_156_21, s_156_22, s_156_23;
wire s_156_24, s_156_25, s_156_26, s_156_27, s_156_28, s_156_29;
wire s_156_30, s_156_31, s_156_32, s_156_33, s_156_34, s_156_35;
wire s_156_36, s_156_37, s_156_38, s_156_39, s_156_40, s_156_41;
wire s_156_42, s_156_43, s_156_44, s_156_45, s_156_46, s_156_47;
wire s_156_48, s_156_49, s_156_50,  s_157_0,  s_157_1,  s_157_2;
wire  s_157_3,  s_157_4,  s_157_5,  s_157_6,  s_157_7,  s_157_8;
wire  s_157_9, s_157_10, s_157_11, s_157_12, s_157_13, s_157_14;
wire s_157_15, s_157_16, s_157_17, s_157_18, s_157_19, s_157_20;
wire s_157_21, s_157_22, s_157_23, s_157_24, s_157_25, s_157_26;
wire s_157_27, s_157_28, s_157_29, s_157_30, s_157_31, s_157_32;
wire s_157_33, s_157_34, s_157_35, s_157_36, s_157_37, s_157_38;
wire s_157_39, s_157_40, s_157_41, s_157_42, s_157_43, s_157_44;
wire s_157_45, s_157_46, s_157_47, s_157_48, s_157_49, s_157_50;
wire  s_158_0,  s_158_1,  s_158_2,  s_158_3,  s_158_4,  s_158_5;
wire  s_158_6,  s_158_7,  s_158_8,  s_158_9, s_158_10, s_158_11;
wire s_158_12, s_158_13, s_158_14, s_158_15, s_158_16, s_158_17;
wire s_158_18, s_158_19, s_158_20, s_158_21, s_158_22, s_158_23;
wire s_158_24, s_158_25, s_158_26, s_158_27, s_158_28, s_158_29;
wire s_158_30, s_158_31, s_158_32, s_158_33, s_158_34, s_158_35;
wire s_158_36, s_158_37, s_158_38, s_158_39, s_158_40, s_158_41;
wire s_158_42, s_158_43, s_158_44, s_158_45, s_158_46, s_158_47;
wire s_158_48, s_158_49,  s_159_0,  s_159_1,  s_159_2,  s_159_3;
wire  s_159_4,  s_159_5,  s_159_6,  s_159_7,  s_159_8,  s_159_9;
wire s_159_10, s_159_11, s_159_12, s_159_13, s_159_14, s_159_15;
wire s_159_16, s_159_17, s_159_18, s_159_19, s_159_20, s_159_21;
wire s_159_22, s_159_23, s_159_24, s_159_25, s_159_26, s_159_27;
wire s_159_28, s_159_29, s_159_30, s_159_31, s_159_32, s_159_33;
wire s_159_34, s_159_35, s_159_36, s_159_37, s_159_38, s_159_39;
wire s_159_40, s_159_41, s_159_42, s_159_43, s_159_44, s_159_45;
wire s_159_46, s_159_47, s_159_48, s_159_49,  s_160_0,  s_160_1;
wire  s_160_2,  s_160_3,  s_160_4,  s_160_5,  s_160_6,  s_160_7;
wire  s_160_8,  s_160_9, s_160_10, s_160_11, s_160_12, s_160_13;
wire s_160_14, s_160_15, s_160_16, s_160_17, s_160_18, s_160_19;
wire s_160_20, s_160_21, s_160_22, s_160_23, s_160_24, s_160_25;
wire s_160_26, s_160_27, s_160_28, s_160_29, s_160_30, s_160_31;
wire s_160_32, s_160_33, s_160_34, s_160_35, s_160_36, s_160_37;
wire s_160_38, s_160_39, s_160_40, s_160_41, s_160_42, s_160_43;
wire s_160_44, s_160_45, s_160_46, s_160_47, s_160_48,  s_161_0;
wire  s_161_1,  s_161_2,  s_161_3,  s_161_4,  s_161_5,  s_161_6;
wire  s_161_7,  s_161_8,  s_161_9, s_161_10, s_161_11, s_161_12;
wire s_161_13, s_161_14, s_161_15, s_161_16, s_161_17, s_161_18;
wire s_161_19, s_161_20, s_161_21, s_161_22, s_161_23, s_161_24;
wire s_161_25, s_161_26, s_161_27, s_161_28, s_161_29, s_161_30;
wire s_161_31, s_161_32, s_161_33, s_161_34, s_161_35, s_161_36;
wire s_161_37, s_161_38, s_161_39, s_161_40, s_161_41, s_161_42;
wire s_161_43, s_161_44, s_161_45, s_161_46, s_161_47, s_161_48;
wire  s_162_0,  s_162_1,  s_162_2,  s_162_3,  s_162_4,  s_162_5;
wire  s_162_6,  s_162_7,  s_162_8,  s_162_9, s_162_10, s_162_11;
wire s_162_12, s_162_13, s_162_14, s_162_15, s_162_16, s_162_17;
wire s_162_18, s_162_19, s_162_20, s_162_21, s_162_22, s_162_23;
wire s_162_24, s_162_25, s_162_26, s_162_27, s_162_28, s_162_29;
wire s_162_30, s_162_31, s_162_32, s_162_33, s_162_34, s_162_35;
wire s_162_36, s_162_37, s_162_38, s_162_39, s_162_40, s_162_41;
wire s_162_42, s_162_43, s_162_44, s_162_45, s_162_46, s_162_47;
wire  s_163_0,  s_163_1,  s_163_2,  s_163_3,  s_163_4,  s_163_5;
wire  s_163_6,  s_163_7,  s_163_8,  s_163_9, s_163_10, s_163_11;
wire s_163_12, s_163_13, s_163_14, s_163_15, s_163_16, s_163_17;
wire s_163_18, s_163_19, s_163_20, s_163_21, s_163_22, s_163_23;
wire s_163_24, s_163_25, s_163_26, s_163_27, s_163_28, s_163_29;
wire s_163_30, s_163_31, s_163_32, s_163_33, s_163_34, s_163_35;
wire s_163_36, s_163_37, s_163_38, s_163_39, s_163_40, s_163_41;
wire s_163_42, s_163_43, s_163_44, s_163_45, s_163_46, s_163_47;
wire  s_164_0,  s_164_1,  s_164_2,  s_164_3,  s_164_4,  s_164_5;
wire  s_164_6,  s_164_7,  s_164_8,  s_164_9, s_164_10, s_164_11;
wire s_164_12, s_164_13, s_164_14, s_164_15, s_164_16, s_164_17;
wire s_164_18, s_164_19, s_164_20, s_164_21, s_164_22, s_164_23;
wire s_164_24, s_164_25, s_164_26, s_164_27, s_164_28, s_164_29;
wire s_164_30, s_164_31, s_164_32, s_164_33, s_164_34, s_164_35;
wire s_164_36, s_164_37, s_164_38, s_164_39, s_164_40, s_164_41;
wire s_164_42, s_164_43, s_164_44, s_164_45, s_164_46,  s_165_0;
wire  s_165_1,  s_165_2,  s_165_3,  s_165_4,  s_165_5,  s_165_6;
wire  s_165_7,  s_165_8,  s_165_9, s_165_10, s_165_11, s_165_12;
wire s_165_13, s_165_14, s_165_15, s_165_16, s_165_17, s_165_18;
wire s_165_19, s_165_20, s_165_21, s_165_22, s_165_23, s_165_24;
wire s_165_25, s_165_26, s_165_27, s_165_28, s_165_29, s_165_30;
wire s_165_31, s_165_32, s_165_33, s_165_34, s_165_35, s_165_36;
wire s_165_37, s_165_38, s_165_39, s_165_40, s_165_41, s_165_42;
wire s_165_43, s_165_44, s_165_45, s_165_46,  s_166_0,  s_166_1;
wire  s_166_2,  s_166_3,  s_166_4,  s_166_5,  s_166_6,  s_166_7;
wire  s_166_8,  s_166_9, s_166_10, s_166_11, s_166_12, s_166_13;
wire s_166_14, s_166_15, s_166_16, s_166_17, s_166_18, s_166_19;
wire s_166_20, s_166_21, s_166_22, s_166_23, s_166_24, s_166_25;
wire s_166_26, s_166_27, s_166_28, s_166_29, s_166_30, s_166_31;
wire s_166_32, s_166_33, s_166_34, s_166_35, s_166_36, s_166_37;
wire s_166_38, s_166_39, s_166_40, s_166_41, s_166_42, s_166_43;
wire s_166_44, s_166_45,  s_167_0,  s_167_1,  s_167_2,  s_167_3;
wire  s_167_4,  s_167_5,  s_167_6,  s_167_7,  s_167_8,  s_167_9;
wire s_167_10, s_167_11, s_167_12, s_167_13, s_167_14, s_167_15;
wire s_167_16, s_167_17, s_167_18, s_167_19, s_167_20, s_167_21;
wire s_167_22, s_167_23, s_167_24, s_167_25, s_167_26, s_167_27;
wire s_167_28, s_167_29, s_167_30, s_167_31, s_167_32, s_167_33;
wire s_167_34, s_167_35, s_167_36, s_167_37, s_167_38, s_167_39;
wire s_167_40, s_167_41, s_167_42, s_167_43, s_167_44, s_167_45;
wire  s_168_0,  s_168_1,  s_168_2,  s_168_3,  s_168_4,  s_168_5;
wire  s_168_6,  s_168_7,  s_168_8,  s_168_9, s_168_10, s_168_11;
wire s_168_12, s_168_13, s_168_14, s_168_15, s_168_16, s_168_17;
wire s_168_18, s_168_19, s_168_20, s_168_21, s_168_22, s_168_23;
wire s_168_24, s_168_25, s_168_26, s_168_27, s_168_28, s_168_29;
wire s_168_30, s_168_31, s_168_32, s_168_33, s_168_34, s_168_35;
wire s_168_36, s_168_37, s_168_38, s_168_39, s_168_40, s_168_41;
wire s_168_42, s_168_43, s_168_44,  s_169_0,  s_169_1,  s_169_2;
wire  s_169_3,  s_169_4,  s_169_5,  s_169_6,  s_169_7,  s_169_8;
wire  s_169_9, s_169_10, s_169_11, s_169_12, s_169_13, s_169_14;
wire s_169_15, s_169_16, s_169_17, s_169_18, s_169_19, s_169_20;
wire s_169_21, s_169_22, s_169_23, s_169_24, s_169_25, s_169_26;
wire s_169_27, s_169_28, s_169_29, s_169_30, s_169_31, s_169_32;
wire s_169_33, s_169_34, s_169_35, s_169_36, s_169_37, s_169_38;
wire s_169_39, s_169_40, s_169_41, s_169_42, s_169_43, s_169_44;
wire  s_170_0,  s_170_1,  s_170_2,  s_170_3,  s_170_4,  s_170_5;
wire  s_170_6,  s_170_7,  s_170_8,  s_170_9, s_170_10, s_170_11;
wire s_170_12, s_170_13, s_170_14, s_170_15, s_170_16, s_170_17;
wire s_170_18, s_170_19, s_170_20, s_170_21, s_170_22, s_170_23;
wire s_170_24, s_170_25, s_170_26, s_170_27, s_170_28, s_170_29;
wire s_170_30, s_170_31, s_170_32, s_170_33, s_170_34, s_170_35;
wire s_170_36, s_170_37, s_170_38, s_170_39, s_170_40, s_170_41;
wire s_170_42, s_170_43,  s_171_0,  s_171_1,  s_171_2,  s_171_3;
wire  s_171_4,  s_171_5,  s_171_6,  s_171_7,  s_171_8,  s_171_9;
wire s_171_10, s_171_11, s_171_12, s_171_13, s_171_14, s_171_15;
wire s_171_16, s_171_17, s_171_18, s_171_19, s_171_20, s_171_21;
wire s_171_22, s_171_23, s_171_24, s_171_25, s_171_26, s_171_27;
wire s_171_28, s_171_29, s_171_30, s_171_31, s_171_32, s_171_33;
wire s_171_34, s_171_35, s_171_36, s_171_37, s_171_38, s_171_39;
wire s_171_40, s_171_41, s_171_42, s_171_43,  s_172_0,  s_172_1;
wire  s_172_2,  s_172_3,  s_172_4,  s_172_5,  s_172_6,  s_172_7;
wire  s_172_8,  s_172_9, s_172_10, s_172_11, s_172_12, s_172_13;
wire s_172_14, s_172_15, s_172_16, s_172_17, s_172_18, s_172_19;
wire s_172_20, s_172_21, s_172_22, s_172_23, s_172_24, s_172_25;
wire s_172_26, s_172_27, s_172_28, s_172_29, s_172_30, s_172_31;
wire s_172_32, s_172_33, s_172_34, s_172_35, s_172_36, s_172_37;
wire s_172_38, s_172_39, s_172_40, s_172_41, s_172_42,  s_173_0;
wire  s_173_1,  s_173_2,  s_173_3,  s_173_4,  s_173_5,  s_173_6;
wire  s_173_7,  s_173_8,  s_173_9, s_173_10, s_173_11, s_173_12;
wire s_173_13, s_173_14, s_173_15, s_173_16, s_173_17, s_173_18;
wire s_173_19, s_173_20, s_173_21, s_173_22, s_173_23, s_173_24;
wire s_173_25, s_173_26, s_173_27, s_173_28, s_173_29, s_173_30;
wire s_173_31, s_173_32, s_173_33, s_173_34, s_173_35, s_173_36;
wire s_173_37, s_173_38, s_173_39, s_173_40, s_173_41, s_173_42;
wire  s_174_0,  s_174_1,  s_174_2,  s_174_3,  s_174_4,  s_174_5;
wire  s_174_6,  s_174_7,  s_174_8,  s_174_9, s_174_10, s_174_11;
wire s_174_12, s_174_13, s_174_14, s_174_15, s_174_16, s_174_17;
wire s_174_18, s_174_19, s_174_20, s_174_21, s_174_22, s_174_23;
wire s_174_24, s_174_25, s_174_26, s_174_27, s_174_28, s_174_29;
wire s_174_30, s_174_31, s_174_32, s_174_33, s_174_34, s_174_35;
wire s_174_36, s_174_37, s_174_38, s_174_39, s_174_40, s_174_41;
wire  s_175_0,  s_175_1,  s_175_2,  s_175_3,  s_175_4,  s_175_5;
wire  s_175_6,  s_175_7,  s_175_8,  s_175_9, s_175_10, s_175_11;
wire s_175_12, s_175_13, s_175_14, s_175_15, s_175_16, s_175_17;
wire s_175_18, s_175_19, s_175_20, s_175_21, s_175_22, s_175_23;
wire s_175_24, s_175_25, s_175_26, s_175_27, s_175_28, s_175_29;
wire s_175_30, s_175_31, s_175_32, s_175_33, s_175_34, s_175_35;
wire s_175_36, s_175_37, s_175_38, s_175_39, s_175_40, s_175_41;
wire  s_176_0,  s_176_1,  s_176_2,  s_176_3,  s_176_4,  s_176_5;
wire  s_176_6,  s_176_7,  s_176_8,  s_176_9, s_176_10, s_176_11;
wire s_176_12, s_176_13, s_176_14, s_176_15, s_176_16, s_176_17;
wire s_176_18, s_176_19, s_176_20, s_176_21, s_176_22, s_176_23;
wire s_176_24, s_176_25, s_176_26, s_176_27, s_176_28, s_176_29;
wire s_176_30, s_176_31, s_176_32, s_176_33, s_176_34, s_176_35;
wire s_176_36, s_176_37, s_176_38, s_176_39, s_176_40,  s_177_0;
wire  s_177_1,  s_177_2,  s_177_3,  s_177_4,  s_177_5,  s_177_6;
wire  s_177_7,  s_177_8,  s_177_9, s_177_10, s_177_11, s_177_12;
wire s_177_13, s_177_14, s_177_15, s_177_16, s_177_17, s_177_18;
wire s_177_19, s_177_20, s_177_21, s_177_22, s_177_23, s_177_24;
wire s_177_25, s_177_26, s_177_27, s_177_28, s_177_29, s_177_30;
wire s_177_31, s_177_32, s_177_33, s_177_34, s_177_35, s_177_36;
wire s_177_37, s_177_38, s_177_39, s_177_40,  s_178_0,  s_178_1;
wire  s_178_2,  s_178_3,  s_178_4,  s_178_5,  s_178_6,  s_178_7;
wire  s_178_8,  s_178_9, s_178_10, s_178_11, s_178_12, s_178_13;
wire s_178_14, s_178_15, s_178_16, s_178_17, s_178_18, s_178_19;
wire s_178_20, s_178_21, s_178_22, s_178_23, s_178_24, s_178_25;
wire s_178_26, s_178_27, s_178_28, s_178_29, s_178_30, s_178_31;
wire s_178_32, s_178_33, s_178_34, s_178_35, s_178_36, s_178_37;
wire s_178_38, s_178_39,  s_179_0,  s_179_1,  s_179_2,  s_179_3;
wire  s_179_4,  s_179_5,  s_179_6,  s_179_7,  s_179_8,  s_179_9;
wire s_179_10, s_179_11, s_179_12, s_179_13, s_179_14, s_179_15;
wire s_179_16, s_179_17, s_179_18, s_179_19, s_179_20, s_179_21;
wire s_179_22, s_179_23, s_179_24, s_179_25, s_179_26, s_179_27;
wire s_179_28, s_179_29, s_179_30, s_179_31, s_179_32, s_179_33;
wire s_179_34, s_179_35, s_179_36, s_179_37, s_179_38, s_179_39;
wire  s_180_0,  s_180_1,  s_180_2,  s_180_3,  s_180_4,  s_180_5;
wire  s_180_6,  s_180_7,  s_180_8,  s_180_9, s_180_10, s_180_11;
wire s_180_12, s_180_13, s_180_14, s_180_15, s_180_16, s_180_17;
wire s_180_18, s_180_19, s_180_20, s_180_21, s_180_22, s_180_23;
wire s_180_24, s_180_25, s_180_26, s_180_27, s_180_28, s_180_29;
wire s_180_30, s_180_31, s_180_32, s_180_33, s_180_34, s_180_35;
wire s_180_36, s_180_37, s_180_38,  s_181_0,  s_181_1,  s_181_2;
wire  s_181_3,  s_181_4,  s_181_5,  s_181_6,  s_181_7,  s_181_8;
wire  s_181_9, s_181_10, s_181_11, s_181_12, s_181_13, s_181_14;
wire s_181_15, s_181_16, s_181_17, s_181_18, s_181_19, s_181_20;
wire s_181_21, s_181_22, s_181_23, s_181_24, s_181_25, s_181_26;
wire s_181_27, s_181_28, s_181_29, s_181_30, s_181_31, s_181_32;
wire s_181_33, s_181_34, s_181_35, s_181_36, s_181_37, s_181_38;
wire  s_182_0,  s_182_1,  s_182_2,  s_182_3,  s_182_4,  s_182_5;
wire  s_182_6,  s_182_7,  s_182_8,  s_182_9, s_182_10, s_182_11;
wire s_182_12, s_182_13, s_182_14, s_182_15, s_182_16, s_182_17;
wire s_182_18, s_182_19, s_182_20, s_182_21, s_182_22, s_182_23;
wire s_182_24, s_182_25, s_182_26, s_182_27, s_182_28, s_182_29;
wire s_182_30, s_182_31, s_182_32, s_182_33, s_182_34, s_182_35;
wire s_182_36, s_182_37,  s_183_0,  s_183_1,  s_183_2,  s_183_3;
wire  s_183_4,  s_183_5,  s_183_6,  s_183_7,  s_183_8,  s_183_9;
wire s_183_10, s_183_11, s_183_12, s_183_13, s_183_14, s_183_15;
wire s_183_16, s_183_17, s_183_18, s_183_19, s_183_20, s_183_21;
wire s_183_22, s_183_23, s_183_24, s_183_25, s_183_26, s_183_27;
wire s_183_28, s_183_29, s_183_30, s_183_31, s_183_32, s_183_33;
wire s_183_34, s_183_35, s_183_36, s_183_37,  s_184_0,  s_184_1;
wire  s_184_2,  s_184_3,  s_184_4,  s_184_5,  s_184_6,  s_184_7;
wire  s_184_8,  s_184_9, s_184_10, s_184_11, s_184_12, s_184_13;
wire s_184_14, s_184_15, s_184_16, s_184_17, s_184_18, s_184_19;
wire s_184_20, s_184_21, s_184_22, s_184_23, s_184_24, s_184_25;
wire s_184_26, s_184_27, s_184_28, s_184_29, s_184_30, s_184_31;
wire s_184_32, s_184_33, s_184_34, s_184_35, s_184_36,  s_185_0;
wire  s_185_1,  s_185_2,  s_185_3,  s_185_4,  s_185_5,  s_185_6;
wire  s_185_7,  s_185_8,  s_185_9, s_185_10, s_185_11, s_185_12;
wire s_185_13, s_185_14, s_185_15, s_185_16, s_185_17, s_185_18;
wire s_185_19, s_185_20, s_185_21, s_185_22, s_185_23, s_185_24;
wire s_185_25, s_185_26, s_185_27, s_185_28, s_185_29, s_185_30;
wire s_185_31, s_185_32, s_185_33, s_185_34, s_185_35, s_185_36;
wire  s_186_0,  s_186_1,  s_186_2,  s_186_3,  s_186_4,  s_186_5;
wire  s_186_6,  s_186_7,  s_186_8,  s_186_9, s_186_10, s_186_11;
wire s_186_12, s_186_13, s_186_14, s_186_15, s_186_16, s_186_17;
wire s_186_18, s_186_19, s_186_20, s_186_21, s_186_22, s_186_23;
wire s_186_24, s_186_25, s_186_26, s_186_27, s_186_28, s_186_29;
wire s_186_30, s_186_31, s_186_32, s_186_33, s_186_34, s_186_35;
wire  s_187_0,  s_187_1,  s_187_2,  s_187_3,  s_187_4,  s_187_5;
wire  s_187_6,  s_187_7,  s_187_8,  s_187_9, s_187_10, s_187_11;
wire s_187_12, s_187_13, s_187_14, s_187_15, s_187_16, s_187_17;
wire s_187_18, s_187_19, s_187_20, s_187_21, s_187_22, s_187_23;
wire s_187_24, s_187_25, s_187_26, s_187_27, s_187_28, s_187_29;
wire s_187_30, s_187_31, s_187_32, s_187_33, s_187_34, s_187_35;
wire  s_188_0,  s_188_1,  s_188_2,  s_188_3,  s_188_4,  s_188_5;
wire  s_188_6,  s_188_7,  s_188_8,  s_188_9, s_188_10, s_188_11;
wire s_188_12, s_188_13, s_188_14, s_188_15, s_188_16, s_188_17;
wire s_188_18, s_188_19, s_188_20, s_188_21, s_188_22, s_188_23;
wire s_188_24, s_188_25, s_188_26, s_188_27, s_188_28, s_188_29;
wire s_188_30, s_188_31, s_188_32, s_188_33, s_188_34,  s_189_0;
wire  s_189_1,  s_189_2,  s_189_3,  s_189_4,  s_189_5,  s_189_6;
wire  s_189_7,  s_189_8,  s_189_9, s_189_10, s_189_11, s_189_12;
wire s_189_13, s_189_14, s_189_15, s_189_16, s_189_17, s_189_18;
wire s_189_19, s_189_20, s_189_21, s_189_22, s_189_23, s_189_24;
wire s_189_25, s_189_26, s_189_27, s_189_28, s_189_29, s_189_30;
wire s_189_31, s_189_32, s_189_33, s_189_34,  s_190_0,  s_190_1;
wire  s_190_2,  s_190_3,  s_190_4,  s_190_5,  s_190_6,  s_190_7;
wire  s_190_8,  s_190_9, s_190_10, s_190_11, s_190_12, s_190_13;
wire s_190_14, s_190_15, s_190_16, s_190_17, s_190_18, s_190_19;
wire s_190_20, s_190_21, s_190_22, s_190_23, s_190_24, s_190_25;
wire s_190_26, s_190_27, s_190_28, s_190_29, s_190_30, s_190_31;
wire s_190_32, s_190_33,  s_191_0,  s_191_1,  s_191_2,  s_191_3;
wire  s_191_4,  s_191_5,  s_191_6,  s_191_7,  s_191_8,  s_191_9;
wire s_191_10, s_191_11, s_191_12, s_191_13, s_191_14, s_191_15;
wire s_191_16, s_191_17, s_191_18, s_191_19, s_191_20, s_191_21;
wire s_191_22, s_191_23, s_191_24, s_191_25, s_191_26, s_191_27;
wire s_191_28, s_191_29, s_191_30, s_191_31, s_191_32, s_191_33;
wire  s_192_0,  s_192_1,  s_192_2,  s_192_3,  s_192_4,  s_192_5;
wire  s_192_6,  s_192_7,  s_192_8,  s_192_9, s_192_10, s_192_11;
wire s_192_12, s_192_13, s_192_14, s_192_15, s_192_16, s_192_17;
wire s_192_18, s_192_19, s_192_20, s_192_21, s_192_22, s_192_23;
wire s_192_24, s_192_25, s_192_26, s_192_27, s_192_28, s_192_29;
wire s_192_30, s_192_31, s_192_32,  s_193_0,  s_193_1,  s_193_2;
wire  s_193_3,  s_193_4,  s_193_5,  s_193_6,  s_193_7,  s_193_8;
wire  s_193_9, s_193_10, s_193_11, s_193_12, s_193_13, s_193_14;
wire s_193_15, s_193_16, s_193_17, s_193_18, s_193_19, s_193_20;
wire s_193_21, s_193_22, s_193_23, s_193_24, s_193_25, s_193_26;
wire s_193_27, s_193_28, s_193_29, s_193_30, s_193_31, s_193_32;
wire  s_194_0,  s_194_1,  s_194_2,  s_194_3,  s_194_4,  s_194_5;
wire  s_194_6,  s_194_7,  s_194_8,  s_194_9, s_194_10, s_194_11;
wire s_194_12, s_194_13, s_194_14, s_194_15, s_194_16, s_194_17;
wire s_194_18, s_194_19, s_194_20, s_194_21, s_194_22, s_194_23;
wire s_194_24, s_194_25, s_194_26, s_194_27, s_194_28, s_194_29;
wire s_194_30, s_194_31,  s_195_0,  s_195_1,  s_195_2,  s_195_3;
wire  s_195_4,  s_195_5,  s_195_6,  s_195_7,  s_195_8,  s_195_9;
wire s_195_10, s_195_11, s_195_12, s_195_13, s_195_14, s_195_15;
wire s_195_16, s_195_17, s_195_18, s_195_19, s_195_20, s_195_21;
wire s_195_22, s_195_23, s_195_24, s_195_25, s_195_26, s_195_27;
wire s_195_28, s_195_29, s_195_30, s_195_31,  s_196_0,  s_196_1;
wire  s_196_2,  s_196_3,  s_196_4,  s_196_5,  s_196_6,  s_196_7;
wire  s_196_8,  s_196_9, s_196_10, s_196_11, s_196_12, s_196_13;
wire s_196_14, s_196_15, s_196_16, s_196_17, s_196_18, s_196_19;
wire s_196_20, s_196_21, s_196_22, s_196_23, s_196_24, s_196_25;
wire s_196_26, s_196_27, s_196_28, s_196_29, s_196_30,  s_197_0;
wire  s_197_1,  s_197_2,  s_197_3,  s_197_4,  s_197_5,  s_197_6;
wire  s_197_7,  s_197_8,  s_197_9, s_197_10, s_197_11, s_197_12;
wire s_197_13, s_197_14, s_197_15, s_197_16, s_197_17, s_197_18;
wire s_197_19, s_197_20, s_197_21, s_197_22, s_197_23, s_197_24;
wire s_197_25, s_197_26, s_197_27, s_197_28, s_197_29, s_197_30;
wire  s_198_0,  s_198_1,  s_198_2,  s_198_3,  s_198_4,  s_198_5;
wire  s_198_6,  s_198_7,  s_198_8,  s_198_9, s_198_10, s_198_11;
wire s_198_12, s_198_13, s_198_14, s_198_15, s_198_16, s_198_17;
wire s_198_18, s_198_19, s_198_20, s_198_21, s_198_22, s_198_23;
wire s_198_24, s_198_25, s_198_26, s_198_27, s_198_28, s_198_29;
wire  s_199_0,  s_199_1,  s_199_2,  s_199_3,  s_199_4,  s_199_5;
wire  s_199_6,  s_199_7,  s_199_8,  s_199_9, s_199_10, s_199_11;
wire s_199_12, s_199_13, s_199_14, s_199_15, s_199_16, s_199_17;
wire s_199_18, s_199_19, s_199_20, s_199_21, s_199_22, s_199_23;
wire s_199_24, s_199_25, s_199_26, s_199_27, s_199_28, s_199_29;
wire  s_200_0,  s_200_1,  s_200_2,  s_200_3,  s_200_4,  s_200_5;
wire  s_200_6,  s_200_7,  s_200_8,  s_200_9, s_200_10, s_200_11;
wire s_200_12, s_200_13, s_200_14, s_200_15, s_200_16, s_200_17;
wire s_200_18, s_200_19, s_200_20, s_200_21, s_200_22, s_200_23;
wire s_200_24, s_200_25, s_200_26, s_200_27, s_200_28,  s_201_0;
wire  s_201_1,  s_201_2,  s_201_3,  s_201_4,  s_201_5,  s_201_6;
wire  s_201_7,  s_201_8,  s_201_9, s_201_10, s_201_11, s_201_12;
wire s_201_13, s_201_14, s_201_15, s_201_16, s_201_17, s_201_18;
wire s_201_19, s_201_20, s_201_21, s_201_22, s_201_23, s_201_24;
wire s_201_25, s_201_26, s_201_27, s_201_28,  s_202_0,  s_202_1;
wire  s_202_2,  s_202_3,  s_202_4,  s_202_5,  s_202_6,  s_202_7;
wire  s_202_8,  s_202_9, s_202_10, s_202_11, s_202_12, s_202_13;
wire s_202_14, s_202_15, s_202_16, s_202_17, s_202_18, s_202_19;
wire s_202_20, s_202_21, s_202_22, s_202_23, s_202_24, s_202_25;
wire s_202_26, s_202_27,  s_203_0,  s_203_1,  s_203_2,  s_203_3;
wire  s_203_4,  s_203_5,  s_203_6,  s_203_7,  s_203_8,  s_203_9;
wire s_203_10, s_203_11, s_203_12, s_203_13, s_203_14, s_203_15;
wire s_203_16, s_203_17, s_203_18, s_203_19, s_203_20, s_203_21;
wire s_203_22, s_203_23, s_203_24, s_203_25, s_203_26, s_203_27;
wire  s_204_0,  s_204_1,  s_204_2,  s_204_3,  s_204_4,  s_204_5;
wire  s_204_6,  s_204_7,  s_204_8,  s_204_9, s_204_10, s_204_11;
wire s_204_12, s_204_13, s_204_14, s_204_15, s_204_16, s_204_17;
wire s_204_18, s_204_19, s_204_20, s_204_21, s_204_22, s_204_23;
wire s_204_24, s_204_25, s_204_26,  s_205_0,  s_205_1,  s_205_2;
wire  s_205_3,  s_205_4,  s_205_5,  s_205_6,  s_205_7,  s_205_8;
wire  s_205_9, s_205_10, s_205_11, s_205_12, s_205_13, s_205_14;
wire s_205_15, s_205_16, s_205_17, s_205_18, s_205_19, s_205_20;
wire s_205_21, s_205_22, s_205_23, s_205_24, s_205_25, s_205_26;
wire  s_206_0,  s_206_1,  s_206_2,  s_206_3,  s_206_4,  s_206_5;
wire  s_206_6,  s_206_7,  s_206_8,  s_206_9, s_206_10, s_206_11;
wire s_206_12, s_206_13, s_206_14, s_206_15, s_206_16, s_206_17;
wire s_206_18, s_206_19, s_206_20, s_206_21, s_206_22, s_206_23;
wire s_206_24, s_206_25,  s_207_0,  s_207_1,  s_207_2,  s_207_3;
wire  s_207_4,  s_207_5,  s_207_6,  s_207_7,  s_207_8,  s_207_9;
wire s_207_10, s_207_11, s_207_12, s_207_13, s_207_14, s_207_15;
wire s_207_16, s_207_17, s_207_18, s_207_19, s_207_20, s_207_21;
wire s_207_22, s_207_23, s_207_24, s_207_25,  s_208_0,  s_208_1;
wire  s_208_2,  s_208_3,  s_208_4,  s_208_5,  s_208_6,  s_208_7;
wire  s_208_8,  s_208_9, s_208_10, s_208_11, s_208_12, s_208_13;
wire s_208_14, s_208_15, s_208_16, s_208_17, s_208_18, s_208_19;
wire s_208_20, s_208_21, s_208_22, s_208_23, s_208_24,  s_209_0;
wire  s_209_1,  s_209_2,  s_209_3,  s_209_4,  s_209_5,  s_209_6;
wire  s_209_7,  s_209_8,  s_209_9, s_209_10, s_209_11, s_209_12;
wire s_209_13, s_209_14, s_209_15, s_209_16, s_209_17, s_209_18;
wire s_209_19, s_209_20, s_209_21, s_209_22, s_209_23, s_209_24;
wire  s_210_0,  s_210_1,  s_210_2,  s_210_3,  s_210_4,  s_210_5;
wire  s_210_6,  s_210_7,  s_210_8,  s_210_9, s_210_10, s_210_11;
wire s_210_12, s_210_13, s_210_14, s_210_15, s_210_16, s_210_17;
wire s_210_18, s_210_19, s_210_20, s_210_21, s_210_22, s_210_23;
wire  s_211_0,  s_211_1,  s_211_2,  s_211_3,  s_211_4,  s_211_5;
wire  s_211_6,  s_211_7,  s_211_8,  s_211_9, s_211_10, s_211_11;
wire s_211_12, s_211_13, s_211_14, s_211_15, s_211_16, s_211_17;
wire s_211_18, s_211_19, s_211_20, s_211_21, s_211_22, s_211_23;
wire  s_212_0,  s_212_1,  s_212_2,  s_212_3,  s_212_4,  s_212_5;
wire  s_212_6,  s_212_7,  s_212_8,  s_212_9, s_212_10, s_212_11;
wire s_212_12, s_212_13, s_212_14, s_212_15, s_212_16, s_212_17;
wire s_212_18, s_212_19, s_212_20, s_212_21, s_212_22,  s_213_0;
wire  s_213_1,  s_213_2,  s_213_3,  s_213_4,  s_213_5,  s_213_6;
wire  s_213_7,  s_213_8,  s_213_9, s_213_10, s_213_11, s_213_12;
wire s_213_13, s_213_14, s_213_15, s_213_16, s_213_17, s_213_18;
wire s_213_19, s_213_20, s_213_21, s_213_22,  s_214_0,  s_214_1;
wire  s_214_2,  s_214_3,  s_214_4,  s_214_5,  s_214_6,  s_214_7;
wire  s_214_8,  s_214_9, s_214_10, s_214_11, s_214_12, s_214_13;
wire s_214_14, s_214_15, s_214_16, s_214_17, s_214_18, s_214_19;
wire s_214_20, s_214_21,  s_215_0,  s_215_1,  s_215_2,  s_215_3;
wire  s_215_4,  s_215_5,  s_215_6,  s_215_7,  s_215_8,  s_215_9;
wire s_215_10, s_215_11, s_215_12, s_215_13, s_215_14, s_215_15;
wire s_215_16, s_215_17, s_215_18, s_215_19, s_215_20, s_215_21;
wire  s_216_0,  s_216_1,  s_216_2,  s_216_3,  s_216_4,  s_216_5;
wire  s_216_6,  s_216_7,  s_216_8,  s_216_9, s_216_10, s_216_11;
wire s_216_12, s_216_13, s_216_14, s_216_15, s_216_16, s_216_17;
wire s_216_18, s_216_19, s_216_20,  s_217_0,  s_217_1,  s_217_2;
wire  s_217_3,  s_217_4,  s_217_5,  s_217_6,  s_217_7,  s_217_8;
wire  s_217_9, s_217_10, s_217_11, s_217_12, s_217_13, s_217_14;
wire s_217_15, s_217_16, s_217_17, s_217_18, s_217_19, s_217_20;
wire  s_218_0,  s_218_1,  s_218_2,  s_218_3,  s_218_4,  s_218_5;
wire  s_218_6,  s_218_7,  s_218_8,  s_218_9, s_218_10, s_218_11;
wire s_218_12, s_218_13, s_218_14, s_218_15, s_218_16, s_218_17;
wire s_218_18, s_218_19,  s_219_0,  s_219_1,  s_219_2,  s_219_3;
wire  s_219_4,  s_219_5,  s_219_6,  s_219_7,  s_219_8,  s_219_9;
wire s_219_10, s_219_11, s_219_12, s_219_13, s_219_14, s_219_15;
wire s_219_16, s_219_17, s_219_18, s_219_19,  s_220_0,  s_220_1;
wire  s_220_2,  s_220_3,  s_220_4,  s_220_5,  s_220_6,  s_220_7;
wire  s_220_8,  s_220_9, s_220_10, s_220_11, s_220_12, s_220_13;
wire s_220_14, s_220_15, s_220_16, s_220_17, s_220_18,  s_221_0;
wire  s_221_1,  s_221_2,  s_221_3,  s_221_4,  s_221_5,  s_221_6;
wire  s_221_7,  s_221_8,  s_221_9, s_221_10, s_221_11, s_221_12;
wire s_221_13, s_221_14, s_221_15, s_221_16, s_221_17, s_221_18;
wire  s_222_0,  s_222_1,  s_222_2,  s_222_3,  s_222_4,  s_222_5;
wire  s_222_6,  s_222_7,  s_222_8,  s_222_9, s_222_10, s_222_11;
wire s_222_12, s_222_13, s_222_14, s_222_15, s_222_16, s_222_17;
wire  s_223_0,  s_223_1,  s_223_2,  s_223_3,  s_223_4,  s_223_5;
wire  s_223_6,  s_223_7,  s_223_8,  s_223_9, s_223_10, s_223_11;
wire s_223_12, s_223_13, s_223_14, s_223_15, s_223_16, s_223_17;
wire  s_224_0,  s_224_1,  s_224_2,  s_224_3,  s_224_4,  s_224_5;
wire  s_224_6,  s_224_7,  s_224_8,  s_224_9, s_224_10, s_224_11;
wire s_224_12, s_224_13, s_224_14, s_224_15, s_224_16,  s_225_0;
wire  s_225_1,  s_225_2,  s_225_3,  s_225_4,  s_225_5,  s_225_6;
wire  s_225_7,  s_225_8,  s_225_9, s_225_10, s_225_11, s_225_12;
wire s_225_13, s_225_14, s_225_15, s_225_16,  s_226_0,  s_226_1;
wire  s_226_2,  s_226_3,  s_226_4,  s_226_5,  s_226_6,  s_226_7;
wire  s_226_8,  s_226_9, s_226_10, s_226_11, s_226_12, s_226_13;
wire s_226_14, s_226_15,  s_227_0,  s_227_1,  s_227_2,  s_227_3;
wire  s_227_4,  s_227_5,  s_227_6,  s_227_7,  s_227_8,  s_227_9;
wire s_227_10, s_227_11, s_227_12, s_227_13, s_227_14, s_227_15;
wire  s_228_0,  s_228_1,  s_228_2,  s_228_3,  s_228_4,  s_228_5;
wire  s_228_6,  s_228_7,  s_228_8,  s_228_9, s_228_10, s_228_11;
wire s_228_12, s_228_13, s_228_14,  s_229_0,  s_229_1,  s_229_2;
wire  s_229_3,  s_229_4,  s_229_5,  s_229_6,  s_229_7,  s_229_8;
wire  s_229_9, s_229_10, s_229_11, s_229_12, s_229_13, s_229_14;
wire  s_230_0,  s_230_1,  s_230_2,  s_230_3,  s_230_4,  s_230_5;
wire  s_230_6,  s_230_7,  s_230_8,  s_230_9, s_230_10, s_230_11;
wire s_230_12, s_230_13,  s_231_0,  s_231_1,  s_231_2,  s_231_3;
wire  s_231_4,  s_231_5,  s_231_6,  s_231_7,  s_231_8,  s_231_9;
wire s_231_10, s_231_11, s_231_12, s_231_13,  s_232_0,  s_232_1;
wire  s_232_2,  s_232_3,  s_232_4,  s_232_5,  s_232_6,  s_232_7;
wire  s_232_8,  s_232_9, s_232_10, s_232_11, s_232_12,  s_233_0;
wire  s_233_1,  s_233_2,  s_233_3,  s_233_4,  s_233_5,  s_233_6;
wire  s_233_7,  s_233_8,  s_233_9, s_233_10, s_233_11, s_233_12;
wire  s_234_0,  s_234_1,  s_234_2,  s_234_3,  s_234_4,  s_234_5;
wire  s_234_6,  s_234_7,  s_234_8,  s_234_9, s_234_10, s_234_11;
wire  s_235_0,  s_235_1,  s_235_2,  s_235_3,  s_235_4,  s_235_5;
wire  s_235_6,  s_235_7,  s_235_8,  s_235_9, s_235_10, s_235_11;
wire  s_236_0,  s_236_1,  s_236_2,  s_236_3,  s_236_4,  s_236_5;
wire  s_236_6,  s_236_7,  s_236_8,  s_236_9, s_236_10,  s_237_0;
wire  s_237_1,  s_237_2,  s_237_3,  s_237_4,  s_237_5,  s_237_6;
wire  s_237_7,  s_237_8,  s_237_9, s_237_10,  s_238_0,  s_238_1;
wire  s_238_2,  s_238_3,  s_238_4,  s_238_5,  s_238_6,  s_238_7;
wire  s_238_8,  s_238_9,  s_239_0,  s_239_1,  s_239_2,  s_239_3;
wire  s_239_4,  s_239_5,  s_239_6,  s_239_7,  s_239_8,  s_239_9;
wire  s_240_0,  s_240_1,  s_240_2,  s_240_3,  s_240_4,  s_240_5;
wire  s_240_6,  s_240_7,  s_240_8,  s_241_0,  s_241_1,  s_241_2;
wire  s_241_3,  s_241_4,  s_241_5,  s_241_6,  s_241_7,  s_241_8;
wire  s_242_0,  s_242_1,  s_242_2,  s_242_3,  s_242_4,  s_242_5;
wire  s_242_6,  s_242_7,  s_243_0,  s_243_1,  s_243_2,  s_243_3;
wire  s_243_4,  s_243_5,  s_243_6,  s_243_7,  s_244_0,  s_244_1;
wire  s_244_2,  s_244_3,  s_244_4,  s_244_5,  s_244_6,  s_245_0;
wire  s_245_1,  s_245_2,  s_245_3,  s_245_4,  s_245_5,  s_245_6;
wire  s_246_0,  s_246_1,  s_246_2,  s_246_3,  s_246_4,  s_246_5;
wire  s_247_0,  s_247_1,  s_247_2,  s_247_3,  s_247_4,  s_247_5;
wire  s_248_0,  s_248_1,  s_248_2,  s_248_3,  s_248_4,  s_249_0;
wire  s_249_1,  s_249_2,  s_249_3,  s_249_4,  s_250_0,  s_250_1;
wire  s_250_2,  s_250_3,  s_251_0,  s_251_1,  s_251_2,  s_251_3;
wire  s_252_0,  s_252_1,  s_252_2,  s_253_0,  s_253_1,  s_253_2;
wire  s_254_0,  s_254_1,  s_255_0,  s_255_1;

assign {
s_126_64, s_124_63, s_122_62, s_120_61, s_118_60, s_116_59, 
s_114_58, s_112_57, s_110_56, s_108_55, s_106_54, s_104_53, 
s_102_52, s_100_51,  s_98_50,  s_96_49,  s_94_48,  s_92_47, 
 s_90_46,  s_88_45,  s_86_44,  s_84_43,  s_82_42,  s_80_41, 
 s_78_40,  s_76_39,  s_74_38,  s_72_37,  s_70_36,  s_68_35, 
 s_66_34,  s_64_33,  s_62_32,  s_60_31,  s_58_30,  s_56_29, 
 s_54_28,  s_52_27,  s_50_26,  s_48_25,  s_46_24,  s_44_23, 
 s_42_22,  s_40_21,  s_38_20,  s_36_19,  s_34_18,  s_32_17, 
 s_30_16,  s_28_15,  s_26_14,  s_24_13,  s_22_12,  s_20_11, 
 s_18_10,   s_16_9,   s_14_8,   s_12_7,   s_10_6,    s_8_5, 
   s_6_4,    s_4_3,    s_2_2,    s_0_1
} = carry;

assign {
 s_129_0,  s_128_0,  s_127_0,  s_126_0,  s_125_0,  s_124_0, 
 s_123_0,  s_122_0,  s_121_0,  s_120_0,  s_119_0,  s_118_0, 
 s_117_0,  s_116_0,  s_115_0,  s_114_0,  s_113_0,  s_112_0, 
 s_111_0,  s_110_0,  s_109_0,  s_108_0,  s_107_0,  s_106_0, 
 s_105_0,  s_104_0,  s_103_0,  s_102_0,  s_101_0,  s_100_0, 
  s_99_0,   s_98_0,   s_97_0,   s_96_0,   s_95_0,   s_94_0, 
  s_93_0,   s_92_0,   s_91_0,   s_90_0,   s_89_0,   s_88_0, 
  s_87_0,   s_86_0,   s_85_0,   s_84_0,   s_83_0,   s_82_0, 
  s_81_0,   s_80_0,   s_79_0,   s_78_0,   s_77_0,   s_76_0, 
  s_75_0,   s_74_0,   s_73_0,   s_72_0,   s_71_0,   s_70_0, 
  s_69_0,   s_68_0,   s_67_0,   s_66_0,   s_65_0,   s_64_0, 
  s_63_0,   s_62_0,   s_61_0,   s_60_0,   s_59_0,   s_58_0, 
  s_57_0,   s_56_0,   s_55_0,   s_54_0,   s_53_0,   s_52_0, 
  s_51_0,   s_50_0,   s_49_0,   s_48_0,   s_47_0,   s_46_0, 
  s_45_0,   s_44_0,   s_43_0,   s_42_0,   s_41_0,   s_40_0, 
  s_39_0,   s_38_0,   s_37_0,   s_36_0,   s_35_0,   s_34_0, 
  s_33_0,   s_32_0,   s_31_0,   s_30_0,   s_29_0,   s_28_0, 
  s_27_0,   s_26_0,   s_25_0,   s_24_0,   s_23_0,   s_22_0, 
  s_21_0,   s_20_0,   s_19_0,   s_18_0,   s_17_0,   s_16_0, 
  s_15_0,   s_14_0,   s_13_0,   s_12_0,   s_11_0,   s_10_0, 
   s_9_0,    s_8_0,    s_7_0,    s_6_0,    s_5_0,    s_4_0, 
   s_3_0,    s_2_0,    s_1_0,    s_0_0
} = partial_products[(width+2)*(0+1)-1:(width+2)*0];

assign {
 s_131_0,  s_130_0,  s_129_1,  s_128_1,  s_127_1,  s_126_1, 
 s_125_1,  s_124_1,  s_123_1,  s_122_1,  s_121_1,  s_120_1, 
 s_119_1,  s_118_1,  s_117_1,  s_116_1,  s_115_1,  s_114_1, 
 s_113_1,  s_112_1,  s_111_1,  s_110_1,  s_109_1,  s_108_1, 
 s_107_1,  s_106_1,  s_105_1,  s_104_1,  s_103_1,  s_102_1, 
 s_101_1,  s_100_1,   s_99_1,   s_98_1,   s_97_1,   s_96_1, 
  s_95_1,   s_94_1,   s_93_1,   s_92_1,   s_91_1,   s_90_1, 
  s_89_1,   s_88_1,   s_87_1,   s_86_1,   s_85_1,   s_84_1, 
  s_83_1,   s_82_1,   s_81_1,   s_80_1,   s_79_1,   s_78_1, 
  s_77_1,   s_76_1,   s_75_1,   s_74_1,   s_73_1,   s_72_1, 
  s_71_1,   s_70_1,   s_69_1,   s_68_1,   s_67_1,   s_66_1, 
  s_65_1,   s_64_1,   s_63_1,   s_62_1,   s_61_1,   s_60_1, 
  s_59_1,   s_58_1,   s_57_1,   s_56_1,   s_55_1,   s_54_1, 
  s_53_1,   s_52_1,   s_51_1,   s_50_1,   s_49_1,   s_48_1, 
  s_47_1,   s_46_1,   s_45_1,   s_44_1,   s_43_1,   s_42_1, 
  s_41_1,   s_40_1,   s_39_1,   s_38_1,   s_37_1,   s_36_1, 
  s_35_1,   s_34_1,   s_33_1,   s_32_1,   s_31_1,   s_30_1, 
  s_29_1,   s_28_1,   s_27_1,   s_26_1,   s_25_1,   s_24_1, 
  s_23_1,   s_22_1,   s_21_1,   s_20_1,   s_19_1,   s_18_1, 
  s_17_1,   s_16_1,   s_15_1,   s_14_1,   s_13_1,   s_12_1, 
  s_11_1,   s_10_1,    s_9_1,    s_8_1,    s_7_1,    s_6_1, 
   s_5_1,    s_4_1,    s_3_1,    s_2_1
} = partial_products[(width+2)*(1+1)-1:(width+2)*1];

assign {
 s_133_0,  s_132_0,  s_131_1,  s_130_1,  s_129_2,  s_128_2, 
 s_127_2,  s_126_2,  s_125_2,  s_124_2,  s_123_2,  s_122_2, 
 s_121_2,  s_120_2,  s_119_2,  s_118_2,  s_117_2,  s_116_2, 
 s_115_2,  s_114_2,  s_113_2,  s_112_2,  s_111_2,  s_110_2, 
 s_109_2,  s_108_2,  s_107_2,  s_106_2,  s_105_2,  s_104_2, 
 s_103_2,  s_102_2,  s_101_2,  s_100_2,   s_99_2,   s_98_2, 
  s_97_2,   s_96_2,   s_95_2,   s_94_2,   s_93_2,   s_92_2, 
  s_91_2,   s_90_2,   s_89_2,   s_88_2,   s_87_2,   s_86_2, 
  s_85_2,   s_84_2,   s_83_2,   s_82_2,   s_81_2,   s_80_2, 
  s_79_2,   s_78_2,   s_77_2,   s_76_2,   s_75_2,   s_74_2, 
  s_73_2,   s_72_2,   s_71_2,   s_70_2,   s_69_2,   s_68_2, 
  s_67_2,   s_66_2,   s_65_2,   s_64_2,   s_63_2,   s_62_2, 
  s_61_2,   s_60_2,   s_59_2,   s_58_2,   s_57_2,   s_56_2, 
  s_55_2,   s_54_2,   s_53_2,   s_52_2,   s_51_2,   s_50_2, 
  s_49_2,   s_48_2,   s_47_2,   s_46_2,   s_45_2,   s_44_2, 
  s_43_2,   s_42_2,   s_41_2,   s_40_2,   s_39_2,   s_38_2, 
  s_37_2,   s_36_2,   s_35_2,   s_34_2,   s_33_2,   s_32_2, 
  s_31_2,   s_30_2,   s_29_2,   s_28_2,   s_27_2,   s_26_2, 
  s_25_2,   s_24_2,   s_23_2,   s_22_2,   s_21_2,   s_20_2, 
  s_19_2,   s_18_2,   s_17_2,   s_16_2,   s_15_2,   s_14_2, 
  s_13_2,   s_12_2,   s_11_2,   s_10_2,    s_9_2,    s_8_2, 
   s_7_2,    s_6_2,    s_5_2,    s_4_2
} = partial_products[(width+2)*(2+1)-1:(width+2)*2];

assign {
 s_135_0,  s_134_0,  s_133_1,  s_132_1,  s_131_2,  s_130_2, 
 s_129_3,  s_128_3,  s_127_3,  s_126_3,  s_125_3,  s_124_3, 
 s_123_3,  s_122_3,  s_121_3,  s_120_3,  s_119_3,  s_118_3, 
 s_117_3,  s_116_3,  s_115_3,  s_114_3,  s_113_3,  s_112_3, 
 s_111_3,  s_110_3,  s_109_3,  s_108_3,  s_107_3,  s_106_3, 
 s_105_3,  s_104_3,  s_103_3,  s_102_3,  s_101_3,  s_100_3, 
  s_99_3,   s_98_3,   s_97_3,   s_96_3,   s_95_3,   s_94_3, 
  s_93_3,   s_92_3,   s_91_3,   s_90_3,   s_89_3,   s_88_3, 
  s_87_3,   s_86_3,   s_85_3,   s_84_3,   s_83_3,   s_82_3, 
  s_81_3,   s_80_3,   s_79_3,   s_78_3,   s_77_3,   s_76_3, 
  s_75_3,   s_74_3,   s_73_3,   s_72_3,   s_71_3,   s_70_3, 
  s_69_3,   s_68_3,   s_67_3,   s_66_3,   s_65_3,   s_64_3, 
  s_63_3,   s_62_3,   s_61_3,   s_60_3,   s_59_3,   s_58_3, 
  s_57_3,   s_56_3,   s_55_3,   s_54_3,   s_53_3,   s_52_3, 
  s_51_3,   s_50_3,   s_49_3,   s_48_3,   s_47_3,   s_46_3, 
  s_45_3,   s_44_3,   s_43_3,   s_42_3,   s_41_3,   s_40_3, 
  s_39_3,   s_38_3,   s_37_3,   s_36_3,   s_35_3,   s_34_3, 
  s_33_3,   s_32_3,   s_31_3,   s_30_3,   s_29_3,   s_28_3, 
  s_27_3,   s_26_3,   s_25_3,   s_24_3,   s_23_3,   s_22_3, 
  s_21_3,   s_20_3,   s_19_3,   s_18_3,   s_17_3,   s_16_3, 
  s_15_3,   s_14_3,   s_13_3,   s_12_3,   s_11_3,   s_10_3, 
   s_9_3,    s_8_3,    s_7_3,    s_6_3
} = partial_products[(width+2)*(3+1)-1:(width+2)*3];

assign {
 s_137_0,  s_136_0,  s_135_1,  s_134_1,  s_133_2,  s_132_2, 
 s_131_3,  s_130_3,  s_129_4,  s_128_4,  s_127_4,  s_126_4, 
 s_125_4,  s_124_4,  s_123_4,  s_122_4,  s_121_4,  s_120_4, 
 s_119_4,  s_118_4,  s_117_4,  s_116_4,  s_115_4,  s_114_4, 
 s_113_4,  s_112_4,  s_111_4,  s_110_4,  s_109_4,  s_108_4, 
 s_107_4,  s_106_4,  s_105_4,  s_104_4,  s_103_4,  s_102_4, 
 s_101_4,  s_100_4,   s_99_4,   s_98_4,   s_97_4,   s_96_4, 
  s_95_4,   s_94_4,   s_93_4,   s_92_4,   s_91_4,   s_90_4, 
  s_89_4,   s_88_4,   s_87_4,   s_86_4,   s_85_4,   s_84_4, 
  s_83_4,   s_82_4,   s_81_4,   s_80_4,   s_79_4,   s_78_4, 
  s_77_4,   s_76_4,   s_75_4,   s_74_4,   s_73_4,   s_72_4, 
  s_71_4,   s_70_4,   s_69_4,   s_68_4,   s_67_4,   s_66_4, 
  s_65_4,   s_64_4,   s_63_4,   s_62_4,   s_61_4,   s_60_4, 
  s_59_4,   s_58_4,   s_57_4,   s_56_4,   s_55_4,   s_54_4, 
  s_53_4,   s_52_4,   s_51_4,   s_50_4,   s_49_4,   s_48_4, 
  s_47_4,   s_46_4,   s_45_4,   s_44_4,   s_43_4,   s_42_4, 
  s_41_4,   s_40_4,   s_39_4,   s_38_4,   s_37_4,   s_36_4, 
  s_35_4,   s_34_4,   s_33_4,   s_32_4,   s_31_4,   s_30_4, 
  s_29_4,   s_28_4,   s_27_4,   s_26_4,   s_25_4,   s_24_4, 
  s_23_4,   s_22_4,   s_21_4,   s_20_4,   s_19_4,   s_18_4, 
  s_17_4,   s_16_4,   s_15_4,   s_14_4,   s_13_4,   s_12_4, 
  s_11_4,   s_10_4,    s_9_4,    s_8_4
} = partial_products[(width+2)*(4+1)-1:(width+2)*4];

assign {
 s_139_0,  s_138_0,  s_137_1,  s_136_1,  s_135_2,  s_134_2, 
 s_133_3,  s_132_3,  s_131_4,  s_130_4,  s_129_5,  s_128_5, 
 s_127_5,  s_126_5,  s_125_5,  s_124_5,  s_123_5,  s_122_5, 
 s_121_5,  s_120_5,  s_119_5,  s_118_5,  s_117_5,  s_116_5, 
 s_115_5,  s_114_5,  s_113_5,  s_112_5,  s_111_5,  s_110_5, 
 s_109_5,  s_108_5,  s_107_5,  s_106_5,  s_105_5,  s_104_5, 
 s_103_5,  s_102_5,  s_101_5,  s_100_5,   s_99_5,   s_98_5, 
  s_97_5,   s_96_5,   s_95_5,   s_94_5,   s_93_5,   s_92_5, 
  s_91_5,   s_90_5,   s_89_5,   s_88_5,   s_87_5,   s_86_5, 
  s_85_5,   s_84_5,   s_83_5,   s_82_5,   s_81_5,   s_80_5, 
  s_79_5,   s_78_5,   s_77_5,   s_76_5,   s_75_5,   s_74_5, 
  s_73_5,   s_72_5,   s_71_5,   s_70_5,   s_69_5,   s_68_5, 
  s_67_5,   s_66_5,   s_65_5,   s_64_5,   s_63_5,   s_62_5, 
  s_61_5,   s_60_5,   s_59_5,   s_58_5,   s_57_5,   s_56_5, 
  s_55_5,   s_54_5,   s_53_5,   s_52_5,   s_51_5,   s_50_5, 
  s_49_5,   s_48_5,   s_47_5,   s_46_5,   s_45_5,   s_44_5, 
  s_43_5,   s_42_5,   s_41_5,   s_40_5,   s_39_5,   s_38_5, 
  s_37_5,   s_36_5,   s_35_5,   s_34_5,   s_33_5,   s_32_5, 
  s_31_5,   s_30_5,   s_29_5,   s_28_5,   s_27_5,   s_26_5, 
  s_25_5,   s_24_5,   s_23_5,   s_22_5,   s_21_5,   s_20_5, 
  s_19_5,   s_18_5,   s_17_5,   s_16_5,   s_15_5,   s_14_5, 
  s_13_5,   s_12_5,   s_11_5,   s_10_5
} = partial_products[(width+2)*(5+1)-1:(width+2)*5];

assign {
 s_141_0,  s_140_0,  s_139_1,  s_138_1,  s_137_2,  s_136_2, 
 s_135_3,  s_134_3,  s_133_4,  s_132_4,  s_131_5,  s_130_5, 
 s_129_6,  s_128_6,  s_127_6,  s_126_6,  s_125_6,  s_124_6, 
 s_123_6,  s_122_6,  s_121_6,  s_120_6,  s_119_6,  s_118_6, 
 s_117_6,  s_116_6,  s_115_6,  s_114_6,  s_113_6,  s_112_6, 
 s_111_6,  s_110_6,  s_109_6,  s_108_6,  s_107_6,  s_106_6, 
 s_105_6,  s_104_6,  s_103_6,  s_102_6,  s_101_6,  s_100_6, 
  s_99_6,   s_98_6,   s_97_6,   s_96_6,   s_95_6,   s_94_6, 
  s_93_6,   s_92_6,   s_91_6,   s_90_6,   s_89_6,   s_88_6, 
  s_87_6,   s_86_6,   s_85_6,   s_84_6,   s_83_6,   s_82_6, 
  s_81_6,   s_80_6,   s_79_6,   s_78_6,   s_77_6,   s_76_6, 
  s_75_6,   s_74_6,   s_73_6,   s_72_6,   s_71_6,   s_70_6, 
  s_69_6,   s_68_6,   s_67_6,   s_66_6,   s_65_6,   s_64_6, 
  s_63_6,   s_62_6,   s_61_6,   s_60_6,   s_59_6,   s_58_6, 
  s_57_6,   s_56_6,   s_55_6,   s_54_6,   s_53_6,   s_52_6, 
  s_51_6,   s_50_6,   s_49_6,   s_48_6,   s_47_6,   s_46_6, 
  s_45_6,   s_44_6,   s_43_6,   s_42_6,   s_41_6,   s_40_6, 
  s_39_6,   s_38_6,   s_37_6,   s_36_6,   s_35_6,   s_34_6, 
  s_33_6,   s_32_6,   s_31_6,   s_30_6,   s_29_6,   s_28_6, 
  s_27_6,   s_26_6,   s_25_6,   s_24_6,   s_23_6,   s_22_6, 
  s_21_6,   s_20_6,   s_19_6,   s_18_6,   s_17_6,   s_16_6, 
  s_15_6,   s_14_6,   s_13_6,   s_12_6
} = partial_products[(width+2)*(6+1)-1:(width+2)*6];

assign {
 s_143_0,  s_142_0,  s_141_1,  s_140_1,  s_139_2,  s_138_2, 
 s_137_3,  s_136_3,  s_135_4,  s_134_4,  s_133_5,  s_132_5, 
 s_131_6,  s_130_6,  s_129_7,  s_128_7,  s_127_7,  s_126_7, 
 s_125_7,  s_124_7,  s_123_7,  s_122_7,  s_121_7,  s_120_7, 
 s_119_7,  s_118_7,  s_117_7,  s_116_7,  s_115_7,  s_114_7, 
 s_113_7,  s_112_7,  s_111_7,  s_110_7,  s_109_7,  s_108_7, 
 s_107_7,  s_106_7,  s_105_7,  s_104_7,  s_103_7,  s_102_7, 
 s_101_7,  s_100_7,   s_99_7,   s_98_7,   s_97_7,   s_96_7, 
  s_95_7,   s_94_7,   s_93_7,   s_92_7,   s_91_7,   s_90_7, 
  s_89_7,   s_88_7,   s_87_7,   s_86_7,   s_85_7,   s_84_7, 
  s_83_7,   s_82_7,   s_81_7,   s_80_7,   s_79_7,   s_78_7, 
  s_77_7,   s_76_7,   s_75_7,   s_74_7,   s_73_7,   s_72_7, 
  s_71_7,   s_70_7,   s_69_7,   s_68_7,   s_67_7,   s_66_7, 
  s_65_7,   s_64_7,   s_63_7,   s_62_7,   s_61_7,   s_60_7, 
  s_59_7,   s_58_7,   s_57_7,   s_56_7,   s_55_7,   s_54_7, 
  s_53_7,   s_52_7,   s_51_7,   s_50_7,   s_49_7,   s_48_7, 
  s_47_7,   s_46_7,   s_45_7,   s_44_7,   s_43_7,   s_42_7, 
  s_41_7,   s_40_7,   s_39_7,   s_38_7,   s_37_7,   s_36_7, 
  s_35_7,   s_34_7,   s_33_7,   s_32_7,   s_31_7,   s_30_7, 
  s_29_7,   s_28_7,   s_27_7,   s_26_7,   s_25_7,   s_24_7, 
  s_23_7,   s_22_7,   s_21_7,   s_20_7,   s_19_7,   s_18_7, 
  s_17_7,   s_16_7,   s_15_7,   s_14_7
} = partial_products[(width+2)*(7+1)-1:(width+2)*7];

assign {
 s_145_0,  s_144_0,  s_143_1,  s_142_1,  s_141_2,  s_140_2, 
 s_139_3,  s_138_3,  s_137_4,  s_136_4,  s_135_5,  s_134_5, 
 s_133_6,  s_132_6,  s_131_7,  s_130_7,  s_129_8,  s_128_8, 
 s_127_8,  s_126_8,  s_125_8,  s_124_8,  s_123_8,  s_122_8, 
 s_121_8,  s_120_8,  s_119_8,  s_118_8,  s_117_8,  s_116_8, 
 s_115_8,  s_114_8,  s_113_8,  s_112_8,  s_111_8,  s_110_8, 
 s_109_8,  s_108_8,  s_107_8,  s_106_8,  s_105_8,  s_104_8, 
 s_103_8,  s_102_8,  s_101_8,  s_100_8,   s_99_8,   s_98_8, 
  s_97_8,   s_96_8,   s_95_8,   s_94_8,   s_93_8,   s_92_8, 
  s_91_8,   s_90_8,   s_89_8,   s_88_8,   s_87_8,   s_86_8, 
  s_85_8,   s_84_8,   s_83_8,   s_82_8,   s_81_8,   s_80_8, 
  s_79_8,   s_78_8,   s_77_8,   s_76_8,   s_75_8,   s_74_8, 
  s_73_8,   s_72_8,   s_71_8,   s_70_8,   s_69_8,   s_68_8, 
  s_67_8,   s_66_8,   s_65_8,   s_64_8,   s_63_8,   s_62_8, 
  s_61_8,   s_60_8,   s_59_8,   s_58_8,   s_57_8,   s_56_8, 
  s_55_8,   s_54_8,   s_53_8,   s_52_8,   s_51_8,   s_50_8, 
  s_49_8,   s_48_8,   s_47_8,   s_46_8,   s_45_8,   s_44_8, 
  s_43_8,   s_42_8,   s_41_8,   s_40_8,   s_39_8,   s_38_8, 
  s_37_8,   s_36_8,   s_35_8,   s_34_8,   s_33_8,   s_32_8, 
  s_31_8,   s_30_8,   s_29_8,   s_28_8,   s_27_8,   s_26_8, 
  s_25_8,   s_24_8,   s_23_8,   s_22_8,   s_21_8,   s_20_8, 
  s_19_8,   s_18_8,   s_17_8,   s_16_8
} = partial_products[(width+2)*(8+1)-1:(width+2)*8];

assign {
 s_147_0,  s_146_0,  s_145_1,  s_144_1,  s_143_2,  s_142_2, 
 s_141_3,  s_140_3,  s_139_4,  s_138_4,  s_137_5,  s_136_5, 
 s_135_6,  s_134_6,  s_133_7,  s_132_7,  s_131_8,  s_130_8, 
 s_129_9,  s_128_9,  s_127_9,  s_126_9,  s_125_9,  s_124_9, 
 s_123_9,  s_122_9,  s_121_9,  s_120_9,  s_119_9,  s_118_9, 
 s_117_9,  s_116_9,  s_115_9,  s_114_9,  s_113_9,  s_112_9, 
 s_111_9,  s_110_9,  s_109_9,  s_108_9,  s_107_9,  s_106_9, 
 s_105_9,  s_104_9,  s_103_9,  s_102_9,  s_101_9,  s_100_9, 
  s_99_9,   s_98_9,   s_97_9,   s_96_9,   s_95_9,   s_94_9, 
  s_93_9,   s_92_9,   s_91_9,   s_90_9,   s_89_9,   s_88_9, 
  s_87_9,   s_86_9,   s_85_9,   s_84_9,   s_83_9,   s_82_9, 
  s_81_9,   s_80_9,   s_79_9,   s_78_9,   s_77_9,   s_76_9, 
  s_75_9,   s_74_9,   s_73_9,   s_72_9,   s_71_9,   s_70_9, 
  s_69_9,   s_68_9,   s_67_9,   s_66_9,   s_65_9,   s_64_9, 
  s_63_9,   s_62_9,   s_61_9,   s_60_9,   s_59_9,   s_58_9, 
  s_57_9,   s_56_9,   s_55_9,   s_54_9,   s_53_9,   s_52_9, 
  s_51_9,   s_50_9,   s_49_9,   s_48_9,   s_47_9,   s_46_9, 
  s_45_9,   s_44_9,   s_43_9,   s_42_9,   s_41_9,   s_40_9, 
  s_39_9,   s_38_9,   s_37_9,   s_36_9,   s_35_9,   s_34_9, 
  s_33_9,   s_32_9,   s_31_9,   s_30_9,   s_29_9,   s_28_9, 
  s_27_9,   s_26_9,   s_25_9,   s_24_9,   s_23_9,   s_22_9, 
  s_21_9,   s_20_9,   s_19_9,   s_18_9
} = partial_products[(width+2)*(9+1)-1:(width+2)*9];

assign {
 s_149_0,  s_148_0,  s_147_1,  s_146_1,  s_145_2,  s_144_2, 
 s_143_3,  s_142_3,  s_141_4,  s_140_4,  s_139_5,  s_138_5, 
 s_137_6,  s_136_6,  s_135_7,  s_134_7,  s_133_8,  s_132_8, 
 s_131_9,  s_130_9, s_129_10, s_128_10, s_127_10, s_126_10, 
s_125_10, s_124_10, s_123_10, s_122_10, s_121_10, s_120_10, 
s_119_10, s_118_10, s_117_10, s_116_10, s_115_10, s_114_10, 
s_113_10, s_112_10, s_111_10, s_110_10, s_109_10, s_108_10, 
s_107_10, s_106_10, s_105_10, s_104_10, s_103_10, s_102_10, 
s_101_10, s_100_10,  s_99_10,  s_98_10,  s_97_10,  s_96_10, 
 s_95_10,  s_94_10,  s_93_10,  s_92_10,  s_91_10,  s_90_10, 
 s_89_10,  s_88_10,  s_87_10,  s_86_10,  s_85_10,  s_84_10, 
 s_83_10,  s_82_10,  s_81_10,  s_80_10,  s_79_10,  s_78_10, 
 s_77_10,  s_76_10,  s_75_10,  s_74_10,  s_73_10,  s_72_10, 
 s_71_10,  s_70_10,  s_69_10,  s_68_10,  s_67_10,  s_66_10, 
 s_65_10,  s_64_10,  s_63_10,  s_62_10,  s_61_10,  s_60_10, 
 s_59_10,  s_58_10,  s_57_10,  s_56_10,  s_55_10,  s_54_10, 
 s_53_10,  s_52_10,  s_51_10,  s_50_10,  s_49_10,  s_48_10, 
 s_47_10,  s_46_10,  s_45_10,  s_44_10,  s_43_10,  s_42_10, 
 s_41_10,  s_40_10,  s_39_10,  s_38_10,  s_37_10,  s_36_10, 
 s_35_10,  s_34_10,  s_33_10,  s_32_10,  s_31_10,  s_30_10, 
 s_29_10,  s_28_10,  s_27_10,  s_26_10,  s_25_10,  s_24_10, 
 s_23_10,  s_22_10,  s_21_10,  s_20_10
} = partial_products[(width+2)*(10+1)-1:(width+2)*10];

assign {
 s_151_0,  s_150_0,  s_149_1,  s_148_1,  s_147_2,  s_146_2, 
 s_145_3,  s_144_3,  s_143_4,  s_142_4,  s_141_5,  s_140_5, 
 s_139_6,  s_138_6,  s_137_7,  s_136_7,  s_135_8,  s_134_8, 
 s_133_9,  s_132_9, s_131_10, s_130_10, s_129_11, s_128_11, 
s_127_11, s_126_11, s_125_11, s_124_11, s_123_11, s_122_11, 
s_121_11, s_120_11, s_119_11, s_118_11, s_117_11, s_116_11, 
s_115_11, s_114_11, s_113_11, s_112_11, s_111_11, s_110_11, 
s_109_11, s_108_11, s_107_11, s_106_11, s_105_11, s_104_11, 
s_103_11, s_102_11, s_101_11, s_100_11,  s_99_11,  s_98_11, 
 s_97_11,  s_96_11,  s_95_11,  s_94_11,  s_93_11,  s_92_11, 
 s_91_11,  s_90_11,  s_89_11,  s_88_11,  s_87_11,  s_86_11, 
 s_85_11,  s_84_11,  s_83_11,  s_82_11,  s_81_11,  s_80_11, 
 s_79_11,  s_78_11,  s_77_11,  s_76_11,  s_75_11,  s_74_11, 
 s_73_11,  s_72_11,  s_71_11,  s_70_11,  s_69_11,  s_68_11, 
 s_67_11,  s_66_11,  s_65_11,  s_64_11,  s_63_11,  s_62_11, 
 s_61_11,  s_60_11,  s_59_11,  s_58_11,  s_57_11,  s_56_11, 
 s_55_11,  s_54_11,  s_53_11,  s_52_11,  s_51_11,  s_50_11, 
 s_49_11,  s_48_11,  s_47_11,  s_46_11,  s_45_11,  s_44_11, 
 s_43_11,  s_42_11,  s_41_11,  s_40_11,  s_39_11,  s_38_11, 
 s_37_11,  s_36_11,  s_35_11,  s_34_11,  s_33_11,  s_32_11, 
 s_31_11,  s_30_11,  s_29_11,  s_28_11,  s_27_11,  s_26_11, 
 s_25_11,  s_24_11,  s_23_11,  s_22_11
} = partial_products[(width+2)*(11+1)-1:(width+2)*11];

assign {
 s_153_0,  s_152_0,  s_151_1,  s_150_1,  s_149_2,  s_148_2, 
 s_147_3,  s_146_3,  s_145_4,  s_144_4,  s_143_5,  s_142_5, 
 s_141_6,  s_140_6,  s_139_7,  s_138_7,  s_137_8,  s_136_8, 
 s_135_9,  s_134_9, s_133_10, s_132_10, s_131_11, s_130_11, 
s_129_12, s_128_12, s_127_12, s_126_12, s_125_12, s_124_12, 
s_123_12, s_122_12, s_121_12, s_120_12, s_119_12, s_118_12, 
s_117_12, s_116_12, s_115_12, s_114_12, s_113_12, s_112_12, 
s_111_12, s_110_12, s_109_12, s_108_12, s_107_12, s_106_12, 
s_105_12, s_104_12, s_103_12, s_102_12, s_101_12, s_100_12, 
 s_99_12,  s_98_12,  s_97_12,  s_96_12,  s_95_12,  s_94_12, 
 s_93_12,  s_92_12,  s_91_12,  s_90_12,  s_89_12,  s_88_12, 
 s_87_12,  s_86_12,  s_85_12,  s_84_12,  s_83_12,  s_82_12, 
 s_81_12,  s_80_12,  s_79_12,  s_78_12,  s_77_12,  s_76_12, 
 s_75_12,  s_74_12,  s_73_12,  s_72_12,  s_71_12,  s_70_12, 
 s_69_12,  s_68_12,  s_67_12,  s_66_12,  s_65_12,  s_64_12, 
 s_63_12,  s_62_12,  s_61_12,  s_60_12,  s_59_12,  s_58_12, 
 s_57_12,  s_56_12,  s_55_12,  s_54_12,  s_53_12,  s_52_12, 
 s_51_12,  s_50_12,  s_49_12,  s_48_12,  s_47_12,  s_46_12, 
 s_45_12,  s_44_12,  s_43_12,  s_42_12,  s_41_12,  s_40_12, 
 s_39_12,  s_38_12,  s_37_12,  s_36_12,  s_35_12,  s_34_12, 
 s_33_12,  s_32_12,  s_31_12,  s_30_12,  s_29_12,  s_28_12, 
 s_27_12,  s_26_12,  s_25_12,  s_24_12
} = partial_products[(width+2)*(12+1)-1:(width+2)*12];

assign {
 s_155_0,  s_154_0,  s_153_1,  s_152_1,  s_151_2,  s_150_2, 
 s_149_3,  s_148_3,  s_147_4,  s_146_4,  s_145_5,  s_144_5, 
 s_143_6,  s_142_6,  s_141_7,  s_140_7,  s_139_8,  s_138_8, 
 s_137_9,  s_136_9, s_135_10, s_134_10, s_133_11, s_132_11, 
s_131_12, s_130_12, s_129_13, s_128_13, s_127_13, s_126_13, 
s_125_13, s_124_13, s_123_13, s_122_13, s_121_13, s_120_13, 
s_119_13, s_118_13, s_117_13, s_116_13, s_115_13, s_114_13, 
s_113_13, s_112_13, s_111_13, s_110_13, s_109_13, s_108_13, 
s_107_13, s_106_13, s_105_13, s_104_13, s_103_13, s_102_13, 
s_101_13, s_100_13,  s_99_13,  s_98_13,  s_97_13,  s_96_13, 
 s_95_13,  s_94_13,  s_93_13,  s_92_13,  s_91_13,  s_90_13, 
 s_89_13,  s_88_13,  s_87_13,  s_86_13,  s_85_13,  s_84_13, 
 s_83_13,  s_82_13,  s_81_13,  s_80_13,  s_79_13,  s_78_13, 
 s_77_13,  s_76_13,  s_75_13,  s_74_13,  s_73_13,  s_72_13, 
 s_71_13,  s_70_13,  s_69_13,  s_68_13,  s_67_13,  s_66_13, 
 s_65_13,  s_64_13,  s_63_13,  s_62_13,  s_61_13,  s_60_13, 
 s_59_13,  s_58_13,  s_57_13,  s_56_13,  s_55_13,  s_54_13, 
 s_53_13,  s_52_13,  s_51_13,  s_50_13,  s_49_13,  s_48_13, 
 s_47_13,  s_46_13,  s_45_13,  s_44_13,  s_43_13,  s_42_13, 
 s_41_13,  s_40_13,  s_39_13,  s_38_13,  s_37_13,  s_36_13, 
 s_35_13,  s_34_13,  s_33_13,  s_32_13,  s_31_13,  s_30_13, 
 s_29_13,  s_28_13,  s_27_13,  s_26_13
} = partial_products[(width+2)*(13+1)-1:(width+2)*13];

assign {
 s_157_0,  s_156_0,  s_155_1,  s_154_1,  s_153_2,  s_152_2, 
 s_151_3,  s_150_3,  s_149_4,  s_148_4,  s_147_5,  s_146_5, 
 s_145_6,  s_144_6,  s_143_7,  s_142_7,  s_141_8,  s_140_8, 
 s_139_9,  s_138_9, s_137_10, s_136_10, s_135_11, s_134_11, 
s_133_12, s_132_12, s_131_13, s_130_13, s_129_14, s_128_14, 
s_127_14, s_126_14, s_125_14, s_124_14, s_123_14, s_122_14, 
s_121_14, s_120_14, s_119_14, s_118_14, s_117_14, s_116_14, 
s_115_14, s_114_14, s_113_14, s_112_14, s_111_14, s_110_14, 
s_109_14, s_108_14, s_107_14, s_106_14, s_105_14, s_104_14, 
s_103_14, s_102_14, s_101_14, s_100_14,  s_99_14,  s_98_14, 
 s_97_14,  s_96_14,  s_95_14,  s_94_14,  s_93_14,  s_92_14, 
 s_91_14,  s_90_14,  s_89_14,  s_88_14,  s_87_14,  s_86_14, 
 s_85_14,  s_84_14,  s_83_14,  s_82_14,  s_81_14,  s_80_14, 
 s_79_14,  s_78_14,  s_77_14,  s_76_14,  s_75_14,  s_74_14, 
 s_73_14,  s_72_14,  s_71_14,  s_70_14,  s_69_14,  s_68_14, 
 s_67_14,  s_66_14,  s_65_14,  s_64_14,  s_63_14,  s_62_14, 
 s_61_14,  s_60_14,  s_59_14,  s_58_14,  s_57_14,  s_56_14, 
 s_55_14,  s_54_14,  s_53_14,  s_52_14,  s_51_14,  s_50_14, 
 s_49_14,  s_48_14,  s_47_14,  s_46_14,  s_45_14,  s_44_14, 
 s_43_14,  s_42_14,  s_41_14,  s_40_14,  s_39_14,  s_38_14, 
 s_37_14,  s_36_14,  s_35_14,  s_34_14,  s_33_14,  s_32_14, 
 s_31_14,  s_30_14,  s_29_14,  s_28_14
} = partial_products[(width+2)*(14+1)-1:(width+2)*14];

assign {
 s_159_0,  s_158_0,  s_157_1,  s_156_1,  s_155_2,  s_154_2, 
 s_153_3,  s_152_3,  s_151_4,  s_150_4,  s_149_5,  s_148_5, 
 s_147_6,  s_146_6,  s_145_7,  s_144_7,  s_143_8,  s_142_8, 
 s_141_9,  s_140_9, s_139_10, s_138_10, s_137_11, s_136_11, 
s_135_12, s_134_12, s_133_13, s_132_13, s_131_14, s_130_14, 
s_129_15, s_128_15, s_127_15, s_126_15, s_125_15, s_124_15, 
s_123_15, s_122_15, s_121_15, s_120_15, s_119_15, s_118_15, 
s_117_15, s_116_15, s_115_15, s_114_15, s_113_15, s_112_15, 
s_111_15, s_110_15, s_109_15, s_108_15, s_107_15, s_106_15, 
s_105_15, s_104_15, s_103_15, s_102_15, s_101_15, s_100_15, 
 s_99_15,  s_98_15,  s_97_15,  s_96_15,  s_95_15,  s_94_15, 
 s_93_15,  s_92_15,  s_91_15,  s_90_15,  s_89_15,  s_88_15, 
 s_87_15,  s_86_15,  s_85_15,  s_84_15,  s_83_15,  s_82_15, 
 s_81_15,  s_80_15,  s_79_15,  s_78_15,  s_77_15,  s_76_15, 
 s_75_15,  s_74_15,  s_73_15,  s_72_15,  s_71_15,  s_70_15, 
 s_69_15,  s_68_15,  s_67_15,  s_66_15,  s_65_15,  s_64_15, 
 s_63_15,  s_62_15,  s_61_15,  s_60_15,  s_59_15,  s_58_15, 
 s_57_15,  s_56_15,  s_55_15,  s_54_15,  s_53_15,  s_52_15, 
 s_51_15,  s_50_15,  s_49_15,  s_48_15,  s_47_15,  s_46_15, 
 s_45_15,  s_44_15,  s_43_15,  s_42_15,  s_41_15,  s_40_15, 
 s_39_15,  s_38_15,  s_37_15,  s_36_15,  s_35_15,  s_34_15, 
 s_33_15,  s_32_15,  s_31_15,  s_30_15
} = partial_products[(width+2)*(15+1)-1:(width+2)*15];

assign {
 s_161_0,  s_160_0,  s_159_1,  s_158_1,  s_157_2,  s_156_2, 
 s_155_3,  s_154_3,  s_153_4,  s_152_4,  s_151_5,  s_150_5, 
 s_149_6,  s_148_6,  s_147_7,  s_146_7,  s_145_8,  s_144_8, 
 s_143_9,  s_142_9, s_141_10, s_140_10, s_139_11, s_138_11, 
s_137_12, s_136_12, s_135_13, s_134_13, s_133_14, s_132_14, 
s_131_15, s_130_15, s_129_16, s_128_16, s_127_16, s_126_16, 
s_125_16, s_124_16, s_123_16, s_122_16, s_121_16, s_120_16, 
s_119_16, s_118_16, s_117_16, s_116_16, s_115_16, s_114_16, 
s_113_16, s_112_16, s_111_16, s_110_16, s_109_16, s_108_16, 
s_107_16, s_106_16, s_105_16, s_104_16, s_103_16, s_102_16, 
s_101_16, s_100_16,  s_99_16,  s_98_16,  s_97_16,  s_96_16, 
 s_95_16,  s_94_16,  s_93_16,  s_92_16,  s_91_16,  s_90_16, 
 s_89_16,  s_88_16,  s_87_16,  s_86_16,  s_85_16,  s_84_16, 
 s_83_16,  s_82_16,  s_81_16,  s_80_16,  s_79_16,  s_78_16, 
 s_77_16,  s_76_16,  s_75_16,  s_74_16,  s_73_16,  s_72_16, 
 s_71_16,  s_70_16,  s_69_16,  s_68_16,  s_67_16,  s_66_16, 
 s_65_16,  s_64_16,  s_63_16,  s_62_16,  s_61_16,  s_60_16, 
 s_59_16,  s_58_16,  s_57_16,  s_56_16,  s_55_16,  s_54_16, 
 s_53_16,  s_52_16,  s_51_16,  s_50_16,  s_49_16,  s_48_16, 
 s_47_16,  s_46_16,  s_45_16,  s_44_16,  s_43_16,  s_42_16, 
 s_41_16,  s_40_16,  s_39_16,  s_38_16,  s_37_16,  s_36_16, 
 s_35_16,  s_34_16,  s_33_16,  s_32_16
} = partial_products[(width+2)*(16+1)-1:(width+2)*16];

assign {
 s_163_0,  s_162_0,  s_161_1,  s_160_1,  s_159_2,  s_158_2, 
 s_157_3,  s_156_3,  s_155_4,  s_154_4,  s_153_5,  s_152_5, 
 s_151_6,  s_150_6,  s_149_7,  s_148_7,  s_147_8,  s_146_8, 
 s_145_9,  s_144_9, s_143_10, s_142_10, s_141_11, s_140_11, 
s_139_12, s_138_12, s_137_13, s_136_13, s_135_14, s_134_14, 
s_133_15, s_132_15, s_131_16, s_130_16, s_129_17, s_128_17, 
s_127_17, s_126_17, s_125_17, s_124_17, s_123_17, s_122_17, 
s_121_17, s_120_17, s_119_17, s_118_17, s_117_17, s_116_17, 
s_115_17, s_114_17, s_113_17, s_112_17, s_111_17, s_110_17, 
s_109_17, s_108_17, s_107_17, s_106_17, s_105_17, s_104_17, 
s_103_17, s_102_17, s_101_17, s_100_17,  s_99_17,  s_98_17, 
 s_97_17,  s_96_17,  s_95_17,  s_94_17,  s_93_17,  s_92_17, 
 s_91_17,  s_90_17,  s_89_17,  s_88_17,  s_87_17,  s_86_17, 
 s_85_17,  s_84_17,  s_83_17,  s_82_17,  s_81_17,  s_80_17, 
 s_79_17,  s_78_17,  s_77_17,  s_76_17,  s_75_17,  s_74_17, 
 s_73_17,  s_72_17,  s_71_17,  s_70_17,  s_69_17,  s_68_17, 
 s_67_17,  s_66_17,  s_65_17,  s_64_17,  s_63_17,  s_62_17, 
 s_61_17,  s_60_17,  s_59_17,  s_58_17,  s_57_17,  s_56_17, 
 s_55_17,  s_54_17,  s_53_17,  s_52_17,  s_51_17,  s_50_17, 
 s_49_17,  s_48_17,  s_47_17,  s_46_17,  s_45_17,  s_44_17, 
 s_43_17,  s_42_17,  s_41_17,  s_40_17,  s_39_17,  s_38_17, 
 s_37_17,  s_36_17,  s_35_17,  s_34_17
} = partial_products[(width+2)*(17+1)-1:(width+2)*17];

assign {
 s_165_0,  s_164_0,  s_163_1,  s_162_1,  s_161_2,  s_160_2, 
 s_159_3,  s_158_3,  s_157_4,  s_156_4,  s_155_5,  s_154_5, 
 s_153_6,  s_152_6,  s_151_7,  s_150_7,  s_149_8,  s_148_8, 
 s_147_9,  s_146_9, s_145_10, s_144_10, s_143_11, s_142_11, 
s_141_12, s_140_12, s_139_13, s_138_13, s_137_14, s_136_14, 
s_135_15, s_134_15, s_133_16, s_132_16, s_131_17, s_130_17, 
s_129_18, s_128_18, s_127_18, s_126_18, s_125_18, s_124_18, 
s_123_18, s_122_18, s_121_18, s_120_18, s_119_18, s_118_18, 
s_117_18, s_116_18, s_115_18, s_114_18, s_113_18, s_112_18, 
s_111_18, s_110_18, s_109_18, s_108_18, s_107_18, s_106_18, 
s_105_18, s_104_18, s_103_18, s_102_18, s_101_18, s_100_18, 
 s_99_18,  s_98_18,  s_97_18,  s_96_18,  s_95_18,  s_94_18, 
 s_93_18,  s_92_18,  s_91_18,  s_90_18,  s_89_18,  s_88_18, 
 s_87_18,  s_86_18,  s_85_18,  s_84_18,  s_83_18,  s_82_18, 
 s_81_18,  s_80_18,  s_79_18,  s_78_18,  s_77_18,  s_76_18, 
 s_75_18,  s_74_18,  s_73_18,  s_72_18,  s_71_18,  s_70_18, 
 s_69_18,  s_68_18,  s_67_18,  s_66_18,  s_65_18,  s_64_18, 
 s_63_18,  s_62_18,  s_61_18,  s_60_18,  s_59_18,  s_58_18, 
 s_57_18,  s_56_18,  s_55_18,  s_54_18,  s_53_18,  s_52_18, 
 s_51_18,  s_50_18,  s_49_18,  s_48_18,  s_47_18,  s_46_18, 
 s_45_18,  s_44_18,  s_43_18,  s_42_18,  s_41_18,  s_40_18, 
 s_39_18,  s_38_18,  s_37_18,  s_36_18
} = partial_products[(width+2)*(18+1)-1:(width+2)*18];

assign {
 s_167_0,  s_166_0,  s_165_1,  s_164_1,  s_163_2,  s_162_2, 
 s_161_3,  s_160_3,  s_159_4,  s_158_4,  s_157_5,  s_156_5, 
 s_155_6,  s_154_6,  s_153_7,  s_152_7,  s_151_8,  s_150_8, 
 s_149_9,  s_148_9, s_147_10, s_146_10, s_145_11, s_144_11, 
s_143_12, s_142_12, s_141_13, s_140_13, s_139_14, s_138_14, 
s_137_15, s_136_15, s_135_16, s_134_16, s_133_17, s_132_17, 
s_131_18, s_130_18, s_129_19, s_128_19, s_127_19, s_126_19, 
s_125_19, s_124_19, s_123_19, s_122_19, s_121_19, s_120_19, 
s_119_19, s_118_19, s_117_19, s_116_19, s_115_19, s_114_19, 
s_113_19, s_112_19, s_111_19, s_110_19, s_109_19, s_108_19, 
s_107_19, s_106_19, s_105_19, s_104_19, s_103_19, s_102_19, 
s_101_19, s_100_19,  s_99_19,  s_98_19,  s_97_19,  s_96_19, 
 s_95_19,  s_94_19,  s_93_19,  s_92_19,  s_91_19,  s_90_19, 
 s_89_19,  s_88_19,  s_87_19,  s_86_19,  s_85_19,  s_84_19, 
 s_83_19,  s_82_19,  s_81_19,  s_80_19,  s_79_19,  s_78_19, 
 s_77_19,  s_76_19,  s_75_19,  s_74_19,  s_73_19,  s_72_19, 
 s_71_19,  s_70_19,  s_69_19,  s_68_19,  s_67_19,  s_66_19, 
 s_65_19,  s_64_19,  s_63_19,  s_62_19,  s_61_19,  s_60_19, 
 s_59_19,  s_58_19,  s_57_19,  s_56_19,  s_55_19,  s_54_19, 
 s_53_19,  s_52_19,  s_51_19,  s_50_19,  s_49_19,  s_48_19, 
 s_47_19,  s_46_19,  s_45_19,  s_44_19,  s_43_19,  s_42_19, 
 s_41_19,  s_40_19,  s_39_19,  s_38_19
} = partial_products[(width+2)*(19+1)-1:(width+2)*19];

assign {
 s_169_0,  s_168_0,  s_167_1,  s_166_1,  s_165_2,  s_164_2, 
 s_163_3,  s_162_3,  s_161_4,  s_160_4,  s_159_5,  s_158_5, 
 s_157_6,  s_156_6,  s_155_7,  s_154_7,  s_153_8,  s_152_8, 
 s_151_9,  s_150_9, s_149_10, s_148_10, s_147_11, s_146_11, 
s_145_12, s_144_12, s_143_13, s_142_13, s_141_14, s_140_14, 
s_139_15, s_138_15, s_137_16, s_136_16, s_135_17, s_134_17, 
s_133_18, s_132_18, s_131_19, s_130_19, s_129_20, s_128_20, 
s_127_20, s_126_20, s_125_20, s_124_20, s_123_20, s_122_20, 
s_121_20, s_120_20, s_119_20, s_118_20, s_117_20, s_116_20, 
s_115_20, s_114_20, s_113_20, s_112_20, s_111_20, s_110_20, 
s_109_20, s_108_20, s_107_20, s_106_20, s_105_20, s_104_20, 
s_103_20, s_102_20, s_101_20, s_100_20,  s_99_20,  s_98_20, 
 s_97_20,  s_96_20,  s_95_20,  s_94_20,  s_93_20,  s_92_20, 
 s_91_20,  s_90_20,  s_89_20,  s_88_20,  s_87_20,  s_86_20, 
 s_85_20,  s_84_20,  s_83_20,  s_82_20,  s_81_20,  s_80_20, 
 s_79_20,  s_78_20,  s_77_20,  s_76_20,  s_75_20,  s_74_20, 
 s_73_20,  s_72_20,  s_71_20,  s_70_20,  s_69_20,  s_68_20, 
 s_67_20,  s_66_20,  s_65_20,  s_64_20,  s_63_20,  s_62_20, 
 s_61_20,  s_60_20,  s_59_20,  s_58_20,  s_57_20,  s_56_20, 
 s_55_20,  s_54_20,  s_53_20,  s_52_20,  s_51_20,  s_50_20, 
 s_49_20,  s_48_20,  s_47_20,  s_46_20,  s_45_20,  s_44_20, 
 s_43_20,  s_42_20,  s_41_20,  s_40_20
} = partial_products[(width+2)*(20+1)-1:(width+2)*20];

assign {
 s_171_0,  s_170_0,  s_169_1,  s_168_1,  s_167_2,  s_166_2, 
 s_165_3,  s_164_3,  s_163_4,  s_162_4,  s_161_5,  s_160_5, 
 s_159_6,  s_158_6,  s_157_7,  s_156_7,  s_155_8,  s_154_8, 
 s_153_9,  s_152_9, s_151_10, s_150_10, s_149_11, s_148_11, 
s_147_12, s_146_12, s_145_13, s_144_13, s_143_14, s_142_14, 
s_141_15, s_140_15, s_139_16, s_138_16, s_137_17, s_136_17, 
s_135_18, s_134_18, s_133_19, s_132_19, s_131_20, s_130_20, 
s_129_21, s_128_21, s_127_21, s_126_21, s_125_21, s_124_21, 
s_123_21, s_122_21, s_121_21, s_120_21, s_119_21, s_118_21, 
s_117_21, s_116_21, s_115_21, s_114_21, s_113_21, s_112_21, 
s_111_21, s_110_21, s_109_21, s_108_21, s_107_21, s_106_21, 
s_105_21, s_104_21, s_103_21, s_102_21, s_101_21, s_100_21, 
 s_99_21,  s_98_21,  s_97_21,  s_96_21,  s_95_21,  s_94_21, 
 s_93_21,  s_92_21,  s_91_21,  s_90_21,  s_89_21,  s_88_21, 
 s_87_21,  s_86_21,  s_85_21,  s_84_21,  s_83_21,  s_82_21, 
 s_81_21,  s_80_21,  s_79_21,  s_78_21,  s_77_21,  s_76_21, 
 s_75_21,  s_74_21,  s_73_21,  s_72_21,  s_71_21,  s_70_21, 
 s_69_21,  s_68_21,  s_67_21,  s_66_21,  s_65_21,  s_64_21, 
 s_63_21,  s_62_21,  s_61_21,  s_60_21,  s_59_21,  s_58_21, 
 s_57_21,  s_56_21,  s_55_21,  s_54_21,  s_53_21,  s_52_21, 
 s_51_21,  s_50_21,  s_49_21,  s_48_21,  s_47_21,  s_46_21, 
 s_45_21,  s_44_21,  s_43_21,  s_42_21
} = partial_products[(width+2)*(21+1)-1:(width+2)*21];

assign {
 s_173_0,  s_172_0,  s_171_1,  s_170_1,  s_169_2,  s_168_2, 
 s_167_3,  s_166_3,  s_165_4,  s_164_4,  s_163_5,  s_162_5, 
 s_161_6,  s_160_6,  s_159_7,  s_158_7,  s_157_8,  s_156_8, 
 s_155_9,  s_154_9, s_153_10, s_152_10, s_151_11, s_150_11, 
s_149_12, s_148_12, s_147_13, s_146_13, s_145_14, s_144_14, 
s_143_15, s_142_15, s_141_16, s_140_16, s_139_17, s_138_17, 
s_137_18, s_136_18, s_135_19, s_134_19, s_133_20, s_132_20, 
s_131_21, s_130_21, s_129_22, s_128_22, s_127_22, s_126_22, 
s_125_22, s_124_22, s_123_22, s_122_22, s_121_22, s_120_22, 
s_119_22, s_118_22, s_117_22, s_116_22, s_115_22, s_114_22, 
s_113_22, s_112_22, s_111_22, s_110_22, s_109_22, s_108_22, 
s_107_22, s_106_22, s_105_22, s_104_22, s_103_22, s_102_22, 
s_101_22, s_100_22,  s_99_22,  s_98_22,  s_97_22,  s_96_22, 
 s_95_22,  s_94_22,  s_93_22,  s_92_22,  s_91_22,  s_90_22, 
 s_89_22,  s_88_22,  s_87_22,  s_86_22,  s_85_22,  s_84_22, 
 s_83_22,  s_82_22,  s_81_22,  s_80_22,  s_79_22,  s_78_22, 
 s_77_22,  s_76_22,  s_75_22,  s_74_22,  s_73_22,  s_72_22, 
 s_71_22,  s_70_22,  s_69_22,  s_68_22,  s_67_22,  s_66_22, 
 s_65_22,  s_64_22,  s_63_22,  s_62_22,  s_61_22,  s_60_22, 
 s_59_22,  s_58_22,  s_57_22,  s_56_22,  s_55_22,  s_54_22, 
 s_53_22,  s_52_22,  s_51_22,  s_50_22,  s_49_22,  s_48_22, 
 s_47_22,  s_46_22,  s_45_22,  s_44_22
} = partial_products[(width+2)*(22+1)-1:(width+2)*22];

assign {
 s_175_0,  s_174_0,  s_173_1,  s_172_1,  s_171_2,  s_170_2, 
 s_169_3,  s_168_3,  s_167_4,  s_166_4,  s_165_5,  s_164_5, 
 s_163_6,  s_162_6,  s_161_7,  s_160_7,  s_159_8,  s_158_8, 
 s_157_9,  s_156_9, s_155_10, s_154_10, s_153_11, s_152_11, 
s_151_12, s_150_12, s_149_13, s_148_13, s_147_14, s_146_14, 
s_145_15, s_144_15, s_143_16, s_142_16, s_141_17, s_140_17, 
s_139_18, s_138_18, s_137_19, s_136_19, s_135_20, s_134_20, 
s_133_21, s_132_21, s_131_22, s_130_22, s_129_23, s_128_23, 
s_127_23, s_126_23, s_125_23, s_124_23, s_123_23, s_122_23, 
s_121_23, s_120_23, s_119_23, s_118_23, s_117_23, s_116_23, 
s_115_23, s_114_23, s_113_23, s_112_23, s_111_23, s_110_23, 
s_109_23, s_108_23, s_107_23, s_106_23, s_105_23, s_104_23, 
s_103_23, s_102_23, s_101_23, s_100_23,  s_99_23,  s_98_23, 
 s_97_23,  s_96_23,  s_95_23,  s_94_23,  s_93_23,  s_92_23, 
 s_91_23,  s_90_23,  s_89_23,  s_88_23,  s_87_23,  s_86_23, 
 s_85_23,  s_84_23,  s_83_23,  s_82_23,  s_81_23,  s_80_23, 
 s_79_23,  s_78_23,  s_77_23,  s_76_23,  s_75_23,  s_74_23, 
 s_73_23,  s_72_23,  s_71_23,  s_70_23,  s_69_23,  s_68_23, 
 s_67_23,  s_66_23,  s_65_23,  s_64_23,  s_63_23,  s_62_23, 
 s_61_23,  s_60_23,  s_59_23,  s_58_23,  s_57_23,  s_56_23, 
 s_55_23,  s_54_23,  s_53_23,  s_52_23,  s_51_23,  s_50_23, 
 s_49_23,  s_48_23,  s_47_23,  s_46_23
} = partial_products[(width+2)*(23+1)-1:(width+2)*23];

assign {
 s_177_0,  s_176_0,  s_175_1,  s_174_1,  s_173_2,  s_172_2, 
 s_171_3,  s_170_3,  s_169_4,  s_168_4,  s_167_5,  s_166_5, 
 s_165_6,  s_164_6,  s_163_7,  s_162_7,  s_161_8,  s_160_8, 
 s_159_9,  s_158_9, s_157_10, s_156_10, s_155_11, s_154_11, 
s_153_12, s_152_12, s_151_13, s_150_13, s_149_14, s_148_14, 
s_147_15, s_146_15, s_145_16, s_144_16, s_143_17, s_142_17, 
s_141_18, s_140_18, s_139_19, s_138_19, s_137_20, s_136_20, 
s_135_21, s_134_21, s_133_22, s_132_22, s_131_23, s_130_23, 
s_129_24, s_128_24, s_127_24, s_126_24, s_125_24, s_124_24, 
s_123_24, s_122_24, s_121_24, s_120_24, s_119_24, s_118_24, 
s_117_24, s_116_24, s_115_24, s_114_24, s_113_24, s_112_24, 
s_111_24, s_110_24, s_109_24, s_108_24, s_107_24, s_106_24, 
s_105_24, s_104_24, s_103_24, s_102_24, s_101_24, s_100_24, 
 s_99_24,  s_98_24,  s_97_24,  s_96_24,  s_95_24,  s_94_24, 
 s_93_24,  s_92_24,  s_91_24,  s_90_24,  s_89_24,  s_88_24, 
 s_87_24,  s_86_24,  s_85_24,  s_84_24,  s_83_24,  s_82_24, 
 s_81_24,  s_80_24,  s_79_24,  s_78_24,  s_77_24,  s_76_24, 
 s_75_24,  s_74_24,  s_73_24,  s_72_24,  s_71_24,  s_70_24, 
 s_69_24,  s_68_24,  s_67_24,  s_66_24,  s_65_24,  s_64_24, 
 s_63_24,  s_62_24,  s_61_24,  s_60_24,  s_59_24,  s_58_24, 
 s_57_24,  s_56_24,  s_55_24,  s_54_24,  s_53_24,  s_52_24, 
 s_51_24,  s_50_24,  s_49_24,  s_48_24
} = partial_products[(width+2)*(24+1)-1:(width+2)*24];

assign {
 s_179_0,  s_178_0,  s_177_1,  s_176_1,  s_175_2,  s_174_2, 
 s_173_3,  s_172_3,  s_171_4,  s_170_4,  s_169_5,  s_168_5, 
 s_167_6,  s_166_6,  s_165_7,  s_164_7,  s_163_8,  s_162_8, 
 s_161_9,  s_160_9, s_159_10, s_158_10, s_157_11, s_156_11, 
s_155_12, s_154_12, s_153_13, s_152_13, s_151_14, s_150_14, 
s_149_15, s_148_15, s_147_16, s_146_16, s_145_17, s_144_17, 
s_143_18, s_142_18, s_141_19, s_140_19, s_139_20, s_138_20, 
s_137_21, s_136_21, s_135_22, s_134_22, s_133_23, s_132_23, 
s_131_24, s_130_24, s_129_25, s_128_25, s_127_25, s_126_25, 
s_125_25, s_124_25, s_123_25, s_122_25, s_121_25, s_120_25, 
s_119_25, s_118_25, s_117_25, s_116_25, s_115_25, s_114_25, 
s_113_25, s_112_25, s_111_25, s_110_25, s_109_25, s_108_25, 
s_107_25, s_106_25, s_105_25, s_104_25, s_103_25, s_102_25, 
s_101_25, s_100_25,  s_99_25,  s_98_25,  s_97_25,  s_96_25, 
 s_95_25,  s_94_25,  s_93_25,  s_92_25,  s_91_25,  s_90_25, 
 s_89_25,  s_88_25,  s_87_25,  s_86_25,  s_85_25,  s_84_25, 
 s_83_25,  s_82_25,  s_81_25,  s_80_25,  s_79_25,  s_78_25, 
 s_77_25,  s_76_25,  s_75_25,  s_74_25,  s_73_25,  s_72_25, 
 s_71_25,  s_70_25,  s_69_25,  s_68_25,  s_67_25,  s_66_25, 
 s_65_25,  s_64_25,  s_63_25,  s_62_25,  s_61_25,  s_60_25, 
 s_59_25,  s_58_25,  s_57_25,  s_56_25,  s_55_25,  s_54_25, 
 s_53_25,  s_52_25,  s_51_25,  s_50_25
} = partial_products[(width+2)*(25+1)-1:(width+2)*25];

assign {
 s_181_0,  s_180_0,  s_179_1,  s_178_1,  s_177_2,  s_176_2, 
 s_175_3,  s_174_3,  s_173_4,  s_172_4,  s_171_5,  s_170_5, 
 s_169_6,  s_168_6,  s_167_7,  s_166_7,  s_165_8,  s_164_8, 
 s_163_9,  s_162_9, s_161_10, s_160_10, s_159_11, s_158_11, 
s_157_12, s_156_12, s_155_13, s_154_13, s_153_14, s_152_14, 
s_151_15, s_150_15, s_149_16, s_148_16, s_147_17, s_146_17, 
s_145_18, s_144_18, s_143_19, s_142_19, s_141_20, s_140_20, 
s_139_21, s_138_21, s_137_22, s_136_22, s_135_23, s_134_23, 
s_133_24, s_132_24, s_131_25, s_130_25, s_129_26, s_128_26, 
s_127_26, s_126_26, s_125_26, s_124_26, s_123_26, s_122_26, 
s_121_26, s_120_26, s_119_26, s_118_26, s_117_26, s_116_26, 
s_115_26, s_114_26, s_113_26, s_112_26, s_111_26, s_110_26, 
s_109_26, s_108_26, s_107_26, s_106_26, s_105_26, s_104_26, 
s_103_26, s_102_26, s_101_26, s_100_26,  s_99_26,  s_98_26, 
 s_97_26,  s_96_26,  s_95_26,  s_94_26,  s_93_26,  s_92_26, 
 s_91_26,  s_90_26,  s_89_26,  s_88_26,  s_87_26,  s_86_26, 
 s_85_26,  s_84_26,  s_83_26,  s_82_26,  s_81_26,  s_80_26, 
 s_79_26,  s_78_26,  s_77_26,  s_76_26,  s_75_26,  s_74_26, 
 s_73_26,  s_72_26,  s_71_26,  s_70_26,  s_69_26,  s_68_26, 
 s_67_26,  s_66_26,  s_65_26,  s_64_26,  s_63_26,  s_62_26, 
 s_61_26,  s_60_26,  s_59_26,  s_58_26,  s_57_26,  s_56_26, 
 s_55_26,  s_54_26,  s_53_26,  s_52_26
} = partial_products[(width+2)*(26+1)-1:(width+2)*26];

assign {
 s_183_0,  s_182_0,  s_181_1,  s_180_1,  s_179_2,  s_178_2, 
 s_177_3,  s_176_3,  s_175_4,  s_174_4,  s_173_5,  s_172_5, 
 s_171_6,  s_170_6,  s_169_7,  s_168_7,  s_167_8,  s_166_8, 
 s_165_9,  s_164_9, s_163_10, s_162_10, s_161_11, s_160_11, 
s_159_12, s_158_12, s_157_13, s_156_13, s_155_14, s_154_14, 
s_153_15, s_152_15, s_151_16, s_150_16, s_149_17, s_148_17, 
s_147_18, s_146_18, s_145_19, s_144_19, s_143_20, s_142_20, 
s_141_21, s_140_21, s_139_22, s_138_22, s_137_23, s_136_23, 
s_135_24, s_134_24, s_133_25, s_132_25, s_131_26, s_130_26, 
s_129_27, s_128_27, s_127_27, s_126_27, s_125_27, s_124_27, 
s_123_27, s_122_27, s_121_27, s_120_27, s_119_27, s_118_27, 
s_117_27, s_116_27, s_115_27, s_114_27, s_113_27, s_112_27, 
s_111_27, s_110_27, s_109_27, s_108_27, s_107_27, s_106_27, 
s_105_27, s_104_27, s_103_27, s_102_27, s_101_27, s_100_27, 
 s_99_27,  s_98_27,  s_97_27,  s_96_27,  s_95_27,  s_94_27, 
 s_93_27,  s_92_27,  s_91_27,  s_90_27,  s_89_27,  s_88_27, 
 s_87_27,  s_86_27,  s_85_27,  s_84_27,  s_83_27,  s_82_27, 
 s_81_27,  s_80_27,  s_79_27,  s_78_27,  s_77_27,  s_76_27, 
 s_75_27,  s_74_27,  s_73_27,  s_72_27,  s_71_27,  s_70_27, 
 s_69_27,  s_68_27,  s_67_27,  s_66_27,  s_65_27,  s_64_27, 
 s_63_27,  s_62_27,  s_61_27,  s_60_27,  s_59_27,  s_58_27, 
 s_57_27,  s_56_27,  s_55_27,  s_54_27
} = partial_products[(width+2)*(27+1)-1:(width+2)*27];

assign {
 s_185_0,  s_184_0,  s_183_1,  s_182_1,  s_181_2,  s_180_2, 
 s_179_3,  s_178_3,  s_177_4,  s_176_4,  s_175_5,  s_174_5, 
 s_173_6,  s_172_6,  s_171_7,  s_170_7,  s_169_8,  s_168_8, 
 s_167_9,  s_166_9, s_165_10, s_164_10, s_163_11, s_162_11, 
s_161_12, s_160_12, s_159_13, s_158_13, s_157_14, s_156_14, 
s_155_15, s_154_15, s_153_16, s_152_16, s_151_17, s_150_17, 
s_149_18, s_148_18, s_147_19, s_146_19, s_145_20, s_144_20, 
s_143_21, s_142_21, s_141_22, s_140_22, s_139_23, s_138_23, 
s_137_24, s_136_24, s_135_25, s_134_25, s_133_26, s_132_26, 
s_131_27, s_130_27, s_129_28, s_128_28, s_127_28, s_126_28, 
s_125_28, s_124_28, s_123_28, s_122_28, s_121_28, s_120_28, 
s_119_28, s_118_28, s_117_28, s_116_28, s_115_28, s_114_28, 
s_113_28, s_112_28, s_111_28, s_110_28, s_109_28, s_108_28, 
s_107_28, s_106_28, s_105_28, s_104_28, s_103_28, s_102_28, 
s_101_28, s_100_28,  s_99_28,  s_98_28,  s_97_28,  s_96_28, 
 s_95_28,  s_94_28,  s_93_28,  s_92_28,  s_91_28,  s_90_28, 
 s_89_28,  s_88_28,  s_87_28,  s_86_28,  s_85_28,  s_84_28, 
 s_83_28,  s_82_28,  s_81_28,  s_80_28,  s_79_28,  s_78_28, 
 s_77_28,  s_76_28,  s_75_28,  s_74_28,  s_73_28,  s_72_28, 
 s_71_28,  s_70_28,  s_69_28,  s_68_28,  s_67_28,  s_66_28, 
 s_65_28,  s_64_28,  s_63_28,  s_62_28,  s_61_28,  s_60_28, 
 s_59_28,  s_58_28,  s_57_28,  s_56_28
} = partial_products[(width+2)*(28+1)-1:(width+2)*28];

assign {
 s_187_0,  s_186_0,  s_185_1,  s_184_1,  s_183_2,  s_182_2, 
 s_181_3,  s_180_3,  s_179_4,  s_178_4,  s_177_5,  s_176_5, 
 s_175_6,  s_174_6,  s_173_7,  s_172_7,  s_171_8,  s_170_8, 
 s_169_9,  s_168_9, s_167_10, s_166_10, s_165_11, s_164_11, 
s_163_12, s_162_12, s_161_13, s_160_13, s_159_14, s_158_14, 
s_157_15, s_156_15, s_155_16, s_154_16, s_153_17, s_152_17, 
s_151_18, s_150_18, s_149_19, s_148_19, s_147_20, s_146_20, 
s_145_21, s_144_21, s_143_22, s_142_22, s_141_23, s_140_23, 
s_139_24, s_138_24, s_137_25, s_136_25, s_135_26, s_134_26, 
s_133_27, s_132_27, s_131_28, s_130_28, s_129_29, s_128_29, 
s_127_29, s_126_29, s_125_29, s_124_29, s_123_29, s_122_29, 
s_121_29, s_120_29, s_119_29, s_118_29, s_117_29, s_116_29, 
s_115_29, s_114_29, s_113_29, s_112_29, s_111_29, s_110_29, 
s_109_29, s_108_29, s_107_29, s_106_29, s_105_29, s_104_29, 
s_103_29, s_102_29, s_101_29, s_100_29,  s_99_29,  s_98_29, 
 s_97_29,  s_96_29,  s_95_29,  s_94_29,  s_93_29,  s_92_29, 
 s_91_29,  s_90_29,  s_89_29,  s_88_29,  s_87_29,  s_86_29, 
 s_85_29,  s_84_29,  s_83_29,  s_82_29,  s_81_29,  s_80_29, 
 s_79_29,  s_78_29,  s_77_29,  s_76_29,  s_75_29,  s_74_29, 
 s_73_29,  s_72_29,  s_71_29,  s_70_29,  s_69_29,  s_68_29, 
 s_67_29,  s_66_29,  s_65_29,  s_64_29,  s_63_29,  s_62_29, 
 s_61_29,  s_60_29,  s_59_29,  s_58_29
} = partial_products[(width+2)*(29+1)-1:(width+2)*29];

assign {
 s_189_0,  s_188_0,  s_187_1,  s_186_1,  s_185_2,  s_184_2, 
 s_183_3,  s_182_3,  s_181_4,  s_180_4,  s_179_5,  s_178_5, 
 s_177_6,  s_176_6,  s_175_7,  s_174_7,  s_173_8,  s_172_8, 
 s_171_9,  s_170_9, s_169_10, s_168_10, s_167_11, s_166_11, 
s_165_12, s_164_12, s_163_13, s_162_13, s_161_14, s_160_14, 
s_159_15, s_158_15, s_157_16, s_156_16, s_155_17, s_154_17, 
s_153_18, s_152_18, s_151_19, s_150_19, s_149_20, s_148_20, 
s_147_21, s_146_21, s_145_22, s_144_22, s_143_23, s_142_23, 
s_141_24, s_140_24, s_139_25, s_138_25, s_137_26, s_136_26, 
s_135_27, s_134_27, s_133_28, s_132_28, s_131_29, s_130_29, 
s_129_30, s_128_30, s_127_30, s_126_30, s_125_30, s_124_30, 
s_123_30, s_122_30, s_121_30, s_120_30, s_119_30, s_118_30, 
s_117_30, s_116_30, s_115_30, s_114_30, s_113_30, s_112_30, 
s_111_30, s_110_30, s_109_30, s_108_30, s_107_30, s_106_30, 
s_105_30, s_104_30, s_103_30, s_102_30, s_101_30, s_100_30, 
 s_99_30,  s_98_30,  s_97_30,  s_96_30,  s_95_30,  s_94_30, 
 s_93_30,  s_92_30,  s_91_30,  s_90_30,  s_89_30,  s_88_30, 
 s_87_30,  s_86_30,  s_85_30,  s_84_30,  s_83_30,  s_82_30, 
 s_81_30,  s_80_30,  s_79_30,  s_78_30,  s_77_30,  s_76_30, 
 s_75_30,  s_74_30,  s_73_30,  s_72_30,  s_71_30,  s_70_30, 
 s_69_30,  s_68_30,  s_67_30,  s_66_30,  s_65_30,  s_64_30, 
 s_63_30,  s_62_30,  s_61_30,  s_60_30
} = partial_products[(width+2)*(30+1)-1:(width+2)*30];

assign {
 s_191_0,  s_190_0,  s_189_1,  s_188_1,  s_187_2,  s_186_2, 
 s_185_3,  s_184_3,  s_183_4,  s_182_4,  s_181_5,  s_180_5, 
 s_179_6,  s_178_6,  s_177_7,  s_176_7,  s_175_8,  s_174_8, 
 s_173_9,  s_172_9, s_171_10, s_170_10, s_169_11, s_168_11, 
s_167_12, s_166_12, s_165_13, s_164_13, s_163_14, s_162_14, 
s_161_15, s_160_15, s_159_16, s_158_16, s_157_17, s_156_17, 
s_155_18, s_154_18, s_153_19, s_152_19, s_151_20, s_150_20, 
s_149_21, s_148_21, s_147_22, s_146_22, s_145_23, s_144_23, 
s_143_24, s_142_24, s_141_25, s_140_25, s_139_26, s_138_26, 
s_137_27, s_136_27, s_135_28, s_134_28, s_133_29, s_132_29, 
s_131_30, s_130_30, s_129_31, s_128_31, s_127_31, s_126_31, 
s_125_31, s_124_31, s_123_31, s_122_31, s_121_31, s_120_31, 
s_119_31, s_118_31, s_117_31, s_116_31, s_115_31, s_114_31, 
s_113_31, s_112_31, s_111_31, s_110_31, s_109_31, s_108_31, 
s_107_31, s_106_31, s_105_31, s_104_31, s_103_31, s_102_31, 
s_101_31, s_100_31,  s_99_31,  s_98_31,  s_97_31,  s_96_31, 
 s_95_31,  s_94_31,  s_93_31,  s_92_31,  s_91_31,  s_90_31, 
 s_89_31,  s_88_31,  s_87_31,  s_86_31,  s_85_31,  s_84_31, 
 s_83_31,  s_82_31,  s_81_31,  s_80_31,  s_79_31,  s_78_31, 
 s_77_31,  s_76_31,  s_75_31,  s_74_31,  s_73_31,  s_72_31, 
 s_71_31,  s_70_31,  s_69_31,  s_68_31,  s_67_31,  s_66_31, 
 s_65_31,  s_64_31,  s_63_31,  s_62_31
} = partial_products[(width+2)*(31+1)-1:(width+2)*31];

assign {
 s_193_0,  s_192_0,  s_191_1,  s_190_1,  s_189_2,  s_188_2, 
 s_187_3,  s_186_3,  s_185_4,  s_184_4,  s_183_5,  s_182_5, 
 s_181_6,  s_180_6,  s_179_7,  s_178_7,  s_177_8,  s_176_8, 
 s_175_9,  s_174_9, s_173_10, s_172_10, s_171_11, s_170_11, 
s_169_12, s_168_12, s_167_13, s_166_13, s_165_14, s_164_14, 
s_163_15, s_162_15, s_161_16, s_160_16, s_159_17, s_158_17, 
s_157_18, s_156_18, s_155_19, s_154_19, s_153_20, s_152_20, 
s_151_21, s_150_21, s_149_22, s_148_22, s_147_23, s_146_23, 
s_145_24, s_144_24, s_143_25, s_142_25, s_141_26, s_140_26, 
s_139_27, s_138_27, s_137_28, s_136_28, s_135_29, s_134_29, 
s_133_30, s_132_30, s_131_31, s_130_31, s_129_32, s_128_32, 
s_127_32, s_126_32, s_125_32, s_124_32, s_123_32, s_122_32, 
s_121_32, s_120_32, s_119_32, s_118_32, s_117_32, s_116_32, 
s_115_32, s_114_32, s_113_32, s_112_32, s_111_32, s_110_32, 
s_109_32, s_108_32, s_107_32, s_106_32, s_105_32, s_104_32, 
s_103_32, s_102_32, s_101_32, s_100_32,  s_99_32,  s_98_32, 
 s_97_32,  s_96_32,  s_95_32,  s_94_32,  s_93_32,  s_92_32, 
 s_91_32,  s_90_32,  s_89_32,  s_88_32,  s_87_32,  s_86_32, 
 s_85_32,  s_84_32,  s_83_32,  s_82_32,  s_81_32,  s_80_32, 
 s_79_32,  s_78_32,  s_77_32,  s_76_32,  s_75_32,  s_74_32, 
 s_73_32,  s_72_32,  s_71_32,  s_70_32,  s_69_32,  s_68_32, 
 s_67_32,  s_66_32,  s_65_32,  s_64_32
} = partial_products[(width+2)*(32+1)-1:(width+2)*32];

assign {
 s_195_0,  s_194_0,  s_193_1,  s_192_1,  s_191_2,  s_190_2, 
 s_189_3,  s_188_3,  s_187_4,  s_186_4,  s_185_5,  s_184_5, 
 s_183_6,  s_182_6,  s_181_7,  s_180_7,  s_179_8,  s_178_8, 
 s_177_9,  s_176_9, s_175_10, s_174_10, s_173_11, s_172_11, 
s_171_12, s_170_12, s_169_13, s_168_13, s_167_14, s_166_14, 
s_165_15, s_164_15, s_163_16, s_162_16, s_161_17, s_160_17, 
s_159_18, s_158_18, s_157_19, s_156_19, s_155_20, s_154_20, 
s_153_21, s_152_21, s_151_22, s_150_22, s_149_23, s_148_23, 
s_147_24, s_146_24, s_145_25, s_144_25, s_143_26, s_142_26, 
s_141_27, s_140_27, s_139_28, s_138_28, s_137_29, s_136_29, 
s_135_30, s_134_30, s_133_31, s_132_31, s_131_32, s_130_32, 
s_129_33, s_128_33, s_127_33, s_126_33, s_125_33, s_124_33, 
s_123_33, s_122_33, s_121_33, s_120_33, s_119_33, s_118_33, 
s_117_33, s_116_33, s_115_33, s_114_33, s_113_33, s_112_33, 
s_111_33, s_110_33, s_109_33, s_108_33, s_107_33, s_106_33, 
s_105_33, s_104_33, s_103_33, s_102_33, s_101_33, s_100_33, 
 s_99_33,  s_98_33,  s_97_33,  s_96_33,  s_95_33,  s_94_33, 
 s_93_33,  s_92_33,  s_91_33,  s_90_33,  s_89_33,  s_88_33, 
 s_87_33,  s_86_33,  s_85_33,  s_84_33,  s_83_33,  s_82_33, 
 s_81_33,  s_80_33,  s_79_33,  s_78_33,  s_77_33,  s_76_33, 
 s_75_33,  s_74_33,  s_73_33,  s_72_33,  s_71_33,  s_70_33, 
 s_69_33,  s_68_33,  s_67_33,  s_66_33
} = partial_products[(width+2)*(33+1)-1:(width+2)*33];

assign {
 s_197_0,  s_196_0,  s_195_1,  s_194_1,  s_193_2,  s_192_2, 
 s_191_3,  s_190_3,  s_189_4,  s_188_4,  s_187_5,  s_186_5, 
 s_185_6,  s_184_6,  s_183_7,  s_182_7,  s_181_8,  s_180_8, 
 s_179_9,  s_178_9, s_177_10, s_176_10, s_175_11, s_174_11, 
s_173_12, s_172_12, s_171_13, s_170_13, s_169_14, s_168_14, 
s_167_15, s_166_15, s_165_16, s_164_16, s_163_17, s_162_17, 
s_161_18, s_160_18, s_159_19, s_158_19, s_157_20, s_156_20, 
s_155_21, s_154_21, s_153_22, s_152_22, s_151_23, s_150_23, 
s_149_24, s_148_24, s_147_25, s_146_25, s_145_26, s_144_26, 
s_143_27, s_142_27, s_141_28, s_140_28, s_139_29, s_138_29, 
s_137_30, s_136_30, s_135_31, s_134_31, s_133_32, s_132_32, 
s_131_33, s_130_33, s_129_34, s_128_34, s_127_34, s_126_34, 
s_125_34, s_124_34, s_123_34, s_122_34, s_121_34, s_120_34, 
s_119_34, s_118_34, s_117_34, s_116_34, s_115_34, s_114_34, 
s_113_34, s_112_34, s_111_34, s_110_34, s_109_34, s_108_34, 
s_107_34, s_106_34, s_105_34, s_104_34, s_103_34, s_102_34, 
s_101_34, s_100_34,  s_99_34,  s_98_34,  s_97_34,  s_96_34, 
 s_95_34,  s_94_34,  s_93_34,  s_92_34,  s_91_34,  s_90_34, 
 s_89_34,  s_88_34,  s_87_34,  s_86_34,  s_85_34,  s_84_34, 
 s_83_34,  s_82_34,  s_81_34,  s_80_34,  s_79_34,  s_78_34, 
 s_77_34,  s_76_34,  s_75_34,  s_74_34,  s_73_34,  s_72_34, 
 s_71_34,  s_70_34,  s_69_34,  s_68_34
} = partial_products[(width+2)*(34+1)-1:(width+2)*34];

assign {
 s_199_0,  s_198_0,  s_197_1,  s_196_1,  s_195_2,  s_194_2, 
 s_193_3,  s_192_3,  s_191_4,  s_190_4,  s_189_5,  s_188_5, 
 s_187_6,  s_186_6,  s_185_7,  s_184_7,  s_183_8,  s_182_8, 
 s_181_9,  s_180_9, s_179_10, s_178_10, s_177_11, s_176_11, 
s_175_12, s_174_12, s_173_13, s_172_13, s_171_14, s_170_14, 
s_169_15, s_168_15, s_167_16, s_166_16, s_165_17, s_164_17, 
s_163_18, s_162_18, s_161_19, s_160_19, s_159_20, s_158_20, 
s_157_21, s_156_21, s_155_22, s_154_22, s_153_23, s_152_23, 
s_151_24, s_150_24, s_149_25, s_148_25, s_147_26, s_146_26, 
s_145_27, s_144_27, s_143_28, s_142_28, s_141_29, s_140_29, 
s_139_30, s_138_30, s_137_31, s_136_31, s_135_32, s_134_32, 
s_133_33, s_132_33, s_131_34, s_130_34, s_129_35, s_128_35, 
s_127_35, s_126_35, s_125_35, s_124_35, s_123_35, s_122_35, 
s_121_35, s_120_35, s_119_35, s_118_35, s_117_35, s_116_35, 
s_115_35, s_114_35, s_113_35, s_112_35, s_111_35, s_110_35, 
s_109_35, s_108_35, s_107_35, s_106_35, s_105_35, s_104_35, 
s_103_35, s_102_35, s_101_35, s_100_35,  s_99_35,  s_98_35, 
 s_97_35,  s_96_35,  s_95_35,  s_94_35,  s_93_35,  s_92_35, 
 s_91_35,  s_90_35,  s_89_35,  s_88_35,  s_87_35,  s_86_35, 
 s_85_35,  s_84_35,  s_83_35,  s_82_35,  s_81_35,  s_80_35, 
 s_79_35,  s_78_35,  s_77_35,  s_76_35,  s_75_35,  s_74_35, 
 s_73_35,  s_72_35,  s_71_35,  s_70_35
} = partial_products[(width+2)*(35+1)-1:(width+2)*35];

assign {
 s_201_0,  s_200_0,  s_199_1,  s_198_1,  s_197_2,  s_196_2, 
 s_195_3,  s_194_3,  s_193_4,  s_192_4,  s_191_5,  s_190_5, 
 s_189_6,  s_188_6,  s_187_7,  s_186_7,  s_185_8,  s_184_8, 
 s_183_9,  s_182_9, s_181_10, s_180_10, s_179_11, s_178_11, 
s_177_12, s_176_12, s_175_13, s_174_13, s_173_14, s_172_14, 
s_171_15, s_170_15, s_169_16, s_168_16, s_167_17, s_166_17, 
s_165_18, s_164_18, s_163_19, s_162_19, s_161_20, s_160_20, 
s_159_21, s_158_21, s_157_22, s_156_22, s_155_23, s_154_23, 
s_153_24, s_152_24, s_151_25, s_150_25, s_149_26, s_148_26, 
s_147_27, s_146_27, s_145_28, s_144_28, s_143_29, s_142_29, 
s_141_30, s_140_30, s_139_31, s_138_31, s_137_32, s_136_32, 
s_135_33, s_134_33, s_133_34, s_132_34, s_131_35, s_130_35, 
s_129_36, s_128_36, s_127_36, s_126_36, s_125_36, s_124_36, 
s_123_36, s_122_36, s_121_36, s_120_36, s_119_36, s_118_36, 
s_117_36, s_116_36, s_115_36, s_114_36, s_113_36, s_112_36, 
s_111_36, s_110_36, s_109_36, s_108_36, s_107_36, s_106_36, 
s_105_36, s_104_36, s_103_36, s_102_36, s_101_36, s_100_36, 
 s_99_36,  s_98_36,  s_97_36,  s_96_36,  s_95_36,  s_94_36, 
 s_93_36,  s_92_36,  s_91_36,  s_90_36,  s_89_36,  s_88_36, 
 s_87_36,  s_86_36,  s_85_36,  s_84_36,  s_83_36,  s_82_36, 
 s_81_36,  s_80_36,  s_79_36,  s_78_36,  s_77_36,  s_76_36, 
 s_75_36,  s_74_36,  s_73_36,  s_72_36
} = partial_products[(width+2)*(36+1)-1:(width+2)*36];

assign {
 s_203_0,  s_202_0,  s_201_1,  s_200_1,  s_199_2,  s_198_2, 
 s_197_3,  s_196_3,  s_195_4,  s_194_4,  s_193_5,  s_192_5, 
 s_191_6,  s_190_6,  s_189_7,  s_188_7,  s_187_8,  s_186_8, 
 s_185_9,  s_184_9, s_183_10, s_182_10, s_181_11, s_180_11, 
s_179_12, s_178_12, s_177_13, s_176_13, s_175_14, s_174_14, 
s_173_15, s_172_15, s_171_16, s_170_16, s_169_17, s_168_17, 
s_167_18, s_166_18, s_165_19, s_164_19, s_163_20, s_162_20, 
s_161_21, s_160_21, s_159_22, s_158_22, s_157_23, s_156_23, 
s_155_24, s_154_24, s_153_25, s_152_25, s_151_26, s_150_26, 
s_149_27, s_148_27, s_147_28, s_146_28, s_145_29, s_144_29, 
s_143_30, s_142_30, s_141_31, s_140_31, s_139_32, s_138_32, 
s_137_33, s_136_33, s_135_34, s_134_34, s_133_35, s_132_35, 
s_131_36, s_130_36, s_129_37, s_128_37, s_127_37, s_126_37, 
s_125_37, s_124_37, s_123_37, s_122_37, s_121_37, s_120_37, 
s_119_37, s_118_37, s_117_37, s_116_37, s_115_37, s_114_37, 
s_113_37, s_112_37, s_111_37, s_110_37, s_109_37, s_108_37, 
s_107_37, s_106_37, s_105_37, s_104_37, s_103_37, s_102_37, 
s_101_37, s_100_37,  s_99_37,  s_98_37,  s_97_37,  s_96_37, 
 s_95_37,  s_94_37,  s_93_37,  s_92_37,  s_91_37,  s_90_37, 
 s_89_37,  s_88_37,  s_87_37,  s_86_37,  s_85_37,  s_84_37, 
 s_83_37,  s_82_37,  s_81_37,  s_80_37,  s_79_37,  s_78_37, 
 s_77_37,  s_76_37,  s_75_37,  s_74_37
} = partial_products[(width+2)*(37+1)-1:(width+2)*37];

assign {
 s_205_0,  s_204_0,  s_203_1,  s_202_1,  s_201_2,  s_200_2, 
 s_199_3,  s_198_3,  s_197_4,  s_196_4,  s_195_5,  s_194_5, 
 s_193_6,  s_192_6,  s_191_7,  s_190_7,  s_189_8,  s_188_8, 
 s_187_9,  s_186_9, s_185_10, s_184_10, s_183_11, s_182_11, 
s_181_12, s_180_12, s_179_13, s_178_13, s_177_14, s_176_14, 
s_175_15, s_174_15, s_173_16, s_172_16, s_171_17, s_170_17, 
s_169_18, s_168_18, s_167_19, s_166_19, s_165_20, s_164_20, 
s_163_21, s_162_21, s_161_22, s_160_22, s_159_23, s_158_23, 
s_157_24, s_156_24, s_155_25, s_154_25, s_153_26, s_152_26, 
s_151_27, s_150_27, s_149_28, s_148_28, s_147_29, s_146_29, 
s_145_30, s_144_30, s_143_31, s_142_31, s_141_32, s_140_32, 
s_139_33, s_138_33, s_137_34, s_136_34, s_135_35, s_134_35, 
s_133_36, s_132_36, s_131_37, s_130_37, s_129_38, s_128_38, 
s_127_38, s_126_38, s_125_38, s_124_38, s_123_38, s_122_38, 
s_121_38, s_120_38, s_119_38, s_118_38, s_117_38, s_116_38, 
s_115_38, s_114_38, s_113_38, s_112_38, s_111_38, s_110_38, 
s_109_38, s_108_38, s_107_38, s_106_38, s_105_38, s_104_38, 
s_103_38, s_102_38, s_101_38, s_100_38,  s_99_38,  s_98_38, 
 s_97_38,  s_96_38,  s_95_38,  s_94_38,  s_93_38,  s_92_38, 
 s_91_38,  s_90_38,  s_89_38,  s_88_38,  s_87_38,  s_86_38, 
 s_85_38,  s_84_38,  s_83_38,  s_82_38,  s_81_38,  s_80_38, 
 s_79_38,  s_78_38,  s_77_38,  s_76_38
} = partial_products[(width+2)*(38+1)-1:(width+2)*38];

assign {
 s_207_0,  s_206_0,  s_205_1,  s_204_1,  s_203_2,  s_202_2, 
 s_201_3,  s_200_3,  s_199_4,  s_198_4,  s_197_5,  s_196_5, 
 s_195_6,  s_194_6,  s_193_7,  s_192_7,  s_191_8,  s_190_8, 
 s_189_9,  s_188_9, s_187_10, s_186_10, s_185_11, s_184_11, 
s_183_12, s_182_12, s_181_13, s_180_13, s_179_14, s_178_14, 
s_177_15, s_176_15, s_175_16, s_174_16, s_173_17, s_172_17, 
s_171_18, s_170_18, s_169_19, s_168_19, s_167_20, s_166_20, 
s_165_21, s_164_21, s_163_22, s_162_22, s_161_23, s_160_23, 
s_159_24, s_158_24, s_157_25, s_156_25, s_155_26, s_154_26, 
s_153_27, s_152_27, s_151_28, s_150_28, s_149_29, s_148_29, 
s_147_30, s_146_30, s_145_31, s_144_31, s_143_32, s_142_32, 
s_141_33, s_140_33, s_139_34, s_138_34, s_137_35, s_136_35, 
s_135_36, s_134_36, s_133_37, s_132_37, s_131_38, s_130_38, 
s_129_39, s_128_39, s_127_39, s_126_39, s_125_39, s_124_39, 
s_123_39, s_122_39, s_121_39, s_120_39, s_119_39, s_118_39, 
s_117_39, s_116_39, s_115_39, s_114_39, s_113_39, s_112_39, 
s_111_39, s_110_39, s_109_39, s_108_39, s_107_39, s_106_39, 
s_105_39, s_104_39, s_103_39, s_102_39, s_101_39, s_100_39, 
 s_99_39,  s_98_39,  s_97_39,  s_96_39,  s_95_39,  s_94_39, 
 s_93_39,  s_92_39,  s_91_39,  s_90_39,  s_89_39,  s_88_39, 
 s_87_39,  s_86_39,  s_85_39,  s_84_39,  s_83_39,  s_82_39, 
 s_81_39,  s_80_39,  s_79_39,  s_78_39
} = partial_products[(width+2)*(39+1)-1:(width+2)*39];

assign {
 s_209_0,  s_208_0,  s_207_1,  s_206_1,  s_205_2,  s_204_2, 
 s_203_3,  s_202_3,  s_201_4,  s_200_4,  s_199_5,  s_198_5, 
 s_197_6,  s_196_6,  s_195_7,  s_194_7,  s_193_8,  s_192_8, 
 s_191_9,  s_190_9, s_189_10, s_188_10, s_187_11, s_186_11, 
s_185_12, s_184_12, s_183_13, s_182_13, s_181_14, s_180_14, 
s_179_15, s_178_15, s_177_16, s_176_16, s_175_17, s_174_17, 
s_173_18, s_172_18, s_171_19, s_170_19, s_169_20, s_168_20, 
s_167_21, s_166_21, s_165_22, s_164_22, s_163_23, s_162_23, 
s_161_24, s_160_24, s_159_25, s_158_25, s_157_26, s_156_26, 
s_155_27, s_154_27, s_153_28, s_152_28, s_151_29, s_150_29, 
s_149_30, s_148_30, s_147_31, s_146_31, s_145_32, s_144_32, 
s_143_33, s_142_33, s_141_34, s_140_34, s_139_35, s_138_35, 
s_137_36, s_136_36, s_135_37, s_134_37, s_133_38, s_132_38, 
s_131_39, s_130_39, s_129_40, s_128_40, s_127_40, s_126_40, 
s_125_40, s_124_40, s_123_40, s_122_40, s_121_40, s_120_40, 
s_119_40, s_118_40, s_117_40, s_116_40, s_115_40, s_114_40, 
s_113_40, s_112_40, s_111_40, s_110_40, s_109_40, s_108_40, 
s_107_40, s_106_40, s_105_40, s_104_40, s_103_40, s_102_40, 
s_101_40, s_100_40,  s_99_40,  s_98_40,  s_97_40,  s_96_40, 
 s_95_40,  s_94_40,  s_93_40,  s_92_40,  s_91_40,  s_90_40, 
 s_89_40,  s_88_40,  s_87_40,  s_86_40,  s_85_40,  s_84_40, 
 s_83_40,  s_82_40,  s_81_40,  s_80_40
} = partial_products[(width+2)*(40+1)-1:(width+2)*40];

assign {
 s_211_0,  s_210_0,  s_209_1,  s_208_1,  s_207_2,  s_206_2, 
 s_205_3,  s_204_3,  s_203_4,  s_202_4,  s_201_5,  s_200_5, 
 s_199_6,  s_198_6,  s_197_7,  s_196_7,  s_195_8,  s_194_8, 
 s_193_9,  s_192_9, s_191_10, s_190_10, s_189_11, s_188_11, 
s_187_12, s_186_12, s_185_13, s_184_13, s_183_14, s_182_14, 
s_181_15, s_180_15, s_179_16, s_178_16, s_177_17, s_176_17, 
s_175_18, s_174_18, s_173_19, s_172_19, s_171_20, s_170_20, 
s_169_21, s_168_21, s_167_22, s_166_22, s_165_23, s_164_23, 
s_163_24, s_162_24, s_161_25, s_160_25, s_159_26, s_158_26, 
s_157_27, s_156_27, s_155_28, s_154_28, s_153_29, s_152_29, 
s_151_30, s_150_30, s_149_31, s_148_31, s_147_32, s_146_32, 
s_145_33, s_144_33, s_143_34, s_142_34, s_141_35, s_140_35, 
s_139_36, s_138_36, s_137_37, s_136_37, s_135_38, s_134_38, 
s_133_39, s_132_39, s_131_40, s_130_40, s_129_41, s_128_41, 
s_127_41, s_126_41, s_125_41, s_124_41, s_123_41, s_122_41, 
s_121_41, s_120_41, s_119_41, s_118_41, s_117_41, s_116_41, 
s_115_41, s_114_41, s_113_41, s_112_41, s_111_41, s_110_41, 
s_109_41, s_108_41, s_107_41, s_106_41, s_105_41, s_104_41, 
s_103_41, s_102_41, s_101_41, s_100_41,  s_99_41,  s_98_41, 
 s_97_41,  s_96_41,  s_95_41,  s_94_41,  s_93_41,  s_92_41, 
 s_91_41,  s_90_41,  s_89_41,  s_88_41,  s_87_41,  s_86_41, 
 s_85_41,  s_84_41,  s_83_41,  s_82_41
} = partial_products[(width+2)*(41+1)-1:(width+2)*41];

assign {
 s_213_0,  s_212_0,  s_211_1,  s_210_1,  s_209_2,  s_208_2, 
 s_207_3,  s_206_3,  s_205_4,  s_204_4,  s_203_5,  s_202_5, 
 s_201_6,  s_200_6,  s_199_7,  s_198_7,  s_197_8,  s_196_8, 
 s_195_9,  s_194_9, s_193_10, s_192_10, s_191_11, s_190_11, 
s_189_12, s_188_12, s_187_13, s_186_13, s_185_14, s_184_14, 
s_183_15, s_182_15, s_181_16, s_180_16, s_179_17, s_178_17, 
s_177_18, s_176_18, s_175_19, s_174_19, s_173_20, s_172_20, 
s_171_21, s_170_21, s_169_22, s_168_22, s_167_23, s_166_23, 
s_165_24, s_164_24, s_163_25, s_162_25, s_161_26, s_160_26, 
s_159_27, s_158_27, s_157_28, s_156_28, s_155_29, s_154_29, 
s_153_30, s_152_30, s_151_31, s_150_31, s_149_32, s_148_32, 
s_147_33, s_146_33, s_145_34, s_144_34, s_143_35, s_142_35, 
s_141_36, s_140_36, s_139_37, s_138_37, s_137_38, s_136_38, 
s_135_39, s_134_39, s_133_40, s_132_40, s_131_41, s_130_41, 
s_129_42, s_128_42, s_127_42, s_126_42, s_125_42, s_124_42, 
s_123_42, s_122_42, s_121_42, s_120_42, s_119_42, s_118_42, 
s_117_42, s_116_42, s_115_42, s_114_42, s_113_42, s_112_42, 
s_111_42, s_110_42, s_109_42, s_108_42, s_107_42, s_106_42, 
s_105_42, s_104_42, s_103_42, s_102_42, s_101_42, s_100_42, 
 s_99_42,  s_98_42,  s_97_42,  s_96_42,  s_95_42,  s_94_42, 
 s_93_42,  s_92_42,  s_91_42,  s_90_42,  s_89_42,  s_88_42, 
 s_87_42,  s_86_42,  s_85_42,  s_84_42
} = partial_products[(width+2)*(42+1)-1:(width+2)*42];

assign {
 s_215_0,  s_214_0,  s_213_1,  s_212_1,  s_211_2,  s_210_2, 
 s_209_3,  s_208_3,  s_207_4,  s_206_4,  s_205_5,  s_204_5, 
 s_203_6,  s_202_6,  s_201_7,  s_200_7,  s_199_8,  s_198_8, 
 s_197_9,  s_196_9, s_195_10, s_194_10, s_193_11, s_192_11, 
s_191_12, s_190_12, s_189_13, s_188_13, s_187_14, s_186_14, 
s_185_15, s_184_15, s_183_16, s_182_16, s_181_17, s_180_17, 
s_179_18, s_178_18, s_177_19, s_176_19, s_175_20, s_174_20, 
s_173_21, s_172_21, s_171_22, s_170_22, s_169_23, s_168_23, 
s_167_24, s_166_24, s_165_25, s_164_25, s_163_26, s_162_26, 
s_161_27, s_160_27, s_159_28, s_158_28, s_157_29, s_156_29, 
s_155_30, s_154_30, s_153_31, s_152_31, s_151_32, s_150_32, 
s_149_33, s_148_33, s_147_34, s_146_34, s_145_35, s_144_35, 
s_143_36, s_142_36, s_141_37, s_140_37, s_139_38, s_138_38, 
s_137_39, s_136_39, s_135_40, s_134_40, s_133_41, s_132_41, 
s_131_42, s_130_42, s_129_43, s_128_43, s_127_43, s_126_43, 
s_125_43, s_124_43, s_123_43, s_122_43, s_121_43, s_120_43, 
s_119_43, s_118_43, s_117_43, s_116_43, s_115_43, s_114_43, 
s_113_43, s_112_43, s_111_43, s_110_43, s_109_43, s_108_43, 
s_107_43, s_106_43, s_105_43, s_104_43, s_103_43, s_102_43, 
s_101_43, s_100_43,  s_99_43,  s_98_43,  s_97_43,  s_96_43, 
 s_95_43,  s_94_43,  s_93_43,  s_92_43,  s_91_43,  s_90_43, 
 s_89_43,  s_88_43,  s_87_43,  s_86_43
} = partial_products[(width+2)*(43+1)-1:(width+2)*43];

assign {
 s_217_0,  s_216_0,  s_215_1,  s_214_1,  s_213_2,  s_212_2, 
 s_211_3,  s_210_3,  s_209_4,  s_208_4,  s_207_5,  s_206_5, 
 s_205_6,  s_204_6,  s_203_7,  s_202_7,  s_201_8,  s_200_8, 
 s_199_9,  s_198_9, s_197_10, s_196_10, s_195_11, s_194_11, 
s_193_12, s_192_12, s_191_13, s_190_13, s_189_14, s_188_14, 
s_187_15, s_186_15, s_185_16, s_184_16, s_183_17, s_182_17, 
s_181_18, s_180_18, s_179_19, s_178_19, s_177_20, s_176_20, 
s_175_21, s_174_21, s_173_22, s_172_22, s_171_23, s_170_23, 
s_169_24, s_168_24, s_167_25, s_166_25, s_165_26, s_164_26, 
s_163_27, s_162_27, s_161_28, s_160_28, s_159_29, s_158_29, 
s_157_30, s_156_30, s_155_31, s_154_31, s_153_32, s_152_32, 
s_151_33, s_150_33, s_149_34, s_148_34, s_147_35, s_146_35, 
s_145_36, s_144_36, s_143_37, s_142_37, s_141_38, s_140_38, 
s_139_39, s_138_39, s_137_40, s_136_40, s_135_41, s_134_41, 
s_133_42, s_132_42, s_131_43, s_130_43, s_129_44, s_128_44, 
s_127_44, s_126_44, s_125_44, s_124_44, s_123_44, s_122_44, 
s_121_44, s_120_44, s_119_44, s_118_44, s_117_44, s_116_44, 
s_115_44, s_114_44, s_113_44, s_112_44, s_111_44, s_110_44, 
s_109_44, s_108_44, s_107_44, s_106_44, s_105_44, s_104_44, 
s_103_44, s_102_44, s_101_44, s_100_44,  s_99_44,  s_98_44, 
 s_97_44,  s_96_44,  s_95_44,  s_94_44,  s_93_44,  s_92_44, 
 s_91_44,  s_90_44,  s_89_44,  s_88_44
} = partial_products[(width+2)*(44+1)-1:(width+2)*44];

assign {
 s_219_0,  s_218_0,  s_217_1,  s_216_1,  s_215_2,  s_214_2, 
 s_213_3,  s_212_3,  s_211_4,  s_210_4,  s_209_5,  s_208_5, 
 s_207_6,  s_206_6,  s_205_7,  s_204_7,  s_203_8,  s_202_8, 
 s_201_9,  s_200_9, s_199_10, s_198_10, s_197_11, s_196_11, 
s_195_12, s_194_12, s_193_13, s_192_13, s_191_14, s_190_14, 
s_189_15, s_188_15, s_187_16, s_186_16, s_185_17, s_184_17, 
s_183_18, s_182_18, s_181_19, s_180_19, s_179_20, s_178_20, 
s_177_21, s_176_21, s_175_22, s_174_22, s_173_23, s_172_23, 
s_171_24, s_170_24, s_169_25, s_168_25, s_167_26, s_166_26, 
s_165_27, s_164_27, s_163_28, s_162_28, s_161_29, s_160_29, 
s_159_30, s_158_30, s_157_31, s_156_31, s_155_32, s_154_32, 
s_153_33, s_152_33, s_151_34, s_150_34, s_149_35, s_148_35, 
s_147_36, s_146_36, s_145_37, s_144_37, s_143_38, s_142_38, 
s_141_39, s_140_39, s_139_40, s_138_40, s_137_41, s_136_41, 
s_135_42, s_134_42, s_133_43, s_132_43, s_131_44, s_130_44, 
s_129_45, s_128_45, s_127_45, s_126_45, s_125_45, s_124_45, 
s_123_45, s_122_45, s_121_45, s_120_45, s_119_45, s_118_45, 
s_117_45, s_116_45, s_115_45, s_114_45, s_113_45, s_112_45, 
s_111_45, s_110_45, s_109_45, s_108_45, s_107_45, s_106_45, 
s_105_45, s_104_45, s_103_45, s_102_45, s_101_45, s_100_45, 
 s_99_45,  s_98_45,  s_97_45,  s_96_45,  s_95_45,  s_94_45, 
 s_93_45,  s_92_45,  s_91_45,  s_90_45
} = partial_products[(width+2)*(45+1)-1:(width+2)*45];

assign {
 s_221_0,  s_220_0,  s_219_1,  s_218_1,  s_217_2,  s_216_2, 
 s_215_3,  s_214_3,  s_213_4,  s_212_4,  s_211_5,  s_210_5, 
 s_209_6,  s_208_6,  s_207_7,  s_206_7,  s_205_8,  s_204_8, 
 s_203_9,  s_202_9, s_201_10, s_200_10, s_199_11, s_198_11, 
s_197_12, s_196_12, s_195_13, s_194_13, s_193_14, s_192_14, 
s_191_15, s_190_15, s_189_16, s_188_16, s_187_17, s_186_17, 
s_185_18, s_184_18, s_183_19, s_182_19, s_181_20, s_180_20, 
s_179_21, s_178_21, s_177_22, s_176_22, s_175_23, s_174_23, 
s_173_24, s_172_24, s_171_25, s_170_25, s_169_26, s_168_26, 
s_167_27, s_166_27, s_165_28, s_164_28, s_163_29, s_162_29, 
s_161_30, s_160_30, s_159_31, s_158_31, s_157_32, s_156_32, 
s_155_33, s_154_33, s_153_34, s_152_34, s_151_35, s_150_35, 
s_149_36, s_148_36, s_147_37, s_146_37, s_145_38, s_144_38, 
s_143_39, s_142_39, s_141_40, s_140_40, s_139_41, s_138_41, 
s_137_42, s_136_42, s_135_43, s_134_43, s_133_44, s_132_44, 
s_131_45, s_130_45, s_129_46, s_128_46, s_127_46, s_126_46, 
s_125_46, s_124_46, s_123_46, s_122_46, s_121_46, s_120_46, 
s_119_46, s_118_46, s_117_46, s_116_46, s_115_46, s_114_46, 
s_113_46, s_112_46, s_111_46, s_110_46, s_109_46, s_108_46, 
s_107_46, s_106_46, s_105_46, s_104_46, s_103_46, s_102_46, 
s_101_46, s_100_46,  s_99_46,  s_98_46,  s_97_46,  s_96_46, 
 s_95_46,  s_94_46,  s_93_46,  s_92_46
} = partial_products[(width+2)*(46+1)-1:(width+2)*46];

assign {
 s_223_0,  s_222_0,  s_221_1,  s_220_1,  s_219_2,  s_218_2, 
 s_217_3,  s_216_3,  s_215_4,  s_214_4,  s_213_5,  s_212_5, 
 s_211_6,  s_210_6,  s_209_7,  s_208_7,  s_207_8,  s_206_8, 
 s_205_9,  s_204_9, s_203_10, s_202_10, s_201_11, s_200_11, 
s_199_12, s_198_12, s_197_13, s_196_13, s_195_14, s_194_14, 
s_193_15, s_192_15, s_191_16, s_190_16, s_189_17, s_188_17, 
s_187_18, s_186_18, s_185_19, s_184_19, s_183_20, s_182_20, 
s_181_21, s_180_21, s_179_22, s_178_22, s_177_23, s_176_23, 
s_175_24, s_174_24, s_173_25, s_172_25, s_171_26, s_170_26, 
s_169_27, s_168_27, s_167_28, s_166_28, s_165_29, s_164_29, 
s_163_30, s_162_30, s_161_31, s_160_31, s_159_32, s_158_32, 
s_157_33, s_156_33, s_155_34, s_154_34, s_153_35, s_152_35, 
s_151_36, s_150_36, s_149_37, s_148_37, s_147_38, s_146_38, 
s_145_39, s_144_39, s_143_40, s_142_40, s_141_41, s_140_41, 
s_139_42, s_138_42, s_137_43, s_136_43, s_135_44, s_134_44, 
s_133_45, s_132_45, s_131_46, s_130_46, s_129_47, s_128_47, 
s_127_47, s_126_47, s_125_47, s_124_47, s_123_47, s_122_47, 
s_121_47, s_120_47, s_119_47, s_118_47, s_117_47, s_116_47, 
s_115_47, s_114_47, s_113_47, s_112_47, s_111_47, s_110_47, 
s_109_47, s_108_47, s_107_47, s_106_47, s_105_47, s_104_47, 
s_103_47, s_102_47, s_101_47, s_100_47,  s_99_47,  s_98_47, 
 s_97_47,  s_96_47,  s_95_47,  s_94_47
} = partial_products[(width+2)*(47+1)-1:(width+2)*47];

assign {
 s_225_0,  s_224_0,  s_223_1,  s_222_1,  s_221_2,  s_220_2, 
 s_219_3,  s_218_3,  s_217_4,  s_216_4,  s_215_5,  s_214_5, 
 s_213_6,  s_212_6,  s_211_7,  s_210_7,  s_209_8,  s_208_8, 
 s_207_9,  s_206_9, s_205_10, s_204_10, s_203_11, s_202_11, 
s_201_12, s_200_12, s_199_13, s_198_13, s_197_14, s_196_14, 
s_195_15, s_194_15, s_193_16, s_192_16, s_191_17, s_190_17, 
s_189_18, s_188_18, s_187_19, s_186_19, s_185_20, s_184_20, 
s_183_21, s_182_21, s_181_22, s_180_22, s_179_23, s_178_23, 
s_177_24, s_176_24, s_175_25, s_174_25, s_173_26, s_172_26, 
s_171_27, s_170_27, s_169_28, s_168_28, s_167_29, s_166_29, 
s_165_30, s_164_30, s_163_31, s_162_31, s_161_32, s_160_32, 
s_159_33, s_158_33, s_157_34, s_156_34, s_155_35, s_154_35, 
s_153_36, s_152_36, s_151_37, s_150_37, s_149_38, s_148_38, 
s_147_39, s_146_39, s_145_40, s_144_40, s_143_41, s_142_41, 
s_141_42, s_140_42, s_139_43, s_138_43, s_137_44, s_136_44, 
s_135_45, s_134_45, s_133_46, s_132_46, s_131_47, s_130_47, 
s_129_48, s_128_48, s_127_48, s_126_48, s_125_48, s_124_48, 
s_123_48, s_122_48, s_121_48, s_120_48, s_119_48, s_118_48, 
s_117_48, s_116_48, s_115_48, s_114_48, s_113_48, s_112_48, 
s_111_48, s_110_48, s_109_48, s_108_48, s_107_48, s_106_48, 
s_105_48, s_104_48, s_103_48, s_102_48, s_101_48, s_100_48, 
 s_99_48,  s_98_48,  s_97_48,  s_96_48
} = partial_products[(width+2)*(48+1)-1:(width+2)*48];

assign {
 s_227_0,  s_226_0,  s_225_1,  s_224_1,  s_223_2,  s_222_2, 
 s_221_3,  s_220_3,  s_219_4,  s_218_4,  s_217_5,  s_216_5, 
 s_215_6,  s_214_6,  s_213_7,  s_212_7,  s_211_8,  s_210_8, 
 s_209_9,  s_208_9, s_207_10, s_206_10, s_205_11, s_204_11, 
s_203_12, s_202_12, s_201_13, s_200_13, s_199_14, s_198_14, 
s_197_15, s_196_15, s_195_16, s_194_16, s_193_17, s_192_17, 
s_191_18, s_190_18, s_189_19, s_188_19, s_187_20, s_186_20, 
s_185_21, s_184_21, s_183_22, s_182_22, s_181_23, s_180_23, 
s_179_24, s_178_24, s_177_25, s_176_25, s_175_26, s_174_26, 
s_173_27, s_172_27, s_171_28, s_170_28, s_169_29, s_168_29, 
s_167_30, s_166_30, s_165_31, s_164_31, s_163_32, s_162_32, 
s_161_33, s_160_33, s_159_34, s_158_34, s_157_35, s_156_35, 
s_155_36, s_154_36, s_153_37, s_152_37, s_151_38, s_150_38, 
s_149_39, s_148_39, s_147_40, s_146_40, s_145_41, s_144_41, 
s_143_42, s_142_42, s_141_43, s_140_43, s_139_44, s_138_44, 
s_137_45, s_136_45, s_135_46, s_134_46, s_133_47, s_132_47, 
s_131_48, s_130_48, s_129_49, s_128_49, s_127_49, s_126_49, 
s_125_49, s_124_49, s_123_49, s_122_49, s_121_49, s_120_49, 
s_119_49, s_118_49, s_117_49, s_116_49, s_115_49, s_114_49, 
s_113_49, s_112_49, s_111_49, s_110_49, s_109_49, s_108_49, 
s_107_49, s_106_49, s_105_49, s_104_49, s_103_49, s_102_49, 
s_101_49, s_100_49,  s_99_49,  s_98_49
} = partial_products[(width+2)*(49+1)-1:(width+2)*49];

assign {
 s_229_0,  s_228_0,  s_227_1,  s_226_1,  s_225_2,  s_224_2, 
 s_223_3,  s_222_3,  s_221_4,  s_220_4,  s_219_5,  s_218_5, 
 s_217_6,  s_216_6,  s_215_7,  s_214_7,  s_213_8,  s_212_8, 
 s_211_9,  s_210_9, s_209_10, s_208_10, s_207_11, s_206_11, 
s_205_12, s_204_12, s_203_13, s_202_13, s_201_14, s_200_14, 
s_199_15, s_198_15, s_197_16, s_196_16, s_195_17, s_194_17, 
s_193_18, s_192_18, s_191_19, s_190_19, s_189_20, s_188_20, 
s_187_21, s_186_21, s_185_22, s_184_22, s_183_23, s_182_23, 
s_181_24, s_180_24, s_179_25, s_178_25, s_177_26, s_176_26, 
s_175_27, s_174_27, s_173_28, s_172_28, s_171_29, s_170_29, 
s_169_30, s_168_30, s_167_31, s_166_31, s_165_32, s_164_32, 
s_163_33, s_162_33, s_161_34, s_160_34, s_159_35, s_158_35, 
s_157_36, s_156_36, s_155_37, s_154_37, s_153_38, s_152_38, 
s_151_39, s_150_39, s_149_40, s_148_40, s_147_41, s_146_41, 
s_145_42, s_144_42, s_143_43, s_142_43, s_141_44, s_140_44, 
s_139_45, s_138_45, s_137_46, s_136_46, s_135_47, s_134_47, 
s_133_48, s_132_48, s_131_49, s_130_49, s_129_50, s_128_50, 
s_127_50, s_126_50, s_125_50, s_124_50, s_123_50, s_122_50, 
s_121_50, s_120_50, s_119_50, s_118_50, s_117_50, s_116_50, 
s_115_50, s_114_50, s_113_50, s_112_50, s_111_50, s_110_50, 
s_109_50, s_108_50, s_107_50, s_106_50, s_105_50, s_104_50, 
s_103_50, s_102_50, s_101_50, s_100_50
} = partial_products[(width+2)*(50+1)-1:(width+2)*50];

assign {
 s_231_0,  s_230_0,  s_229_1,  s_228_1,  s_227_2,  s_226_2, 
 s_225_3,  s_224_3,  s_223_4,  s_222_4,  s_221_5,  s_220_5, 
 s_219_6,  s_218_6,  s_217_7,  s_216_7,  s_215_8,  s_214_8, 
 s_213_9,  s_212_9, s_211_10, s_210_10, s_209_11, s_208_11, 
s_207_12, s_206_12, s_205_13, s_204_13, s_203_14, s_202_14, 
s_201_15, s_200_15, s_199_16, s_198_16, s_197_17, s_196_17, 
s_195_18, s_194_18, s_193_19, s_192_19, s_191_20, s_190_20, 
s_189_21, s_188_21, s_187_22, s_186_22, s_185_23, s_184_23, 
s_183_24, s_182_24, s_181_25, s_180_25, s_179_26, s_178_26, 
s_177_27, s_176_27, s_175_28, s_174_28, s_173_29, s_172_29, 
s_171_30, s_170_30, s_169_31, s_168_31, s_167_32, s_166_32, 
s_165_33, s_164_33, s_163_34, s_162_34, s_161_35, s_160_35, 
s_159_36, s_158_36, s_157_37, s_156_37, s_155_38, s_154_38, 
s_153_39, s_152_39, s_151_40, s_150_40, s_149_41, s_148_41, 
s_147_42, s_146_42, s_145_43, s_144_43, s_143_44, s_142_44, 
s_141_45, s_140_45, s_139_46, s_138_46, s_137_47, s_136_47, 
s_135_48, s_134_48, s_133_49, s_132_49, s_131_50, s_130_50, 
s_129_51, s_128_51, s_127_51, s_126_51, s_125_51, s_124_51, 
s_123_51, s_122_51, s_121_51, s_120_51, s_119_51, s_118_51, 
s_117_51, s_116_51, s_115_51, s_114_51, s_113_51, s_112_51, 
s_111_51, s_110_51, s_109_51, s_108_51, s_107_51, s_106_51, 
s_105_51, s_104_51, s_103_51, s_102_51
} = partial_products[(width+2)*(51+1)-1:(width+2)*51];

assign {
 s_233_0,  s_232_0,  s_231_1,  s_230_1,  s_229_2,  s_228_2, 
 s_227_3,  s_226_3,  s_225_4,  s_224_4,  s_223_5,  s_222_5, 
 s_221_6,  s_220_6,  s_219_7,  s_218_7,  s_217_8,  s_216_8, 
 s_215_9,  s_214_9, s_213_10, s_212_10, s_211_11, s_210_11, 
s_209_12, s_208_12, s_207_13, s_206_13, s_205_14, s_204_14, 
s_203_15, s_202_15, s_201_16, s_200_16, s_199_17, s_198_17, 
s_197_18, s_196_18, s_195_19, s_194_19, s_193_20, s_192_20, 
s_191_21, s_190_21, s_189_22, s_188_22, s_187_23, s_186_23, 
s_185_24, s_184_24, s_183_25, s_182_25, s_181_26, s_180_26, 
s_179_27, s_178_27, s_177_28, s_176_28, s_175_29, s_174_29, 
s_173_30, s_172_30, s_171_31, s_170_31, s_169_32, s_168_32, 
s_167_33, s_166_33, s_165_34, s_164_34, s_163_35, s_162_35, 
s_161_36, s_160_36, s_159_37, s_158_37, s_157_38, s_156_38, 
s_155_39, s_154_39, s_153_40, s_152_40, s_151_41, s_150_41, 
s_149_42, s_148_42, s_147_43, s_146_43, s_145_44, s_144_44, 
s_143_45, s_142_45, s_141_46, s_140_46, s_139_47, s_138_47, 
s_137_48, s_136_48, s_135_49, s_134_49, s_133_50, s_132_50, 
s_131_51, s_130_51, s_129_52, s_128_52, s_127_52, s_126_52, 
s_125_52, s_124_52, s_123_52, s_122_52, s_121_52, s_120_52, 
s_119_52, s_118_52, s_117_52, s_116_52, s_115_52, s_114_52, 
s_113_52, s_112_52, s_111_52, s_110_52, s_109_52, s_108_52, 
s_107_52, s_106_52, s_105_52, s_104_52
} = partial_products[(width+2)*(52+1)-1:(width+2)*52];

assign {
 s_235_0,  s_234_0,  s_233_1,  s_232_1,  s_231_2,  s_230_2, 
 s_229_3,  s_228_3,  s_227_4,  s_226_4,  s_225_5,  s_224_5, 
 s_223_6,  s_222_6,  s_221_7,  s_220_7,  s_219_8,  s_218_8, 
 s_217_9,  s_216_9, s_215_10, s_214_10, s_213_11, s_212_11, 
s_211_12, s_210_12, s_209_13, s_208_13, s_207_14, s_206_14, 
s_205_15, s_204_15, s_203_16, s_202_16, s_201_17, s_200_17, 
s_199_18, s_198_18, s_197_19, s_196_19, s_195_20, s_194_20, 
s_193_21, s_192_21, s_191_22, s_190_22, s_189_23, s_188_23, 
s_187_24, s_186_24, s_185_25, s_184_25, s_183_26, s_182_26, 
s_181_27, s_180_27, s_179_28, s_178_28, s_177_29, s_176_29, 
s_175_30, s_174_30, s_173_31, s_172_31, s_171_32, s_170_32, 
s_169_33, s_168_33, s_167_34, s_166_34, s_165_35, s_164_35, 
s_163_36, s_162_36, s_161_37, s_160_37, s_159_38, s_158_38, 
s_157_39, s_156_39, s_155_40, s_154_40, s_153_41, s_152_41, 
s_151_42, s_150_42, s_149_43, s_148_43, s_147_44, s_146_44, 
s_145_45, s_144_45, s_143_46, s_142_46, s_141_47, s_140_47, 
s_139_48, s_138_48, s_137_49, s_136_49, s_135_50, s_134_50, 
s_133_51, s_132_51, s_131_52, s_130_52, s_129_53, s_128_53, 
s_127_53, s_126_53, s_125_53, s_124_53, s_123_53, s_122_53, 
s_121_53, s_120_53, s_119_53, s_118_53, s_117_53, s_116_53, 
s_115_53, s_114_53, s_113_53, s_112_53, s_111_53, s_110_53, 
s_109_53, s_108_53, s_107_53, s_106_53
} = partial_products[(width+2)*(53+1)-1:(width+2)*53];

assign {
 s_237_0,  s_236_0,  s_235_1,  s_234_1,  s_233_2,  s_232_2, 
 s_231_3,  s_230_3,  s_229_4,  s_228_4,  s_227_5,  s_226_5, 
 s_225_6,  s_224_6,  s_223_7,  s_222_7,  s_221_8,  s_220_8, 
 s_219_9,  s_218_9, s_217_10, s_216_10, s_215_11, s_214_11, 
s_213_12, s_212_12, s_211_13, s_210_13, s_209_14, s_208_14, 
s_207_15, s_206_15, s_205_16, s_204_16, s_203_17, s_202_17, 
s_201_18, s_200_18, s_199_19, s_198_19, s_197_20, s_196_20, 
s_195_21, s_194_21, s_193_22, s_192_22, s_191_23, s_190_23, 
s_189_24, s_188_24, s_187_25, s_186_25, s_185_26, s_184_26, 
s_183_27, s_182_27, s_181_28, s_180_28, s_179_29, s_178_29, 
s_177_30, s_176_30, s_175_31, s_174_31, s_173_32, s_172_32, 
s_171_33, s_170_33, s_169_34, s_168_34, s_167_35, s_166_35, 
s_165_36, s_164_36, s_163_37, s_162_37, s_161_38, s_160_38, 
s_159_39, s_158_39, s_157_40, s_156_40, s_155_41, s_154_41, 
s_153_42, s_152_42, s_151_43, s_150_43, s_149_44, s_148_44, 
s_147_45, s_146_45, s_145_46, s_144_46, s_143_47, s_142_47, 
s_141_48, s_140_48, s_139_49, s_138_49, s_137_50, s_136_50, 
s_135_51, s_134_51, s_133_52, s_132_52, s_131_53, s_130_53, 
s_129_54, s_128_54, s_127_54, s_126_54, s_125_54, s_124_54, 
s_123_54, s_122_54, s_121_54, s_120_54, s_119_54, s_118_54, 
s_117_54, s_116_54, s_115_54, s_114_54, s_113_54, s_112_54, 
s_111_54, s_110_54, s_109_54, s_108_54
} = partial_products[(width+2)*(54+1)-1:(width+2)*54];

assign {
 s_239_0,  s_238_0,  s_237_1,  s_236_1,  s_235_2,  s_234_2, 
 s_233_3,  s_232_3,  s_231_4,  s_230_4,  s_229_5,  s_228_5, 
 s_227_6,  s_226_6,  s_225_7,  s_224_7,  s_223_8,  s_222_8, 
 s_221_9,  s_220_9, s_219_10, s_218_10, s_217_11, s_216_11, 
s_215_12, s_214_12, s_213_13, s_212_13, s_211_14, s_210_14, 
s_209_15, s_208_15, s_207_16, s_206_16, s_205_17, s_204_17, 
s_203_18, s_202_18, s_201_19, s_200_19, s_199_20, s_198_20, 
s_197_21, s_196_21, s_195_22, s_194_22, s_193_23, s_192_23, 
s_191_24, s_190_24, s_189_25, s_188_25, s_187_26, s_186_26, 
s_185_27, s_184_27, s_183_28, s_182_28, s_181_29, s_180_29, 
s_179_30, s_178_30, s_177_31, s_176_31, s_175_32, s_174_32, 
s_173_33, s_172_33, s_171_34, s_170_34, s_169_35, s_168_35, 
s_167_36, s_166_36, s_165_37, s_164_37, s_163_38, s_162_38, 
s_161_39, s_160_39, s_159_40, s_158_40, s_157_41, s_156_41, 
s_155_42, s_154_42, s_153_43, s_152_43, s_151_44, s_150_44, 
s_149_45, s_148_45, s_147_46, s_146_46, s_145_47, s_144_47, 
s_143_48, s_142_48, s_141_49, s_140_49, s_139_50, s_138_50, 
s_137_51, s_136_51, s_135_52, s_134_52, s_133_53, s_132_53, 
s_131_54, s_130_54, s_129_55, s_128_55, s_127_55, s_126_55, 
s_125_55, s_124_55, s_123_55, s_122_55, s_121_55, s_120_55, 
s_119_55, s_118_55, s_117_55, s_116_55, s_115_55, s_114_55, 
s_113_55, s_112_55, s_111_55, s_110_55
} = partial_products[(width+2)*(55+1)-1:(width+2)*55];

assign {
 s_241_0,  s_240_0,  s_239_1,  s_238_1,  s_237_2,  s_236_2, 
 s_235_3,  s_234_3,  s_233_4,  s_232_4,  s_231_5,  s_230_5, 
 s_229_6,  s_228_6,  s_227_7,  s_226_7,  s_225_8,  s_224_8, 
 s_223_9,  s_222_9, s_221_10, s_220_10, s_219_11, s_218_11, 
s_217_12, s_216_12, s_215_13, s_214_13, s_213_14, s_212_14, 
s_211_15, s_210_15, s_209_16, s_208_16, s_207_17, s_206_17, 
s_205_18, s_204_18, s_203_19, s_202_19, s_201_20, s_200_20, 
s_199_21, s_198_21, s_197_22, s_196_22, s_195_23, s_194_23, 
s_193_24, s_192_24, s_191_25, s_190_25, s_189_26, s_188_26, 
s_187_27, s_186_27, s_185_28, s_184_28, s_183_29, s_182_29, 
s_181_30, s_180_30, s_179_31, s_178_31, s_177_32, s_176_32, 
s_175_33, s_174_33, s_173_34, s_172_34, s_171_35, s_170_35, 
s_169_36, s_168_36, s_167_37, s_166_37, s_165_38, s_164_38, 
s_163_39, s_162_39, s_161_40, s_160_40, s_159_41, s_158_41, 
s_157_42, s_156_42, s_155_43, s_154_43, s_153_44, s_152_44, 
s_151_45, s_150_45, s_149_46, s_148_46, s_147_47, s_146_47, 
s_145_48, s_144_48, s_143_49, s_142_49, s_141_50, s_140_50, 
s_139_51, s_138_51, s_137_52, s_136_52, s_135_53, s_134_53, 
s_133_54, s_132_54, s_131_55, s_130_55, s_129_56, s_128_56, 
s_127_56, s_126_56, s_125_56, s_124_56, s_123_56, s_122_56, 
s_121_56, s_120_56, s_119_56, s_118_56, s_117_56, s_116_56, 
s_115_56, s_114_56, s_113_56, s_112_56
} = partial_products[(width+2)*(56+1)-1:(width+2)*56];

assign {
 s_243_0,  s_242_0,  s_241_1,  s_240_1,  s_239_2,  s_238_2, 
 s_237_3,  s_236_3,  s_235_4,  s_234_4,  s_233_5,  s_232_5, 
 s_231_6,  s_230_6,  s_229_7,  s_228_7,  s_227_8,  s_226_8, 
 s_225_9,  s_224_9, s_223_10, s_222_10, s_221_11, s_220_11, 
s_219_12, s_218_12, s_217_13, s_216_13, s_215_14, s_214_14, 
s_213_15, s_212_15, s_211_16, s_210_16, s_209_17, s_208_17, 
s_207_18, s_206_18, s_205_19, s_204_19, s_203_20, s_202_20, 
s_201_21, s_200_21, s_199_22, s_198_22, s_197_23, s_196_23, 
s_195_24, s_194_24, s_193_25, s_192_25, s_191_26, s_190_26, 
s_189_27, s_188_27, s_187_28, s_186_28, s_185_29, s_184_29, 
s_183_30, s_182_30, s_181_31, s_180_31, s_179_32, s_178_32, 
s_177_33, s_176_33, s_175_34, s_174_34, s_173_35, s_172_35, 
s_171_36, s_170_36, s_169_37, s_168_37, s_167_38, s_166_38, 
s_165_39, s_164_39, s_163_40, s_162_40, s_161_41, s_160_41, 
s_159_42, s_158_42, s_157_43, s_156_43, s_155_44, s_154_44, 
s_153_45, s_152_45, s_151_46, s_150_46, s_149_47, s_148_47, 
s_147_48, s_146_48, s_145_49, s_144_49, s_143_50, s_142_50, 
s_141_51, s_140_51, s_139_52, s_138_52, s_137_53, s_136_53, 
s_135_54, s_134_54, s_133_55, s_132_55, s_131_56, s_130_56, 
s_129_57, s_128_57, s_127_57, s_126_57, s_125_57, s_124_57, 
s_123_57, s_122_57, s_121_57, s_120_57, s_119_57, s_118_57, 
s_117_57, s_116_57, s_115_57, s_114_57
} = partial_products[(width+2)*(57+1)-1:(width+2)*57];

assign {
 s_245_0,  s_244_0,  s_243_1,  s_242_1,  s_241_2,  s_240_2, 
 s_239_3,  s_238_3,  s_237_4,  s_236_4,  s_235_5,  s_234_5, 
 s_233_6,  s_232_6,  s_231_7,  s_230_7,  s_229_8,  s_228_8, 
 s_227_9,  s_226_9, s_225_10, s_224_10, s_223_11, s_222_11, 
s_221_12, s_220_12, s_219_13, s_218_13, s_217_14, s_216_14, 
s_215_15, s_214_15, s_213_16, s_212_16, s_211_17, s_210_17, 
s_209_18, s_208_18, s_207_19, s_206_19, s_205_20, s_204_20, 
s_203_21, s_202_21, s_201_22, s_200_22, s_199_23, s_198_23, 
s_197_24, s_196_24, s_195_25, s_194_25, s_193_26, s_192_26, 
s_191_27, s_190_27, s_189_28, s_188_28, s_187_29, s_186_29, 
s_185_30, s_184_30, s_183_31, s_182_31, s_181_32, s_180_32, 
s_179_33, s_178_33, s_177_34, s_176_34, s_175_35, s_174_35, 
s_173_36, s_172_36, s_171_37, s_170_37, s_169_38, s_168_38, 
s_167_39, s_166_39, s_165_40, s_164_40, s_163_41, s_162_41, 
s_161_42, s_160_42, s_159_43, s_158_43, s_157_44, s_156_44, 
s_155_45, s_154_45, s_153_46, s_152_46, s_151_47, s_150_47, 
s_149_48, s_148_48, s_147_49, s_146_49, s_145_50, s_144_50, 
s_143_51, s_142_51, s_141_52, s_140_52, s_139_53, s_138_53, 
s_137_54, s_136_54, s_135_55, s_134_55, s_133_56, s_132_56, 
s_131_57, s_130_57, s_129_58, s_128_58, s_127_58, s_126_58, 
s_125_58, s_124_58, s_123_58, s_122_58, s_121_58, s_120_58, 
s_119_58, s_118_58, s_117_58, s_116_58
} = partial_products[(width+2)*(58+1)-1:(width+2)*58];

assign {
 s_247_0,  s_246_0,  s_245_1,  s_244_1,  s_243_2,  s_242_2, 
 s_241_3,  s_240_3,  s_239_4,  s_238_4,  s_237_5,  s_236_5, 
 s_235_6,  s_234_6,  s_233_7,  s_232_7,  s_231_8,  s_230_8, 
 s_229_9,  s_228_9, s_227_10, s_226_10, s_225_11, s_224_11, 
s_223_12, s_222_12, s_221_13, s_220_13, s_219_14, s_218_14, 
s_217_15, s_216_15, s_215_16, s_214_16, s_213_17, s_212_17, 
s_211_18, s_210_18, s_209_19, s_208_19, s_207_20, s_206_20, 
s_205_21, s_204_21, s_203_22, s_202_22, s_201_23, s_200_23, 
s_199_24, s_198_24, s_197_25, s_196_25, s_195_26, s_194_26, 
s_193_27, s_192_27, s_191_28, s_190_28, s_189_29, s_188_29, 
s_187_30, s_186_30, s_185_31, s_184_31, s_183_32, s_182_32, 
s_181_33, s_180_33, s_179_34, s_178_34, s_177_35, s_176_35, 
s_175_36, s_174_36, s_173_37, s_172_37, s_171_38, s_170_38, 
s_169_39, s_168_39, s_167_40, s_166_40, s_165_41, s_164_41, 
s_163_42, s_162_42, s_161_43, s_160_43, s_159_44, s_158_44, 
s_157_45, s_156_45, s_155_46, s_154_46, s_153_47, s_152_47, 
s_151_48, s_150_48, s_149_49, s_148_49, s_147_50, s_146_50, 
s_145_51, s_144_51, s_143_52, s_142_52, s_141_53, s_140_53, 
s_139_54, s_138_54, s_137_55, s_136_55, s_135_56, s_134_56, 
s_133_57, s_132_57, s_131_58, s_130_58, s_129_59, s_128_59, 
s_127_59, s_126_59, s_125_59, s_124_59, s_123_59, s_122_59, 
s_121_59, s_120_59, s_119_59, s_118_59
} = partial_products[(width+2)*(59+1)-1:(width+2)*59];

assign {
 s_249_0,  s_248_0,  s_247_1,  s_246_1,  s_245_2,  s_244_2, 
 s_243_3,  s_242_3,  s_241_4,  s_240_4,  s_239_5,  s_238_5, 
 s_237_6,  s_236_6,  s_235_7,  s_234_7,  s_233_8,  s_232_8, 
 s_231_9,  s_230_9, s_229_10, s_228_10, s_227_11, s_226_11, 
s_225_12, s_224_12, s_223_13, s_222_13, s_221_14, s_220_14, 
s_219_15, s_218_15, s_217_16, s_216_16, s_215_17, s_214_17, 
s_213_18, s_212_18, s_211_19, s_210_19, s_209_20, s_208_20, 
s_207_21, s_206_21, s_205_22, s_204_22, s_203_23, s_202_23, 
s_201_24, s_200_24, s_199_25, s_198_25, s_197_26, s_196_26, 
s_195_27, s_194_27, s_193_28, s_192_28, s_191_29, s_190_29, 
s_189_30, s_188_30, s_187_31, s_186_31, s_185_32, s_184_32, 
s_183_33, s_182_33, s_181_34, s_180_34, s_179_35, s_178_35, 
s_177_36, s_176_36, s_175_37, s_174_37, s_173_38, s_172_38, 
s_171_39, s_170_39, s_169_40, s_168_40, s_167_41, s_166_41, 
s_165_42, s_164_42, s_163_43, s_162_43, s_161_44, s_160_44, 
s_159_45, s_158_45, s_157_46, s_156_46, s_155_47, s_154_47, 
s_153_48, s_152_48, s_151_49, s_150_49, s_149_50, s_148_50, 
s_147_51, s_146_51, s_145_52, s_144_52, s_143_53, s_142_53, 
s_141_54, s_140_54, s_139_55, s_138_55, s_137_56, s_136_56, 
s_135_57, s_134_57, s_133_58, s_132_58, s_131_59, s_130_59, 
s_129_60, s_128_60, s_127_60, s_126_60, s_125_60, s_124_60, 
s_123_60, s_122_60, s_121_60, s_120_60
} = partial_products[(width+2)*(60+1)-1:(width+2)*60];

assign {
 s_251_0,  s_250_0,  s_249_1,  s_248_1,  s_247_2,  s_246_2, 
 s_245_3,  s_244_3,  s_243_4,  s_242_4,  s_241_5,  s_240_5, 
 s_239_6,  s_238_6,  s_237_7,  s_236_7,  s_235_8,  s_234_8, 
 s_233_9,  s_232_9, s_231_10, s_230_10, s_229_11, s_228_11, 
s_227_12, s_226_12, s_225_13, s_224_13, s_223_14, s_222_14, 
s_221_15, s_220_15, s_219_16, s_218_16, s_217_17, s_216_17, 
s_215_18, s_214_18, s_213_19, s_212_19, s_211_20, s_210_20, 
s_209_21, s_208_21, s_207_22, s_206_22, s_205_23, s_204_23, 
s_203_24, s_202_24, s_201_25, s_200_25, s_199_26, s_198_26, 
s_197_27, s_196_27, s_195_28, s_194_28, s_193_29, s_192_29, 
s_191_30, s_190_30, s_189_31, s_188_31, s_187_32, s_186_32, 
s_185_33, s_184_33, s_183_34, s_182_34, s_181_35, s_180_35, 
s_179_36, s_178_36, s_177_37, s_176_37, s_175_38, s_174_38, 
s_173_39, s_172_39, s_171_40, s_170_40, s_169_41, s_168_41, 
s_167_42, s_166_42, s_165_43, s_164_43, s_163_44, s_162_44, 
s_161_45, s_160_45, s_159_46, s_158_46, s_157_47, s_156_47, 
s_155_48, s_154_48, s_153_49, s_152_49, s_151_50, s_150_50, 
s_149_51, s_148_51, s_147_52, s_146_52, s_145_53, s_144_53, 
s_143_54, s_142_54, s_141_55, s_140_55, s_139_56, s_138_56, 
s_137_57, s_136_57, s_135_58, s_134_58, s_133_59, s_132_59, 
s_131_60, s_130_60, s_129_61, s_128_61, s_127_61, s_126_61, 
s_125_61, s_124_61, s_123_61, s_122_61
} = partial_products[(width+2)*(61+1)-1:(width+2)*61];

assign {
 s_253_0,  s_252_0,  s_251_1,  s_250_1,  s_249_2,  s_248_2, 
 s_247_3,  s_246_3,  s_245_4,  s_244_4,  s_243_5,  s_242_5, 
 s_241_6,  s_240_6,  s_239_7,  s_238_7,  s_237_8,  s_236_8, 
 s_235_9,  s_234_9, s_233_10, s_232_10, s_231_11, s_230_11, 
s_229_12, s_228_12, s_227_13, s_226_13, s_225_14, s_224_14, 
s_223_15, s_222_15, s_221_16, s_220_16, s_219_17, s_218_17, 
s_217_18, s_216_18, s_215_19, s_214_19, s_213_20, s_212_20, 
s_211_21, s_210_21, s_209_22, s_208_22, s_207_23, s_206_23, 
s_205_24, s_204_24, s_203_25, s_202_25, s_201_26, s_200_26, 
s_199_27, s_198_27, s_197_28, s_196_28, s_195_29, s_194_29, 
s_193_30, s_192_30, s_191_31, s_190_31, s_189_32, s_188_32, 
s_187_33, s_186_33, s_185_34, s_184_34, s_183_35, s_182_35, 
s_181_36, s_180_36, s_179_37, s_178_37, s_177_38, s_176_38, 
s_175_39, s_174_39, s_173_40, s_172_40, s_171_41, s_170_41, 
s_169_42, s_168_42, s_167_43, s_166_43, s_165_44, s_164_44, 
s_163_45, s_162_45, s_161_46, s_160_46, s_159_47, s_158_47, 
s_157_48, s_156_48, s_155_49, s_154_49, s_153_50, s_152_50, 
s_151_51, s_150_51, s_149_52, s_148_52, s_147_53, s_146_53, 
s_145_54, s_144_54, s_143_55, s_142_55, s_141_56, s_140_56, 
s_139_57, s_138_57, s_137_58, s_136_58, s_135_59, s_134_59, 
s_133_60, s_132_60, s_131_61, s_130_61, s_129_62, s_128_62, 
s_127_62, s_126_62, s_125_62, s_124_62
} = partial_products[(width+2)*(62+1)-1:(width+2)*62];

assign {
 s_255_0,  s_254_0,  s_253_1,  s_252_1,  s_251_2,  s_250_2, 
 s_249_3,  s_248_3,  s_247_4,  s_246_4,  s_245_5,  s_244_5, 
 s_243_6,  s_242_6,  s_241_7,  s_240_7,  s_239_8,  s_238_8, 
 s_237_9,  s_236_9, s_235_10, s_234_10, s_233_11, s_232_11, 
s_231_12, s_230_12, s_229_13, s_228_13, s_227_14, s_226_14, 
s_225_15, s_224_15, s_223_16, s_222_16, s_221_17, s_220_17, 
s_219_18, s_218_18, s_217_19, s_216_19, s_215_20, s_214_20, 
s_213_21, s_212_21, s_211_22, s_210_22, s_209_23, s_208_23, 
s_207_24, s_206_24, s_205_25, s_204_25, s_203_26, s_202_26, 
s_201_27, s_200_27, s_199_28, s_198_28, s_197_29, s_196_29, 
s_195_30, s_194_30, s_193_31, s_192_31, s_191_32, s_190_32, 
s_189_33, s_188_33, s_187_34, s_186_34, s_185_35, s_184_35, 
s_183_36, s_182_36, s_181_37, s_180_37, s_179_38, s_178_38, 
s_177_39, s_176_39, s_175_40, s_174_40, s_173_41, s_172_41, 
s_171_42, s_170_42, s_169_43, s_168_43, s_167_44, s_166_44, 
s_165_45, s_164_45, s_163_46, s_162_46, s_161_47, s_160_47, 
s_159_48, s_158_48, s_157_49, s_156_49, s_155_50, s_154_50, 
s_153_51, s_152_51, s_151_52, s_150_52, s_149_53, s_148_53, 
s_147_54, s_146_54, s_145_55, s_144_55, s_143_56, s_142_56, 
s_141_57, s_140_57, s_139_58, s_138_58, s_137_59, s_136_59, 
s_135_60, s_134_60, s_133_61, s_132_61, s_131_62, s_130_62, 
s_129_63, s_128_63, s_127_63, s_126_63
} = partial_products[(width+2)*(63+1)-1:(width+2)*63];

assign {
 s_255_1,  s_254_1,  s_253_2,  s_252_2,  s_251_3,  s_250_3, 
 s_249_4,  s_248_4,  s_247_5,  s_246_5,  s_245_6,  s_244_6, 
 s_243_7,  s_242_7,  s_241_8,  s_240_8,  s_239_9,  s_238_9, 
s_237_10, s_236_10, s_235_11, s_234_11, s_233_12, s_232_12, 
s_231_13, s_230_13, s_229_14, s_228_14, s_227_15, s_226_15, 
s_225_16, s_224_16, s_223_17, s_222_17, s_221_18, s_220_18, 
s_219_19, s_218_19, s_217_20, s_216_20, s_215_21, s_214_21, 
s_213_22, s_212_22, s_211_23, s_210_23, s_209_24, s_208_24, 
s_207_25, s_206_25, s_205_26, s_204_26, s_203_27, s_202_27, 
s_201_28, s_200_28, s_199_29, s_198_29, s_197_30, s_196_30, 
s_195_31, s_194_31, s_193_32, s_192_32, s_191_33, s_190_33, 
s_189_34, s_188_34, s_187_35, s_186_35, s_185_36, s_184_36, 
s_183_37, s_182_37, s_181_38, s_180_38, s_179_39, s_178_39, 
s_177_40, s_176_40, s_175_41, s_174_41, s_173_42, s_172_42, 
s_171_43, s_170_43, s_169_44, s_168_44, s_167_45, s_166_45, 
s_165_46, s_164_46, s_163_47, s_162_47, s_161_48, s_160_48, 
s_159_49, s_158_49, s_157_50, s_156_50, s_155_51, s_154_51, 
s_153_52, s_152_52, s_151_53, s_150_53, s_149_54, s_148_54, 
s_147_55, s_146_55, s_145_56, s_144_56, s_143_57, s_142_57, 
s_141_58, s_140_58, s_139_59, s_138_59, s_137_60, s_136_60, 
s_135_61, s_134_61, s_133_62, s_132_62, s_131_63, s_130_63, 
s_129_64, s_128_64
} = partial_products[(width+2)*(width/2+1)-1:(width+2)*width/2+2];

/* u0_1 Output nets */
wire t_0,      t_1;
/* u1_2 Output nets */
wire t_2,      t_3;
/* u0_3 Output nets */
wire t_4,      t_5;
/* u2_4 Output nets */
wire t_6,      t_7,      t_8;
/* u1_5 Output nets */
wire t_9,     t_10;
/* u2_6 Output nets */
wire t_11,     t_12,     t_13;
/* u2_7 Output nets */
wire t_14,     t_15,     t_16;
/* u2_8 Output nets */
wire t_17,     t_18,     t_19;
/* u0_9 Output nets */
wire t_20,     t_21;
/* u2_10 Output nets */
wire t_22,     t_23,     t_24;
/* u0_11 Output nets */
wire t_25,     t_26;
/* u2_12 Output nets */
wire t_27,     t_28,     t_29;
/* u1_13 Output nets */
wire t_30,     t_31;
/* u2_14 Output nets */
wire t_32,     t_33,     t_34;
/* u1_15 Output nets */
wire t_35,     t_36;
/* u2_16 Output nets */
wire t_37,     t_38,     t_39;
/* u2_17 Output nets */
wire t_40,     t_41,     t_42;
/* u2_18 Output nets */
wire t_43,     t_44,     t_45;
/* u1_19 Output nets */
wire t_46,     t_47;
/* u2_20 Output nets */
wire t_48,     t_49,     t_50;
/* u2_21 Output nets */
wire t_51,     t_52,     t_53;
/* u2_22 Output nets */
wire t_54,     t_55,     t_56;
/* u2_23 Output nets */
wire t_57,     t_58,     t_59;
/* u2_24 Output nets */
wire t_60,     t_61,     t_62;
/* u2_25 Output nets */
wire t_63,     t_64,     t_65;
/* u0_26 Output nets */
wire t_66,     t_67;
/* u2_27 Output nets */
wire t_68,     t_69,     t_70;
/* u2_28 Output nets */
wire t_71,     t_72,     t_73;
/* u0_29 Output nets */
wire t_74,     t_75;
/* u2_30 Output nets */
wire t_76,     t_77,     t_78;
/* u2_31 Output nets */
wire t_79,     t_80,     t_81;
/* u1_32 Output nets */
wire t_82,     t_83;
/* u2_33 Output nets */
wire t_84,     t_85,     t_86;
/* u2_34 Output nets */
wire t_87,     t_88,     t_89;
/* u1_35 Output nets */
wire t_90,     t_91;
/* u2_36 Output nets */
wire t_92,     t_93,     t_94;
/* u2_37 Output nets */
wire t_95,     t_96,     t_97;
/* u2_38 Output nets */
wire t_98,     t_99,    t_100;
/* u2_39 Output nets */
wire t_101,    t_102,    t_103;
/* u2_40 Output nets */
wire t_104,    t_105,    t_106;
/* u1_41 Output nets */
wire t_107,    t_108;
/* u2_42 Output nets */
wire t_109,    t_110,    t_111;
/* u2_43 Output nets */
wire t_112,    t_113,    t_114;
/* u2_44 Output nets */
wire t_115,    t_116,    t_117;
/* u2_45 Output nets */
wire t_118,    t_119,    t_120;
/* u2_46 Output nets */
wire t_121,    t_122,    t_123;
/* u2_47 Output nets */
wire t_124,    t_125,    t_126;
/* u2_48 Output nets */
wire t_127,    t_128,    t_129;
/* u2_49 Output nets */
wire t_130,    t_131,    t_132;
/* u2_50 Output nets */
wire t_133,    t_134,    t_135;
/* u0_51 Output nets */
wire t_136,    t_137;
/* u2_52 Output nets */
wire t_138,    t_139,    t_140;
/* u2_53 Output nets */
wire t_141,    t_142,    t_143;
/* u2_54 Output nets */
wire t_144,    t_145,    t_146;
/* u0_55 Output nets */
wire t_147,    t_148;
/* u2_56 Output nets */
wire t_149,    t_150,    t_151;
/* u2_57 Output nets */
wire t_152,    t_153,    t_154;
/* u2_58 Output nets */
wire t_155,    t_156,    t_157;
/* u1_59 Output nets */
wire t_158,    t_159;
/* u2_60 Output nets */
wire t_160,    t_161,    t_162;
/* u2_61 Output nets */
wire t_163,    t_164,    t_165;
/* u2_62 Output nets */
wire t_166,    t_167,    t_168;
/* u1_63 Output nets */
wire t_169,    t_170;
/* u2_64 Output nets */
wire t_171,    t_172,    t_173;
/* u2_65 Output nets */
wire t_174,    t_175,    t_176;
/* u2_66 Output nets */
wire t_177,    t_178,    t_179;
/* u2_67 Output nets */
wire t_180,    t_181,    t_182;
/* u2_68 Output nets */
wire t_183,    t_184,    t_185;
/* u2_69 Output nets */
wire t_186,    t_187,    t_188;
/* u2_70 Output nets */
wire t_189,    t_190,    t_191;
/* u1_71 Output nets */
wire t_192,    t_193;
/* u2_72 Output nets */
wire t_194,    t_195,    t_196;
/* u2_73 Output nets */
wire t_197,    t_198,    t_199;
/* u2_74 Output nets */
wire t_200,    t_201,    t_202;
/* u2_75 Output nets */
wire t_203,    t_204,    t_205;
/* u2_76 Output nets */
wire t_206,    t_207,    t_208;
/* u2_77 Output nets */
wire t_209,    t_210,    t_211;
/* u2_78 Output nets */
wire t_212,    t_213,    t_214;
/* u2_79 Output nets */
wire t_215,    t_216,    t_217;
/* u2_80 Output nets */
wire t_218,    t_219,    t_220;
/* u2_81 Output nets */
wire t_221,    t_222,    t_223;
/* u2_82 Output nets */
wire t_224,    t_225,    t_226;
/* u2_83 Output nets */
wire t_227,    t_228,    t_229;
/* u0_84 Output nets */
wire t_230,    t_231;
/* u2_85 Output nets */
wire t_232,    t_233,    t_234;
/* u2_86 Output nets */
wire t_235,    t_236,    t_237;
/* u2_87 Output nets */
wire t_238,    t_239,    t_240;
/* u2_88 Output nets */
wire t_241,    t_242,    t_243;
/* u0_89 Output nets */
wire t_244,    t_245;
/* u2_90 Output nets */
wire t_246,    t_247,    t_248;
/* u2_91 Output nets */
wire t_249,    t_250,    t_251;
/* u2_92 Output nets */
wire t_252,    t_253,    t_254;
/* u2_93 Output nets */
wire t_255,    t_256,    t_257;
/* u1_94 Output nets */
wire t_258,    t_259;
/* u2_95 Output nets */
wire t_260,    t_261,    t_262;
/* u2_96 Output nets */
wire t_263,    t_264,    t_265;
/* u2_97 Output nets */
wire t_266,    t_267,    t_268;
/* u2_98 Output nets */
wire t_269,    t_270,    t_271;
/* u1_99 Output nets */
wire t_272,    t_273;
/* u2_100 Output nets */
wire t_274,    t_275,    t_276;
/* u2_101 Output nets */
wire t_277,    t_278,    t_279;
/* u2_102 Output nets */
wire t_280,    t_281,    t_282;
/* u2_103 Output nets */
wire t_283,    t_284,    t_285;
/* u2_104 Output nets */
wire t_286,    t_287,    t_288;
/* u2_105 Output nets */
wire t_289,    t_290,    t_291;
/* u2_106 Output nets */
wire t_292,    t_293,    t_294;
/* u2_107 Output nets */
wire t_295,    t_296,    t_297;
/* u2_108 Output nets */
wire t_298,    t_299,    t_300;
/* u1_109 Output nets */
wire t_301,    t_302;
/* u2_110 Output nets */
wire t_303,    t_304,    t_305;
/* u2_111 Output nets */
wire t_306,    t_307,    t_308;
/* u2_112 Output nets */
wire t_309,    t_310,    t_311;
/* u2_113 Output nets */
wire t_312,    t_313,    t_314;
/* u2_114 Output nets */
wire t_315,    t_316,    t_317;
/* u2_115 Output nets */
wire t_318,    t_319,    t_320;
/* u2_116 Output nets */
wire t_321,    t_322,    t_323;
/* u2_117 Output nets */
wire t_324,    t_325,    t_326;
/* u2_118 Output nets */
wire t_327,    t_328,    t_329;
/* u2_119 Output nets */
wire t_330,    t_331,    t_332;
/* u2_120 Output nets */
wire t_333,    t_334,    t_335;
/* u2_121 Output nets */
wire t_336,    t_337,    t_338;
/* u2_122 Output nets */
wire t_339,    t_340,    t_341;
/* u2_123 Output nets */
wire t_342,    t_343,    t_344;
/* u2_124 Output nets */
wire t_345,    t_346,    t_347;
/* u0_125 Output nets */
wire t_348,    t_349;
/* u2_126 Output nets */
wire t_350,    t_351,    t_352;
/* u2_127 Output nets */
wire t_353,    t_354,    t_355;
/* u2_128 Output nets */
wire t_356,    t_357,    t_358;
/* u2_129 Output nets */
wire t_359,    t_360,    t_361;
/* u2_130 Output nets */
wire t_362,    t_363,    t_364;
/* u0_131 Output nets */
wire t_365,    t_366;
/* u2_132 Output nets */
wire t_367,    t_368,    t_369;
/* u2_133 Output nets */
wire t_370,    t_371,    t_372;
/* u2_134 Output nets */
wire t_373,    t_374,    t_375;
/* u2_135 Output nets */
wire t_376,    t_377,    t_378;
/* u2_136 Output nets */
wire t_379,    t_380,    t_381;
/* u1_137 Output nets */
wire t_382,    t_383;
/* u2_138 Output nets */
wire t_384,    t_385,    t_386;
/* u2_139 Output nets */
wire t_387,    t_388,    t_389;
/* u2_140 Output nets */
wire t_390,    t_391,    t_392;
/* u2_141 Output nets */
wire t_393,    t_394,    t_395;
/* u2_142 Output nets */
wire t_396,    t_397,    t_398;
/* u1_143 Output nets */
wire t_399,    t_400;
/* u2_144 Output nets */
wire t_401,    t_402,    t_403;
/* u2_145 Output nets */
wire t_404,    t_405,    t_406;
/* u2_146 Output nets */
wire t_407,    t_408,    t_409;
/* u2_147 Output nets */
wire t_410,    t_411,    t_412;
/* u2_148 Output nets */
wire t_413,    t_414,    t_415;
/* u2_149 Output nets */
wire t_416,    t_417,    t_418;
/* u2_150 Output nets */
wire t_419,    t_420,    t_421;
/* u2_151 Output nets */
wire t_422,    t_423,    t_424;
/* u2_152 Output nets */
wire t_425,    t_426,    t_427;
/* u2_153 Output nets */
wire t_428,    t_429,    t_430;
/* u2_154 Output nets */
wire t_431,    t_432,    t_433;
/* u1_155 Output nets */
wire t_434,    t_435;
/* u2_156 Output nets */
wire t_436,    t_437,    t_438;
/* u2_157 Output nets */
wire t_439,    t_440,    t_441;
/* u2_158 Output nets */
wire t_442,    t_443,    t_444;
/* u2_159 Output nets */
wire t_445,    t_446,    t_447;
/* u2_160 Output nets */
wire t_448,    t_449,    t_450;
/* u2_161 Output nets */
wire t_451,    t_452,    t_453;
/* u2_162 Output nets */
wire t_454,    t_455,    t_456;
/* u2_163 Output nets */
wire t_457,    t_458,    t_459;
/* u2_164 Output nets */
wire t_460,    t_461,    t_462;
/* u2_165 Output nets */
wire t_463,    t_464,    t_465;
/* u2_166 Output nets */
wire t_466,    t_467,    t_468;
/* u2_167 Output nets */
wire t_469,    t_470,    t_471;
/* u2_168 Output nets */
wire t_472,    t_473,    t_474;
/* u2_169 Output nets */
wire t_475,    t_476,    t_477;
/* u2_170 Output nets */
wire t_478,    t_479,    t_480;
/* u2_171 Output nets */
wire t_481,    t_482,    t_483;
/* u2_172 Output nets */
wire t_484,    t_485,    t_486;
/* u2_173 Output nets */
wire t_487,    t_488,    t_489;
/* u0_174 Output nets */
wire t_490,    t_491;
/* u2_175 Output nets */
wire t_492,    t_493,    t_494;
/* u2_176 Output nets */
wire t_495,    t_496,    t_497;
/* u2_177 Output nets */
wire t_498,    t_499,    t_500;
/* u2_178 Output nets */
wire t_501,    t_502,    t_503;
/* u2_179 Output nets */
wire t_504,    t_505,    t_506;
/* u2_180 Output nets */
wire t_507,    t_508,    t_509;
/* u0_181 Output nets */
wire t_510,    t_511;
/* u2_182 Output nets */
wire t_512,    t_513,    t_514;
/* u2_183 Output nets */
wire t_515,    t_516,    t_517;
/* u2_184 Output nets */
wire t_518,    t_519,    t_520;
/* u2_185 Output nets */
wire t_521,    t_522,    t_523;
/* u2_186 Output nets */
wire t_524,    t_525,    t_526;
/* u2_187 Output nets */
wire t_527,    t_528,    t_529;
/* u1_188 Output nets */
wire t_530,    t_531;
/* u2_189 Output nets */
wire t_532,    t_533,    t_534;
/* u2_190 Output nets */
wire t_535,    t_536,    t_537;
/* u2_191 Output nets */
wire t_538,    t_539,    t_540;
/* u2_192 Output nets */
wire t_541,    t_542,    t_543;
/* u2_193 Output nets */
wire t_544,    t_545,    t_546;
/* u2_194 Output nets */
wire t_547,    t_548,    t_549;
/* u1_195 Output nets */
wire t_550,    t_551;
/* u2_196 Output nets */
wire t_552,    t_553,    t_554;
/* u2_197 Output nets */
wire t_555,    t_556,    t_557;
/* u2_198 Output nets */
wire t_558,    t_559,    t_560;
/* u2_199 Output nets */
wire t_561,    t_562,    t_563;
/* u2_200 Output nets */
wire t_564,    t_565,    t_566;
/* u2_201 Output nets */
wire t_567,    t_568,    t_569;
/* u2_202 Output nets */
wire t_570,    t_571,    t_572;
/* u2_203 Output nets */
wire t_573,    t_574,    t_575;
/* u2_204 Output nets */
wire t_576,    t_577,    t_578;
/* u2_205 Output nets */
wire t_579,    t_580,    t_581;
/* u2_206 Output nets */
wire t_582,    t_583,    t_584;
/* u2_207 Output nets */
wire t_585,    t_586,    t_587;
/* u2_208 Output nets */
wire t_588,    t_589,    t_590;
/* u1_209 Output nets */
wire t_591,    t_592;
/* u2_210 Output nets */
wire t_593,    t_594,    t_595;
/* u2_211 Output nets */
wire t_596,    t_597,    t_598;
/* u2_212 Output nets */
wire t_599,    t_600,    t_601;
/* u2_213 Output nets */
wire t_602,    t_603,    t_604;
/* u2_214 Output nets */
wire t_605,    t_606,    t_607;
/* u2_215 Output nets */
wire t_608,    t_609,    t_610;
/* u2_216 Output nets */
wire t_611,    t_612,    t_613;
/* u2_217 Output nets */
wire t_614,    t_615,    t_616;
/* u2_218 Output nets */
wire t_617,    t_618,    t_619;
/* u2_219 Output nets */
wire t_620,    t_621,    t_622;
/* u2_220 Output nets */
wire t_623,    t_624,    t_625;
/* u2_221 Output nets */
wire t_626,    t_627,    t_628;
/* u2_222 Output nets */
wire t_629,    t_630,    t_631;
/* u2_223 Output nets */
wire t_632,    t_633,    t_634;
/* u2_224 Output nets */
wire t_635,    t_636,    t_637;
/* u2_225 Output nets */
wire t_638,    t_639,    t_640;
/* u2_226 Output nets */
wire t_641,    t_642,    t_643;
/* u2_227 Output nets */
wire t_644,    t_645,    t_646;
/* u2_228 Output nets */
wire t_647,    t_648,    t_649;
/* u2_229 Output nets */
wire t_650,    t_651,    t_652;
/* u2_230 Output nets */
wire t_653,    t_654,    t_655;
/* u0_231 Output nets */
wire t_656,    t_657;
/* u2_232 Output nets */
wire t_658,    t_659,    t_660;
/* u2_233 Output nets */
wire t_661,    t_662,    t_663;
/* u2_234 Output nets */
wire t_664,    t_665,    t_666;
/* u2_235 Output nets */
wire t_667,    t_668,    t_669;
/* u2_236 Output nets */
wire t_670,    t_671,    t_672;
/* u2_237 Output nets */
wire t_673,    t_674,    t_675;
/* u2_238 Output nets */
wire t_676,    t_677,    t_678;
/* u0_239 Output nets */
wire t_679,    t_680;
/* u2_240 Output nets */
wire t_681,    t_682,    t_683;
/* u2_241 Output nets */
wire t_684,    t_685,    t_686;
/* u2_242 Output nets */
wire t_687,    t_688,    t_689;
/* u2_243 Output nets */
wire t_690,    t_691,    t_692;
/* u2_244 Output nets */
wire t_693,    t_694,    t_695;
/* u2_245 Output nets */
wire t_696,    t_697,    t_698;
/* u2_246 Output nets */
wire t_699,    t_700,    t_701;
/* u1_247 Output nets */
wire t_702,    t_703;
/* u2_248 Output nets */
wire t_704,    t_705,    t_706;
/* u2_249 Output nets */
wire t_707,    t_708,    t_709;
/* u2_250 Output nets */
wire t_710,    t_711,    t_712;
/* u2_251 Output nets */
wire t_713,    t_714,    t_715;
/* u2_252 Output nets */
wire t_716,    t_717,    t_718;
/* u2_253 Output nets */
wire t_719,    t_720,    t_721;
/* u2_254 Output nets */
wire t_722,    t_723,    t_724;
/* u1_255 Output nets */
wire t_725,    t_726;
/* u2_256 Output nets */
wire t_727,    t_728,    t_729;
/* u2_257 Output nets */
wire t_730,    t_731,    t_732;
/* u2_258 Output nets */
wire t_733,    t_734,    t_735;
/* u2_259 Output nets */
wire t_736,    t_737,    t_738;
/* u2_260 Output nets */
wire t_739,    t_740,    t_741;
/* u2_261 Output nets */
wire t_742,    t_743,    t_744;
/* u2_262 Output nets */
wire t_745,    t_746,    t_747;
/* u2_263 Output nets */
wire t_748,    t_749,    t_750;
/* u2_264 Output nets */
wire t_751,    t_752,    t_753;
/* u2_265 Output nets */
wire t_754,    t_755,    t_756;
/* u2_266 Output nets */
wire t_757,    t_758,    t_759;
/* u2_267 Output nets */
wire t_760,    t_761,    t_762;
/* u2_268 Output nets */
wire t_763,    t_764,    t_765;
/* u2_269 Output nets */
wire t_766,    t_767,    t_768;
/* u2_270 Output nets */
wire t_769,    t_770,    t_771;
/* u1_271 Output nets */
wire t_772,    t_773;
/* u2_272 Output nets */
wire t_774,    t_775,    t_776;
/* u2_273 Output nets */
wire t_777,    t_778,    t_779;
/* u2_274 Output nets */
wire t_780,    t_781,    t_782;
/* u2_275 Output nets */
wire t_783,    t_784,    t_785;
/* u2_276 Output nets */
wire t_786,    t_787,    t_788;
/* u2_277 Output nets */
wire t_789,    t_790,    t_791;
/* u2_278 Output nets */
wire t_792,    t_793,    t_794;
/* u2_279 Output nets */
wire t_795,    t_796,    t_797;
/* u2_280 Output nets */
wire t_798,    t_799,    t_800;
/* u2_281 Output nets */
wire t_801,    t_802,    t_803;
/* u2_282 Output nets */
wire t_804,    t_805,    t_806;
/* u2_283 Output nets */
wire t_807,    t_808,    t_809;
/* u2_284 Output nets */
wire t_810,    t_811,    t_812;
/* u2_285 Output nets */
wire t_813,    t_814,    t_815;
/* u2_286 Output nets */
wire t_816,    t_817,    t_818;
/* u2_287 Output nets */
wire t_819,    t_820,    t_821;
/* u2_288 Output nets */
wire t_822,    t_823,    t_824;
/* u2_289 Output nets */
wire t_825,    t_826,    t_827;
/* u2_290 Output nets */
wire t_828,    t_829,    t_830;
/* u2_291 Output nets */
wire t_831,    t_832,    t_833;
/* u2_292 Output nets */
wire t_834,    t_835,    t_836;
/* u2_293 Output nets */
wire t_837,    t_838,    t_839;
/* u2_294 Output nets */
wire t_840,    t_841,    t_842;
/* u2_295 Output nets */
wire t_843,    t_844,    t_845;
/* u0_296 Output nets */
wire t_846,    t_847;
/* u2_297 Output nets */
wire t_848,    t_849,    t_850;
/* u2_298 Output nets */
wire t_851,    t_852,    t_853;
/* u2_299 Output nets */
wire t_854,    t_855,    t_856;
/* u2_300 Output nets */
wire t_857,    t_858,    t_859;
/* u2_301 Output nets */
wire t_860,    t_861,    t_862;
/* u2_302 Output nets */
wire t_863,    t_864,    t_865;
/* u2_303 Output nets */
wire t_866,    t_867,    t_868;
/* u2_304 Output nets */
wire t_869,    t_870,    t_871;
/* u0_305 Output nets */
wire t_872,    t_873;
/* u2_306 Output nets */
wire t_874,    t_875,    t_876;
/* u2_307 Output nets */
wire t_877,    t_878,    t_879;
/* u2_308 Output nets */
wire t_880,    t_881,    t_882;
/* u2_309 Output nets */
wire t_883,    t_884,    t_885;
/* u2_310 Output nets */
wire t_886,    t_887,    t_888;
/* u2_311 Output nets */
wire t_889,    t_890,    t_891;
/* u2_312 Output nets */
wire t_892,    t_893,    t_894;
/* u2_313 Output nets */
wire t_895,    t_896,    t_897;
/* u1_314 Output nets */
wire t_898,    t_899;
/* u2_315 Output nets */
wire t_900,    t_901,    t_902;
/* u2_316 Output nets */
wire t_903,    t_904,    t_905;
/* u2_317 Output nets */
wire t_906,    t_907,    t_908;
/* u2_318 Output nets */
wire t_909,    t_910,    t_911;
/* u2_319 Output nets */
wire t_912,    t_913,    t_914;
/* u2_320 Output nets */
wire t_915,    t_916,    t_917;
/* u2_321 Output nets */
wire t_918,    t_919,    t_920;
/* u2_322 Output nets */
wire t_921,    t_922,    t_923;
/* u1_323 Output nets */
wire t_924,    t_925;
/* u2_324 Output nets */
wire t_926,    t_927,    t_928;
/* u2_325 Output nets */
wire t_929,    t_930,    t_931;
/* u2_326 Output nets */
wire t_932,    t_933,    t_934;
/* u2_327 Output nets */
wire t_935,    t_936,    t_937;
/* u2_328 Output nets */
wire t_938,    t_939,    t_940;
/* u2_329 Output nets */
wire t_941,    t_942,    t_943;
/* u2_330 Output nets */
wire t_944,    t_945,    t_946;
/* u2_331 Output nets */
wire t_947,    t_948,    t_949;
/* u2_332 Output nets */
wire t_950,    t_951,    t_952;
/* u2_333 Output nets */
wire t_953,    t_954,    t_955;
/* u2_334 Output nets */
wire t_956,    t_957,    t_958;
/* u2_335 Output nets */
wire t_959,    t_960,    t_961;
/* u2_336 Output nets */
wire t_962,    t_963,    t_964;
/* u2_337 Output nets */
wire t_965,    t_966,    t_967;
/* u2_338 Output nets */
wire t_968,    t_969,    t_970;
/* u2_339 Output nets */
wire t_971,    t_972,    t_973;
/* u2_340 Output nets */
wire t_974,    t_975,    t_976;
/* u1_341 Output nets */
wire t_977,    t_978;
/* u2_342 Output nets */
wire t_979,    t_980,    t_981;
/* u2_343 Output nets */
wire t_982,    t_983,    t_984;
/* u2_344 Output nets */
wire t_985,    t_986,    t_987;
/* u2_345 Output nets */
wire t_988,    t_989,    t_990;
/* u2_346 Output nets */
wire t_991,    t_992,    t_993;
/* u2_347 Output nets */
wire t_994,    t_995,    t_996;
/* u2_348 Output nets */
wire t_997,    t_998,    t_999;
/* u2_349 Output nets */
wire t_1000,   t_1001,   t_1002;
/* u2_350 Output nets */
wire t_1003,   t_1004,   t_1005;
/* u2_351 Output nets */
wire t_1006,   t_1007,   t_1008;
/* u2_352 Output nets */
wire t_1009,   t_1010,   t_1011;
/* u2_353 Output nets */
wire t_1012,   t_1013,   t_1014;
/* u2_354 Output nets */
wire t_1015,   t_1016,   t_1017;
/* u2_355 Output nets */
wire t_1018,   t_1019,   t_1020;
/* u2_356 Output nets */
wire t_1021,   t_1022,   t_1023;
/* u2_357 Output nets */
wire t_1024,   t_1025,   t_1026;
/* u2_358 Output nets */
wire t_1027,   t_1028,   t_1029;
/* u2_359 Output nets */
wire t_1030,   t_1031,   t_1032;
/* u2_360 Output nets */
wire t_1033,   t_1034,   t_1035;
/* u2_361 Output nets */
wire t_1036,   t_1037,   t_1038;
/* u2_362 Output nets */
wire t_1039,   t_1040,   t_1041;
/* u2_363 Output nets */
wire t_1042,   t_1043,   t_1044;
/* u2_364 Output nets */
wire t_1045,   t_1046,   t_1047;
/* u2_365 Output nets */
wire t_1048,   t_1049,   t_1050;
/* u2_366 Output nets */
wire t_1051,   t_1052,   t_1053;
/* u2_367 Output nets */
wire t_1054,   t_1055,   t_1056;
/* u2_368 Output nets */
wire t_1057,   t_1058,   t_1059;
/* u0_369 Output nets */
wire t_1060,   t_1061;
/* u2_370 Output nets */
wire t_1062,   t_1063,   t_1064;
/* u2_371 Output nets */
wire t_1065,   t_1066,   t_1067;
/* u2_372 Output nets */
wire t_1068,   t_1069,   t_1070;
/* u2_373 Output nets */
wire t_1071,   t_1072,   t_1073;
/* u2_374 Output nets */
wire t_1074,   t_1075,   t_1076;
/* u2_375 Output nets */
wire t_1077,   t_1078,   t_1079;
/* u2_376 Output nets */
wire t_1080,   t_1081,   t_1082;
/* u2_377 Output nets */
wire t_1083,   t_1084,   t_1085;
/* u2_378 Output nets */
wire t_1086,   t_1087,   t_1088;
/* u0_379 Output nets */
wire t_1089,   t_1090;
/* u2_380 Output nets */
wire t_1091,   t_1092,   t_1093;
/* u2_381 Output nets */
wire t_1094,   t_1095,   t_1096;
/* u2_382 Output nets */
wire t_1097,   t_1098,   t_1099;
/* u2_383 Output nets */
wire t_1100,   t_1101,   t_1102;
/* u2_384 Output nets */
wire t_1103,   t_1104,   t_1105;
/* u2_385 Output nets */
wire t_1106,   t_1107,   t_1108;
/* u2_386 Output nets */
wire t_1109,   t_1110,   t_1111;
/* u2_387 Output nets */
wire t_1112,   t_1113,   t_1114;
/* u2_388 Output nets */
wire t_1115,   t_1116,   t_1117;
/* u1_389 Output nets */
wire t_1118,   t_1119;
/* u2_390 Output nets */
wire t_1120,   t_1121,   t_1122;
/* u2_391 Output nets */
wire t_1123,   t_1124,   t_1125;
/* u2_392 Output nets */
wire t_1126,   t_1127,   t_1128;
/* u2_393 Output nets */
wire t_1129,   t_1130,   t_1131;
/* u2_394 Output nets */
wire t_1132,   t_1133,   t_1134;
/* u2_395 Output nets */
wire t_1135,   t_1136,   t_1137;
/* u2_396 Output nets */
wire t_1138,   t_1139,   t_1140;
/* u2_397 Output nets */
wire t_1141,   t_1142,   t_1143;
/* u2_398 Output nets */
wire t_1144,   t_1145,   t_1146;
/* u1_399 Output nets */
wire t_1147,   t_1148;
/* u2_400 Output nets */
wire t_1149,   t_1150,   t_1151;
/* u2_401 Output nets */
wire t_1152,   t_1153,   t_1154;
/* u2_402 Output nets */
wire t_1155,   t_1156,   t_1157;
/* u2_403 Output nets */
wire t_1158,   t_1159,   t_1160;
/* u2_404 Output nets */
wire t_1161,   t_1162,   t_1163;
/* u2_405 Output nets */
wire t_1164,   t_1165,   t_1166;
/* u2_406 Output nets */
wire t_1167,   t_1168,   t_1169;
/* u2_407 Output nets */
wire t_1170,   t_1171,   t_1172;
/* u2_408 Output nets */
wire t_1173,   t_1174,   t_1175;
/* u2_409 Output nets */
wire t_1176,   t_1177,   t_1178;
/* u2_410 Output nets */
wire t_1179,   t_1180,   t_1181;
/* u2_411 Output nets */
wire t_1182,   t_1183,   t_1184;
/* u2_412 Output nets */
wire t_1185,   t_1186,   t_1187;
/* u2_413 Output nets */
wire t_1188,   t_1189,   t_1190;
/* u2_414 Output nets */
wire t_1191,   t_1192,   t_1193;
/* u2_415 Output nets */
wire t_1194,   t_1195,   t_1196;
/* u2_416 Output nets */
wire t_1197,   t_1198,   t_1199;
/* u2_417 Output nets */
wire t_1200,   t_1201,   t_1202;
/* u2_418 Output nets */
wire t_1203,   t_1204,   t_1205;
/* u1_419 Output nets */
wire t_1206,   t_1207;
/* u2_420 Output nets */
wire t_1208,   t_1209,   t_1210;
/* u2_421 Output nets */
wire t_1211,   t_1212,   t_1213;
/* u2_422 Output nets */
wire t_1214,   t_1215,   t_1216;
/* u2_423 Output nets */
wire t_1217,   t_1218,   t_1219;
/* u2_424 Output nets */
wire t_1220,   t_1221,   t_1222;
/* u2_425 Output nets */
wire t_1223,   t_1224,   t_1225;
/* u2_426 Output nets */
wire t_1226,   t_1227,   t_1228;
/* u2_427 Output nets */
wire t_1229,   t_1230,   t_1231;
/* u2_428 Output nets */
wire t_1232,   t_1233,   t_1234;
/* u2_429 Output nets */
wire t_1235,   t_1236,   t_1237;
/* u2_430 Output nets */
wire t_1238,   t_1239,   t_1240;
/* u2_431 Output nets */
wire t_1241,   t_1242,   t_1243;
/* u2_432 Output nets */
wire t_1244,   t_1245,   t_1246;
/* u2_433 Output nets */
wire t_1247,   t_1248,   t_1249;
/* u2_434 Output nets */
wire t_1250,   t_1251,   t_1252;
/* u2_435 Output nets */
wire t_1253,   t_1254,   t_1255;
/* u2_436 Output nets */
wire t_1256,   t_1257,   t_1258;
/* u2_437 Output nets */
wire t_1259,   t_1260,   t_1261;
/* u2_438 Output nets */
wire t_1262,   t_1263,   t_1264;
/* u2_439 Output nets */
wire t_1265,   t_1266,   t_1267;
/* u2_440 Output nets */
wire t_1268,   t_1269,   t_1270;
/* u2_441 Output nets */
wire t_1271,   t_1272,   t_1273;
/* u2_442 Output nets */
wire t_1274,   t_1275,   t_1276;
/* u2_443 Output nets */
wire t_1277,   t_1278,   t_1279;
/* u2_444 Output nets */
wire t_1280,   t_1281,   t_1282;
/* u2_445 Output nets */
wire t_1283,   t_1284,   t_1285;
/* u2_446 Output nets */
wire t_1286,   t_1287,   t_1288;
/* u2_447 Output nets */
wire t_1289,   t_1290,   t_1291;
/* u2_448 Output nets */
wire t_1292,   t_1293,   t_1294;
/* u2_449 Output nets */
wire t_1295,   t_1296,   t_1297;
/* u0_450 Output nets */
wire t_1298,   t_1299;
/* u2_451 Output nets */
wire t_1300,   t_1301,   t_1302;
/* u2_452 Output nets */
wire t_1303,   t_1304,   t_1305;
/* u2_453 Output nets */
wire t_1306,   t_1307,   t_1308;
/* u2_454 Output nets */
wire t_1309,   t_1310,   t_1311;
/* u2_455 Output nets */
wire t_1312,   t_1313,   t_1314;
/* u2_456 Output nets */
wire t_1315,   t_1316,   t_1317;
/* u2_457 Output nets */
wire t_1318,   t_1319,   t_1320;
/* u2_458 Output nets */
wire t_1321,   t_1322,   t_1323;
/* u2_459 Output nets */
wire t_1324,   t_1325,   t_1326;
/* u2_460 Output nets */
wire t_1327,   t_1328,   t_1329;
/* u0_461 Output nets */
wire t_1330,   t_1331;
/* u2_462 Output nets */
wire t_1332,   t_1333,   t_1334;
/* u2_463 Output nets */
wire t_1335,   t_1336,   t_1337;
/* u2_464 Output nets */
wire t_1338,   t_1339,   t_1340;
/* u2_465 Output nets */
wire t_1341,   t_1342,   t_1343;
/* u2_466 Output nets */
wire t_1344,   t_1345,   t_1346;
/* u2_467 Output nets */
wire t_1347,   t_1348,   t_1349;
/* u2_468 Output nets */
wire t_1350,   t_1351,   t_1352;
/* u2_469 Output nets */
wire t_1353,   t_1354,   t_1355;
/* u2_470 Output nets */
wire t_1356,   t_1357,   t_1358;
/* u2_471 Output nets */
wire t_1359,   t_1360,   t_1361;
/* u1_472 Output nets */
wire t_1362,   t_1363;
/* u2_473 Output nets */
wire t_1364,   t_1365,   t_1366;
/* u2_474 Output nets */
wire t_1367,   t_1368,   t_1369;
/* u2_475 Output nets */
wire t_1370,   t_1371,   t_1372;
/* u2_476 Output nets */
wire t_1373,   t_1374,   t_1375;
/* u2_477 Output nets */
wire t_1376,   t_1377,   t_1378;
/* u2_478 Output nets */
wire t_1379,   t_1380,   t_1381;
/* u2_479 Output nets */
wire t_1382,   t_1383,   t_1384;
/* u2_480 Output nets */
wire t_1385,   t_1386,   t_1387;
/* u2_481 Output nets */
wire t_1388,   t_1389,   t_1390;
/* u2_482 Output nets */
wire t_1391,   t_1392,   t_1393;
/* u1_483 Output nets */
wire t_1394,   t_1395;
/* u2_484 Output nets */
wire t_1396,   t_1397,   t_1398;
/* u2_485 Output nets */
wire t_1399,   t_1400,   t_1401;
/* u2_486 Output nets */
wire t_1402,   t_1403,   t_1404;
/* u2_487 Output nets */
wire t_1405,   t_1406,   t_1407;
/* u2_488 Output nets */
wire t_1408,   t_1409,   t_1410;
/* u2_489 Output nets */
wire t_1411,   t_1412,   t_1413;
/* u2_490 Output nets */
wire t_1414,   t_1415,   t_1416;
/* u2_491 Output nets */
wire t_1417,   t_1418,   t_1419;
/* u2_492 Output nets */
wire t_1420,   t_1421,   t_1422;
/* u2_493 Output nets */
wire t_1423,   t_1424,   t_1425;
/* u2_494 Output nets */
wire t_1426,   t_1427,   t_1428;
/* u2_495 Output nets */
wire t_1429,   t_1430,   t_1431;
/* u2_496 Output nets */
wire t_1432,   t_1433,   t_1434;
/* u2_497 Output nets */
wire t_1435,   t_1436,   t_1437;
/* u2_498 Output nets */
wire t_1438,   t_1439,   t_1440;
/* u2_499 Output nets */
wire t_1441,   t_1442,   t_1443;
/* u2_500 Output nets */
wire t_1444,   t_1445,   t_1446;
/* u2_501 Output nets */
wire t_1447,   t_1448,   t_1449;
/* u2_502 Output nets */
wire t_1450,   t_1451,   t_1452;
/* u2_503 Output nets */
wire t_1453,   t_1454,   t_1455;
/* u2_504 Output nets */
wire t_1456,   t_1457,   t_1458;
/* u1_505 Output nets */
wire t_1459,   t_1460;
/* u2_506 Output nets */
wire t_1461,   t_1462,   t_1463;
/* u2_507 Output nets */
wire t_1464,   t_1465,   t_1466;
/* u2_508 Output nets */
wire t_1467,   t_1468,   t_1469;
/* u2_509 Output nets */
wire t_1470,   t_1471,   t_1472;
/* u2_510 Output nets */
wire t_1473,   t_1474,   t_1475;
/* u2_511 Output nets */
wire t_1476,   t_1477,   t_1478;
/* u2_512 Output nets */
wire t_1479,   t_1480,   t_1481;
/* u2_513 Output nets */
wire t_1482,   t_1483,   t_1484;
/* u2_514 Output nets */
wire t_1485,   t_1486,   t_1487;
/* u2_515 Output nets */
wire t_1488,   t_1489,   t_1490;
/* u2_516 Output nets */
wire t_1491,   t_1492,   t_1493;
/* u2_517 Output nets */
wire t_1494,   t_1495,   t_1496;
/* u2_518 Output nets */
wire t_1497,   t_1498,   t_1499;
/* u2_519 Output nets */
wire t_1500,   t_1501,   t_1502;
/* u2_520 Output nets */
wire t_1503,   t_1504,   t_1505;
/* u2_521 Output nets */
wire t_1506,   t_1507,   t_1508;
/* u2_522 Output nets */
wire t_1509,   t_1510,   t_1511;
/* u2_523 Output nets */
wire t_1512,   t_1513,   t_1514;
/* u2_524 Output nets */
wire t_1515,   t_1516,   t_1517;
/* u2_525 Output nets */
wire t_1518,   t_1519,   t_1520;
/* u2_526 Output nets */
wire t_1521,   t_1522,   t_1523;
/* u2_527 Output nets */
wire t_1524,   t_1525,   t_1526;
/* u2_528 Output nets */
wire t_1527,   t_1528,   t_1529;
/* u2_529 Output nets */
wire t_1530,   t_1531,   t_1532;
/* u2_530 Output nets */
wire t_1533,   t_1534,   t_1535;
/* u2_531 Output nets */
wire t_1536,   t_1537,   t_1538;
/* u2_532 Output nets */
wire t_1539,   t_1540,   t_1541;
/* u2_533 Output nets */
wire t_1542,   t_1543,   t_1544;
/* u2_534 Output nets */
wire t_1545,   t_1546,   t_1547;
/* u2_535 Output nets */
wire t_1548,   t_1549,   t_1550;
/* u2_536 Output nets */
wire t_1551,   t_1552,   t_1553;
/* u2_537 Output nets */
wire t_1554,   t_1555,   t_1556;
/* u2_538 Output nets */
wire t_1557,   t_1558,   t_1559;
/* u0_539 Output nets */
wire t_1560,   t_1561;
/* u2_540 Output nets */
wire t_1562,   t_1563,   t_1564;
/* u2_541 Output nets */
wire t_1565,   t_1566,   t_1567;
/* u2_542 Output nets */
wire t_1568,   t_1569,   t_1570;
/* u2_543 Output nets */
wire t_1571,   t_1572,   t_1573;
/* u2_544 Output nets */
wire t_1574,   t_1575,   t_1576;
/* u2_545 Output nets */
wire t_1577,   t_1578,   t_1579;
/* u2_546 Output nets */
wire t_1580,   t_1581,   t_1582;
/* u2_547 Output nets */
wire t_1583,   t_1584,   t_1585;
/* u2_548 Output nets */
wire t_1586,   t_1587,   t_1588;
/* u2_549 Output nets */
wire t_1589,   t_1590,   t_1591;
/* u2_550 Output nets */
wire t_1592,   t_1593,   t_1594;
/* u0_551 Output nets */
wire t_1595,   t_1596;
/* u2_552 Output nets */
wire t_1597,   t_1598,   t_1599;
/* u2_553 Output nets */
wire t_1600,   t_1601,   t_1602;
/* u2_554 Output nets */
wire t_1603,   t_1604,   t_1605;
/* u2_555 Output nets */
wire t_1606,   t_1607,   t_1608;
/* u2_556 Output nets */
wire t_1609,   t_1610,   t_1611;
/* u2_557 Output nets */
wire t_1612,   t_1613,   t_1614;
/* u2_558 Output nets */
wire t_1615,   t_1616,   t_1617;
/* u2_559 Output nets */
wire t_1618,   t_1619,   t_1620;
/* u2_560 Output nets */
wire t_1621,   t_1622,   t_1623;
/* u2_561 Output nets */
wire t_1624,   t_1625,   t_1626;
/* u2_562 Output nets */
wire t_1627,   t_1628,   t_1629;
/* u1_563 Output nets */
wire t_1630,   t_1631;
/* u2_564 Output nets */
wire t_1632,   t_1633,   t_1634;
/* u2_565 Output nets */
wire t_1635,   t_1636,   t_1637;
/* u2_566 Output nets */
wire t_1638,   t_1639,   t_1640;
/* u2_567 Output nets */
wire t_1641,   t_1642,   t_1643;
/* u2_568 Output nets */
wire t_1644,   t_1645,   t_1646;
/* u2_569 Output nets */
wire t_1647,   t_1648,   t_1649;
/* u2_570 Output nets */
wire t_1650,   t_1651,   t_1652;
/* u2_571 Output nets */
wire t_1653,   t_1654,   t_1655;
/* u2_572 Output nets */
wire t_1656,   t_1657,   t_1658;
/* u2_573 Output nets */
wire t_1659,   t_1660,   t_1661;
/* u2_574 Output nets */
wire t_1662,   t_1663,   t_1664;
/* u1_575 Output nets */
wire t_1665,   t_1666;
/* u2_576 Output nets */
wire t_1667,   t_1668,   t_1669;
/* u2_577 Output nets */
wire t_1670,   t_1671,   t_1672;
/* u2_578 Output nets */
wire t_1673,   t_1674,   t_1675;
/* u2_579 Output nets */
wire t_1676,   t_1677,   t_1678;
/* u2_580 Output nets */
wire t_1679,   t_1680,   t_1681;
/* u2_581 Output nets */
wire t_1682,   t_1683,   t_1684;
/* u2_582 Output nets */
wire t_1685,   t_1686,   t_1687;
/* u2_583 Output nets */
wire t_1688,   t_1689,   t_1690;
/* u2_584 Output nets */
wire t_1691,   t_1692,   t_1693;
/* u2_585 Output nets */
wire t_1694,   t_1695,   t_1696;
/* u2_586 Output nets */
wire t_1697,   t_1698,   t_1699;
/* u2_587 Output nets */
wire t_1700,   t_1701,   t_1702;
/* u2_588 Output nets */
wire t_1703,   t_1704,   t_1705;
/* u2_589 Output nets */
wire t_1706,   t_1707,   t_1708;
/* u2_590 Output nets */
wire t_1709,   t_1710,   t_1711;
/* u2_591 Output nets */
wire t_1712,   t_1713,   t_1714;
/* u2_592 Output nets */
wire t_1715,   t_1716,   t_1717;
/* u2_593 Output nets */
wire t_1718,   t_1719,   t_1720;
/* u2_594 Output nets */
wire t_1721,   t_1722,   t_1723;
/* u2_595 Output nets */
wire t_1724,   t_1725,   t_1726;
/* u2_596 Output nets */
wire t_1727,   t_1728,   t_1729;
/* u2_597 Output nets */
wire t_1730,   t_1731,   t_1732;
/* u2_598 Output nets */
wire t_1733,   t_1734,   t_1735;
/* u1_599 Output nets */
wire t_1736,   t_1737;
/* u2_600 Output nets */
wire t_1738,   t_1739,   t_1740;
/* u2_601 Output nets */
wire t_1741,   t_1742,   t_1743;
/* u2_602 Output nets */
wire t_1744,   t_1745,   t_1746;
/* u2_603 Output nets */
wire t_1747,   t_1748,   t_1749;
/* u2_604 Output nets */
wire t_1750,   t_1751,   t_1752;
/* u2_605 Output nets */
wire t_1753,   t_1754,   t_1755;
/* u2_606 Output nets */
wire t_1756,   t_1757,   t_1758;
/* u2_607 Output nets */
wire t_1759,   t_1760,   t_1761;
/* u2_608 Output nets */
wire t_1762,   t_1763,   t_1764;
/* u2_609 Output nets */
wire t_1765,   t_1766,   t_1767;
/* u2_610 Output nets */
wire t_1768,   t_1769,   t_1770;
/* u2_611 Output nets */
wire t_1771,   t_1772,   t_1773;
/* u2_612 Output nets */
wire t_1774,   t_1775,   t_1776;
/* u2_613 Output nets */
wire t_1777,   t_1778,   t_1779;
/* u2_614 Output nets */
wire t_1780,   t_1781,   t_1782;
/* u2_615 Output nets */
wire t_1783,   t_1784,   t_1785;
/* u2_616 Output nets */
wire t_1786,   t_1787,   t_1788;
/* u2_617 Output nets */
wire t_1789,   t_1790,   t_1791;
/* u2_618 Output nets */
wire t_1792,   t_1793,   t_1794;
/* u2_619 Output nets */
wire t_1795,   t_1796,   t_1797;
/* u2_620 Output nets */
wire t_1798,   t_1799,   t_1800;
/* u2_621 Output nets */
wire t_1801,   t_1802,   t_1803;
/* u2_622 Output nets */
wire t_1804,   t_1805,   t_1806;
/* u2_623 Output nets */
wire t_1807,   t_1808,   t_1809;
/* u2_624 Output nets */
wire t_1810,   t_1811,   t_1812;
/* u2_625 Output nets */
wire t_1813,   t_1814,   t_1815;
/* u2_626 Output nets */
wire t_1816,   t_1817,   t_1818;
/* u2_627 Output nets */
wire t_1819,   t_1820,   t_1821;
/* u2_628 Output nets */
wire t_1822,   t_1823,   t_1824;
/* u2_629 Output nets */
wire t_1825,   t_1826,   t_1827;
/* u2_630 Output nets */
wire t_1828,   t_1829,   t_1830;
/* u2_631 Output nets */
wire t_1831,   t_1832,   t_1833;
/* u2_632 Output nets */
wire t_1834,   t_1835,   t_1836;
/* u2_633 Output nets */
wire t_1837,   t_1838,   t_1839;
/* u2_634 Output nets */
wire t_1840,   t_1841,   t_1842;
/* u2_635 Output nets */
wire t_1843,   t_1844,   t_1845;
/* u0_636 Output nets */
wire t_1846,   t_1847;
/* u2_637 Output nets */
wire t_1848,   t_1849,   t_1850;
/* u2_638 Output nets */
wire t_1851,   t_1852,   t_1853;
/* u2_639 Output nets */
wire t_1854,   t_1855,   t_1856;
/* u2_640 Output nets */
wire t_1857,   t_1858,   t_1859;
/* u2_641 Output nets */
wire t_1860,   t_1861,   t_1862;
/* u2_642 Output nets */
wire t_1863,   t_1864,   t_1865;
/* u2_643 Output nets */
wire t_1866,   t_1867,   t_1868;
/* u2_644 Output nets */
wire t_1869,   t_1870,   t_1871;
/* u2_645 Output nets */
wire t_1872,   t_1873,   t_1874;
/* u2_646 Output nets */
wire t_1875,   t_1876,   t_1877;
/* u2_647 Output nets */
wire t_1878,   t_1879,   t_1880;
/* u2_648 Output nets */
wire t_1881,   t_1882,   t_1883;
/* u0_649 Output nets */
wire t_1884,   t_1885;
/* u2_650 Output nets */
wire t_1886,   t_1887,   t_1888;
/* u2_651 Output nets */
wire t_1889,   t_1890,   t_1891;
/* u2_652 Output nets */
wire t_1892,   t_1893,   t_1894;
/* u2_653 Output nets */
wire t_1895,   t_1896,   t_1897;
/* u2_654 Output nets */
wire t_1898,   t_1899,   t_1900;
/* u2_655 Output nets */
wire t_1901,   t_1902,   t_1903;
/* u2_656 Output nets */
wire t_1904,   t_1905,   t_1906;
/* u2_657 Output nets */
wire t_1907,   t_1908,   t_1909;
/* u2_658 Output nets */
wire t_1910,   t_1911,   t_1912;
/* u2_659 Output nets */
wire t_1913,   t_1914,   t_1915;
/* u2_660 Output nets */
wire t_1916,   t_1917,   t_1918;
/* u2_661 Output nets */
wire t_1919,   t_1920,   t_1921;
/* u1_662 Output nets */
wire t_1922,   t_1923;
/* u2_663 Output nets */
wire t_1924,   t_1925,   t_1926;
/* u2_664 Output nets */
wire t_1927,   t_1928,   t_1929;
/* u2_665 Output nets */
wire t_1930,   t_1931,   t_1932;
/* u2_666 Output nets */
wire t_1933,   t_1934,   t_1935;
/* u2_667 Output nets */
wire t_1936,   t_1937,   t_1938;
/* u2_668 Output nets */
wire t_1939,   t_1940,   t_1941;
/* u2_669 Output nets */
wire t_1942,   t_1943,   t_1944;
/* u2_670 Output nets */
wire t_1945,   t_1946,   t_1947;
/* u2_671 Output nets */
wire t_1948,   t_1949,   t_1950;
/* u2_672 Output nets */
wire t_1951,   t_1952,   t_1953;
/* u2_673 Output nets */
wire t_1954,   t_1955,   t_1956;
/* u2_674 Output nets */
wire t_1957,   t_1958,   t_1959;
/* u1_675 Output nets */
wire t_1960,   t_1961;
/* u2_676 Output nets */
wire t_1962,   t_1963,   t_1964;
/* u2_677 Output nets */
wire t_1965,   t_1966,   t_1967;
/* u2_678 Output nets */
wire t_1968,   t_1969,   t_1970;
/* u2_679 Output nets */
wire t_1971,   t_1972,   t_1973;
/* u2_680 Output nets */
wire t_1974,   t_1975,   t_1976;
/* u2_681 Output nets */
wire t_1977,   t_1978,   t_1979;
/* u2_682 Output nets */
wire t_1980,   t_1981,   t_1982;
/* u2_683 Output nets */
wire t_1983,   t_1984,   t_1985;
/* u2_684 Output nets */
wire t_1986,   t_1987,   t_1988;
/* u2_685 Output nets */
wire t_1989,   t_1990,   t_1991;
/* u2_686 Output nets */
wire t_1992,   t_1993,   t_1994;
/* u2_687 Output nets */
wire t_1995,   t_1996,   t_1997;
/* u2_688 Output nets */
wire t_1998,   t_1999,   t_2000;
/* u2_689 Output nets */
wire t_2001,   t_2002,   t_2003;
/* u2_690 Output nets */
wire t_2004,   t_2005,   t_2006;
/* u2_691 Output nets */
wire t_2007,   t_2008,   t_2009;
/* u2_692 Output nets */
wire t_2010,   t_2011,   t_2012;
/* u2_693 Output nets */
wire t_2013,   t_2014,   t_2015;
/* u2_694 Output nets */
wire t_2016,   t_2017,   t_2018;
/* u2_695 Output nets */
wire t_2019,   t_2020,   t_2021;
/* u2_696 Output nets */
wire t_2022,   t_2023,   t_2024;
/* u2_697 Output nets */
wire t_2025,   t_2026,   t_2027;
/* u2_698 Output nets */
wire t_2028,   t_2029,   t_2030;
/* u2_699 Output nets */
wire t_2031,   t_2032,   t_2033;
/* u2_700 Output nets */
wire t_2034,   t_2035,   t_2036;
/* u1_701 Output nets */
wire t_2037,   t_2038;
/* u2_702 Output nets */
wire t_2039,   t_2040,   t_2041;
/* u2_703 Output nets */
wire t_2042,   t_2043,   t_2044;
/* u2_704 Output nets */
wire t_2045,   t_2046,   t_2047;
/* u2_705 Output nets */
wire t_2048,   t_2049,   t_2050;
/* u2_706 Output nets */
wire t_2051,   t_2052,   t_2053;
/* u2_707 Output nets */
wire t_2054,   t_2055,   t_2056;
/* u2_708 Output nets */
wire t_2057,   t_2058,   t_2059;
/* u2_709 Output nets */
wire t_2060,   t_2061,   t_2062;
/* u2_710 Output nets */
wire t_2063,   t_2064,   t_2065;
/* u2_711 Output nets */
wire t_2066,   t_2067,   t_2068;
/* u2_712 Output nets */
wire t_2069,   t_2070,   t_2071;
/* u2_713 Output nets */
wire t_2072,   t_2073,   t_2074;
/* u2_714 Output nets */
wire t_2075,   t_2076,   t_2077;
/* u2_715 Output nets */
wire t_2078,   t_2079,   t_2080;
/* u2_716 Output nets */
wire t_2081,   t_2082,   t_2083;
/* u2_717 Output nets */
wire t_2084,   t_2085,   t_2086;
/* u2_718 Output nets */
wire t_2087,   t_2088,   t_2089;
/* u2_719 Output nets */
wire t_2090,   t_2091,   t_2092;
/* u2_720 Output nets */
wire t_2093,   t_2094,   t_2095;
/* u2_721 Output nets */
wire t_2096,   t_2097,   t_2098;
/* u2_722 Output nets */
wire t_2099,   t_2100,   t_2101;
/* u2_723 Output nets */
wire t_2102,   t_2103,   t_2104;
/* u2_724 Output nets */
wire t_2105,   t_2106,   t_2107;
/* u2_725 Output nets */
wire t_2108,   t_2109,   t_2110;
/* u2_726 Output nets */
wire t_2111,   t_2112,   t_2113;
/* u2_727 Output nets */
wire t_2114,   t_2115,   t_2116;
/* u2_728 Output nets */
wire t_2117,   t_2118,   t_2119;
/* u2_729 Output nets */
wire t_2120,   t_2121,   t_2122;
/* u2_730 Output nets */
wire t_2123,   t_2124,   t_2125;
/* u2_731 Output nets */
wire t_2126,   t_2127,   t_2128;
/* u2_732 Output nets */
wire t_2129,   t_2130,   t_2131;
/* u2_733 Output nets */
wire t_2132,   t_2133,   t_2134;
/* u2_734 Output nets */
wire t_2135,   t_2136,   t_2137;
/* u2_735 Output nets */
wire t_2138,   t_2139,   t_2140;
/* u2_736 Output nets */
wire t_2141,   t_2142,   t_2143;
/* u2_737 Output nets */
wire t_2144,   t_2145,   t_2146;
/* u2_738 Output nets */
wire t_2147,   t_2148,   t_2149;
/* u2_739 Output nets */
wire t_2150,   t_2151,   t_2152;
/* u2_740 Output nets */
wire t_2153,   t_2154,   t_2155;
/* u0_741 Output nets */
wire t_2156,   t_2157;
/* u2_742 Output nets */
wire t_2158,   t_2159,   t_2160;
/* u2_743 Output nets */
wire t_2161,   t_2162,   t_2163;
/* u2_744 Output nets */
wire t_2164,   t_2165,   t_2166;
/* u2_745 Output nets */
wire t_2167,   t_2168,   t_2169;
/* u2_746 Output nets */
wire t_2170,   t_2171,   t_2172;
/* u2_747 Output nets */
wire t_2173,   t_2174,   t_2175;
/* u2_748 Output nets */
wire t_2176,   t_2177,   t_2178;
/* u2_749 Output nets */
wire t_2179,   t_2180,   t_2181;
/* u2_750 Output nets */
wire t_2182,   t_2183,   t_2184;
/* u2_751 Output nets */
wire t_2185,   t_2186,   t_2187;
/* u2_752 Output nets */
wire t_2188,   t_2189,   t_2190;
/* u2_753 Output nets */
wire t_2191,   t_2192,   t_2193;
/* u2_754 Output nets */
wire t_2194,   t_2195,   t_2196;
/* u0_755 Output nets */
wire t_2197,   t_2198;
/* u2_756 Output nets */
wire t_2199,   t_2200,   t_2201;
/* u2_757 Output nets */
wire t_2202,   t_2203,   t_2204;
/* u2_758 Output nets */
wire t_2205,   t_2206,   t_2207;
/* u2_759 Output nets */
wire t_2208,   t_2209,   t_2210;
/* u2_760 Output nets */
wire t_2211,   t_2212,   t_2213;
/* u2_761 Output nets */
wire t_2214,   t_2215,   t_2216;
/* u2_762 Output nets */
wire t_2217,   t_2218,   t_2219;
/* u2_763 Output nets */
wire t_2220,   t_2221,   t_2222;
/* u2_764 Output nets */
wire t_2223,   t_2224,   t_2225;
/* u2_765 Output nets */
wire t_2226,   t_2227,   t_2228;
/* u2_766 Output nets */
wire t_2229,   t_2230,   t_2231;
/* u2_767 Output nets */
wire t_2232,   t_2233,   t_2234;
/* u2_768 Output nets */
wire t_2235,   t_2236,   t_2237;
/* u1_769 Output nets */
wire t_2238,   t_2239;
/* u2_770 Output nets */
wire t_2240,   t_2241,   t_2242;
/* u2_771 Output nets */
wire t_2243,   t_2244,   t_2245;
/* u2_772 Output nets */
wire t_2246,   t_2247,   t_2248;
/* u2_773 Output nets */
wire t_2249,   t_2250,   t_2251;
/* u2_774 Output nets */
wire t_2252,   t_2253,   t_2254;
/* u2_775 Output nets */
wire t_2255,   t_2256,   t_2257;
/* u2_776 Output nets */
wire t_2258,   t_2259,   t_2260;
/* u2_777 Output nets */
wire t_2261,   t_2262,   t_2263;
/* u2_778 Output nets */
wire t_2264,   t_2265,   t_2266;
/* u2_779 Output nets */
wire t_2267,   t_2268,   t_2269;
/* u2_780 Output nets */
wire t_2270,   t_2271,   t_2272;
/* u2_781 Output nets */
wire t_2273,   t_2274,   t_2275;
/* u2_782 Output nets */
wire t_2276,   t_2277,   t_2278;
/* u1_783 Output nets */
wire t_2279,   t_2280;
/* u2_784 Output nets */
wire t_2281,   t_2282,   t_2283;
/* u2_785 Output nets */
wire t_2284,   t_2285,   t_2286;
/* u2_786 Output nets */
wire t_2287,   t_2288,   t_2289;
/* u2_787 Output nets */
wire t_2290,   t_2291,   t_2292;
/* u2_788 Output nets */
wire t_2293,   t_2294,   t_2295;
/* u2_789 Output nets */
wire t_2296,   t_2297,   t_2298;
/* u2_790 Output nets */
wire t_2299,   t_2300,   t_2301;
/* u2_791 Output nets */
wire t_2302,   t_2303,   t_2304;
/* u2_792 Output nets */
wire t_2305,   t_2306,   t_2307;
/* u2_793 Output nets */
wire t_2308,   t_2309,   t_2310;
/* u2_794 Output nets */
wire t_2311,   t_2312,   t_2313;
/* u2_795 Output nets */
wire t_2314,   t_2315,   t_2316;
/* u2_796 Output nets */
wire t_2317,   t_2318,   t_2319;
/* u2_797 Output nets */
wire t_2320,   t_2321,   t_2322;
/* u2_798 Output nets */
wire t_2323,   t_2324,   t_2325;
/* u2_799 Output nets */
wire t_2326,   t_2327,   t_2328;
/* u2_800 Output nets */
wire t_2329,   t_2330,   t_2331;
/* u2_801 Output nets */
wire t_2332,   t_2333,   t_2334;
/* u2_802 Output nets */
wire t_2335,   t_2336,   t_2337;
/* u2_803 Output nets */
wire t_2338,   t_2339,   t_2340;
/* u2_804 Output nets */
wire t_2341,   t_2342,   t_2343;
/* u2_805 Output nets */
wire t_2344,   t_2345,   t_2346;
/* u2_806 Output nets */
wire t_2347,   t_2348,   t_2349;
/* u2_807 Output nets */
wire t_2350,   t_2351,   t_2352;
/* u2_808 Output nets */
wire t_2353,   t_2354,   t_2355;
/* u2_809 Output nets */
wire t_2356,   t_2357,   t_2358;
/* u2_810 Output nets */
wire t_2359,   t_2360,   t_2361;
/* u1_811 Output nets */
wire t_2362,   t_2363;
/* u2_812 Output nets */
wire t_2364,   t_2365,   t_2366;
/* u2_813 Output nets */
wire t_2367,   t_2368,   t_2369;
/* u2_814 Output nets */
wire t_2370,   t_2371,   t_2372;
/* u2_815 Output nets */
wire t_2373,   t_2374,   t_2375;
/* u2_816 Output nets */
wire t_2376,   t_2377,   t_2378;
/* u2_817 Output nets */
wire t_2379,   t_2380,   t_2381;
/* u2_818 Output nets */
wire t_2382,   t_2383,   t_2384;
/* u2_819 Output nets */
wire t_2385,   t_2386,   t_2387;
/* u2_820 Output nets */
wire t_2388,   t_2389,   t_2390;
/* u2_821 Output nets */
wire t_2391,   t_2392,   t_2393;
/* u2_822 Output nets */
wire t_2394,   t_2395,   t_2396;
/* u2_823 Output nets */
wire t_2397,   t_2398,   t_2399;
/* u2_824 Output nets */
wire t_2400,   t_2401,   t_2402;
/* u2_825 Output nets */
wire t_2403,   t_2404,   t_2405;
/* u2_826 Output nets */
wire t_2406,   t_2407,   t_2408;
/* u2_827 Output nets */
wire t_2409,   t_2410,   t_2411;
/* u2_828 Output nets */
wire t_2412,   t_2413,   t_2414;
/* u2_829 Output nets */
wire t_2415,   t_2416,   t_2417;
/* u2_830 Output nets */
wire t_2418,   t_2419,   t_2420;
/* u2_831 Output nets */
wire t_2421,   t_2422,   t_2423;
/* u2_832 Output nets */
wire t_2424,   t_2425,   t_2426;
/* u2_833 Output nets */
wire t_2427,   t_2428,   t_2429;
/* u2_834 Output nets */
wire t_2430,   t_2431,   t_2432;
/* u2_835 Output nets */
wire t_2433,   t_2434,   t_2435;
/* u2_836 Output nets */
wire t_2436,   t_2437,   t_2438;
/* u2_837 Output nets */
wire t_2439,   t_2440,   t_2441;
/* u2_838 Output nets */
wire t_2442,   t_2443,   t_2444;
/* u2_839 Output nets */
wire t_2445,   t_2446,   t_2447;
/* u2_840 Output nets */
wire t_2448,   t_2449,   t_2450;
/* u2_841 Output nets */
wire t_2451,   t_2452,   t_2453;
/* u2_842 Output nets */
wire t_2454,   t_2455,   t_2456;
/* u2_843 Output nets */
wire t_2457,   t_2458,   t_2459;
/* u2_844 Output nets */
wire t_2460,   t_2461,   t_2462;
/* u2_845 Output nets */
wire t_2463,   t_2464,   t_2465;
/* u2_846 Output nets */
wire t_2466,   t_2467,   t_2468;
/* u2_847 Output nets */
wire t_2469,   t_2470,   t_2471;
/* u2_848 Output nets */
wire t_2472,   t_2473,   t_2474;
/* u2_849 Output nets */
wire t_2475,   t_2476,   t_2477;
/* u2_850 Output nets */
wire t_2478,   t_2479,   t_2480;
/* u2_851 Output nets */
wire t_2481,   t_2482,   t_2483;
/* u2_852 Output nets */
wire t_2484,   t_2485,   t_2486;
/* u2_853 Output nets */
wire t_2487,   t_2488,   t_2489;
/* u0_854 Output nets */
wire t_2490,   t_2491;
/* u2_855 Output nets */
wire t_2492,   t_2493,   t_2494;
/* u2_856 Output nets */
wire t_2495,   t_2496,   t_2497;
/* u2_857 Output nets */
wire t_2498,   t_2499,   t_2500;
/* u2_858 Output nets */
wire t_2501,   t_2502,   t_2503;
/* u2_859 Output nets */
wire t_2504,   t_2505,   t_2506;
/* u2_860 Output nets */
wire t_2507,   t_2508,   t_2509;
/* u2_861 Output nets */
wire t_2510,   t_2511,   t_2512;
/* u2_862 Output nets */
wire t_2513,   t_2514,   t_2515;
/* u2_863 Output nets */
wire t_2516,   t_2517,   t_2518;
/* u2_864 Output nets */
wire t_2519,   t_2520,   t_2521;
/* u2_865 Output nets */
wire t_2522,   t_2523,   t_2524;
/* u2_866 Output nets */
wire t_2525,   t_2526,   t_2527;
/* u2_867 Output nets */
wire t_2528,   t_2529,   t_2530;
/* u2_868 Output nets */
wire t_2531,   t_2532,   t_2533;
/* u0_869 Output nets */
wire t_2534,   t_2535;
/* u2_870 Output nets */
wire t_2536,   t_2537,   t_2538;
/* u2_871 Output nets */
wire t_2539,   t_2540,   t_2541;
/* u2_872 Output nets */
wire t_2542,   t_2543,   t_2544;
/* u2_873 Output nets */
wire t_2545,   t_2546,   t_2547;
/* u2_874 Output nets */
wire t_2548,   t_2549,   t_2550;
/* u2_875 Output nets */
wire t_2551,   t_2552,   t_2553;
/* u2_876 Output nets */
wire t_2554,   t_2555,   t_2556;
/* u2_877 Output nets */
wire t_2557,   t_2558,   t_2559;
/* u2_878 Output nets */
wire t_2560,   t_2561,   t_2562;
/* u2_879 Output nets */
wire t_2563,   t_2564,   t_2565;
/* u2_880 Output nets */
wire t_2566,   t_2567,   t_2568;
/* u2_881 Output nets */
wire t_2569,   t_2570,   t_2571;
/* u2_882 Output nets */
wire t_2572,   t_2573,   t_2574;
/* u2_883 Output nets */
wire t_2575,   t_2576,   t_2577;
/* u1_884 Output nets */
wire t_2578,   t_2579;
/* u2_885 Output nets */
wire t_2580,   t_2581,   t_2582;
/* u2_886 Output nets */
wire t_2583,   t_2584,   t_2585;
/* u2_887 Output nets */
wire t_2586,   t_2587,   t_2588;
/* u2_888 Output nets */
wire t_2589,   t_2590,   t_2591;
/* u2_889 Output nets */
wire t_2592,   t_2593,   t_2594;
/* u2_890 Output nets */
wire t_2595,   t_2596,   t_2597;
/* u2_891 Output nets */
wire t_2598,   t_2599,   t_2600;
/* u2_892 Output nets */
wire t_2601,   t_2602,   t_2603;
/* u2_893 Output nets */
wire t_2604,   t_2605,   t_2606;
/* u2_894 Output nets */
wire t_2607,   t_2608,   t_2609;
/* u2_895 Output nets */
wire t_2610,   t_2611,   t_2612;
/* u2_896 Output nets */
wire t_2613,   t_2614,   t_2615;
/* u2_897 Output nets */
wire t_2616,   t_2617,   t_2618;
/* u2_898 Output nets */
wire t_2619,   t_2620,   t_2621;
/* u1_899 Output nets */
wire t_2622,   t_2623;
/* u2_900 Output nets */
wire t_2624,   t_2625,   t_2626;
/* u2_901 Output nets */
wire t_2627,   t_2628,   t_2629;
/* u2_902 Output nets */
wire t_2630,   t_2631,   t_2632;
/* u2_903 Output nets */
wire t_2633,   t_2634,   t_2635;
/* u2_904 Output nets */
wire t_2636,   t_2637,   t_2638;
/* u2_905 Output nets */
wire t_2639,   t_2640,   t_2641;
/* u2_906 Output nets */
wire t_2642,   t_2643,   t_2644;
/* u2_907 Output nets */
wire t_2645,   t_2646,   t_2647;
/* u2_908 Output nets */
wire t_2648,   t_2649,   t_2650;
/* u2_909 Output nets */
wire t_2651,   t_2652,   t_2653;
/* u2_910 Output nets */
wire t_2654,   t_2655,   t_2656;
/* u2_911 Output nets */
wire t_2657,   t_2658,   t_2659;
/* u2_912 Output nets */
wire t_2660,   t_2661,   t_2662;
/* u2_913 Output nets */
wire t_2663,   t_2664,   t_2665;
/* u2_914 Output nets */
wire t_2666,   t_2667,   t_2668;
/* u2_915 Output nets */
wire t_2669,   t_2670,   t_2671;
/* u2_916 Output nets */
wire t_2672,   t_2673,   t_2674;
/* u2_917 Output nets */
wire t_2675,   t_2676,   t_2677;
/* u2_918 Output nets */
wire t_2678,   t_2679,   t_2680;
/* u2_919 Output nets */
wire t_2681,   t_2682,   t_2683;
/* u2_920 Output nets */
wire t_2684,   t_2685,   t_2686;
/* u2_921 Output nets */
wire t_2687,   t_2688,   t_2689;
/* u2_922 Output nets */
wire t_2690,   t_2691,   t_2692;
/* u2_923 Output nets */
wire t_2693,   t_2694,   t_2695;
/* u2_924 Output nets */
wire t_2696,   t_2697,   t_2698;
/* u2_925 Output nets */
wire t_2699,   t_2700,   t_2701;
/* u2_926 Output nets */
wire t_2702,   t_2703,   t_2704;
/* u2_927 Output nets */
wire t_2705,   t_2706,   t_2707;
/* u2_928 Output nets */
wire t_2708,   t_2709,   t_2710;
/* u1_929 Output nets */
wire t_2711,   t_2712;
/* u2_930 Output nets */
wire t_2713,   t_2714,   t_2715;
/* u2_931 Output nets */
wire t_2716,   t_2717,   t_2718;
/* u2_932 Output nets */
wire t_2719,   t_2720,   t_2721;
/* u2_933 Output nets */
wire t_2722,   t_2723,   t_2724;
/* u2_934 Output nets */
wire t_2725,   t_2726,   t_2727;
/* u2_935 Output nets */
wire t_2728,   t_2729,   t_2730;
/* u2_936 Output nets */
wire t_2731,   t_2732,   t_2733;
/* u2_937 Output nets */
wire t_2734,   t_2735,   t_2736;
/* u2_938 Output nets */
wire t_2737,   t_2738,   t_2739;
/* u2_939 Output nets */
wire t_2740,   t_2741,   t_2742;
/* u2_940 Output nets */
wire t_2743,   t_2744,   t_2745;
/* u2_941 Output nets */
wire t_2746,   t_2747,   t_2748;
/* u2_942 Output nets */
wire t_2749,   t_2750,   t_2751;
/* u2_943 Output nets */
wire t_2752,   t_2753,   t_2754;
/* u2_944 Output nets */
wire t_2755,   t_2756,   t_2757;
/* u2_945 Output nets */
wire t_2758,   t_2759,   t_2760;
/* u2_946 Output nets */
wire t_2761,   t_2762,   t_2763;
/* u2_947 Output nets */
wire t_2764,   t_2765,   t_2766;
/* u2_948 Output nets */
wire t_2767,   t_2768,   t_2769;
/* u2_949 Output nets */
wire t_2770,   t_2771,   t_2772;
/* u2_950 Output nets */
wire t_2773,   t_2774,   t_2775;
/* u2_951 Output nets */
wire t_2776,   t_2777,   t_2778;
/* u2_952 Output nets */
wire t_2779,   t_2780,   t_2781;
/* u2_953 Output nets */
wire t_2782,   t_2783,   t_2784;
/* u2_954 Output nets */
wire t_2785,   t_2786,   t_2787;
/* u2_955 Output nets */
wire t_2788,   t_2789,   t_2790;
/* u2_956 Output nets */
wire t_2791,   t_2792,   t_2793;
/* u2_957 Output nets */
wire t_2794,   t_2795,   t_2796;
/* u2_958 Output nets */
wire t_2797,   t_2798,   t_2799;
/* u2_959 Output nets */
wire t_2800,   t_2801,   t_2802;
/* u2_960 Output nets */
wire t_2803,   t_2804,   t_2805;
/* u2_961 Output nets */
wire t_2806,   t_2807,   t_2808;
/* u2_962 Output nets */
wire t_2809,   t_2810,   t_2811;
/* u2_963 Output nets */
wire t_2812,   t_2813,   t_2814;
/* u2_964 Output nets */
wire t_2815,   t_2816,   t_2817;
/* u2_965 Output nets */
wire t_2818,   t_2819,   t_2820;
/* u2_966 Output nets */
wire t_2821,   t_2822,   t_2823;
/* u2_967 Output nets */
wire t_2824,   t_2825,   t_2826;
/* u2_968 Output nets */
wire t_2827,   t_2828,   t_2829;
/* u2_969 Output nets */
wire t_2830,   t_2831,   t_2832;
/* u2_970 Output nets */
wire t_2833,   t_2834,   t_2835;
/* u2_971 Output nets */
wire t_2836,   t_2837,   t_2838;
/* u2_972 Output nets */
wire t_2839,   t_2840,   t_2841;
/* u2_973 Output nets */
wire t_2842,   t_2843,   t_2844;
/* u2_974 Output nets */
wire t_2845,   t_2846,   t_2847;
/* u0_975 Output nets */
wire t_2848,   t_2849;
/* u2_976 Output nets */
wire t_2850,   t_2851,   t_2852;
/* u2_977 Output nets */
wire t_2853,   t_2854,   t_2855;
/* u2_978 Output nets */
wire t_2856,   t_2857,   t_2858;
/* u2_979 Output nets */
wire t_2859,   t_2860,   t_2861;
/* u2_980 Output nets */
wire t_2862,   t_2863,   t_2864;
/* u2_981 Output nets */
wire t_2865,   t_2866,   t_2867;
/* u2_982 Output nets */
wire t_2868,   t_2869,   t_2870;
/* u2_983 Output nets */
wire t_2871,   t_2872,   t_2873;
/* u2_984 Output nets */
wire t_2874,   t_2875,   t_2876;
/* u2_985 Output nets */
wire t_2877,   t_2878,   t_2879;
/* u2_986 Output nets */
wire t_2880,   t_2881,   t_2882;
/* u2_987 Output nets */
wire t_2883,   t_2884,   t_2885;
/* u2_988 Output nets */
wire t_2886,   t_2887,   t_2888;
/* u2_989 Output nets */
wire t_2889,   t_2890,   t_2891;
/* u2_990 Output nets */
wire t_2892,   t_2893,   t_2894;
/* u0_991 Output nets */
wire t_2895,   t_2896;
/* u2_992 Output nets */
wire t_2897,   t_2898,   t_2899;
/* u2_993 Output nets */
wire t_2900,   t_2901,   t_2902;
/* u2_994 Output nets */
wire t_2903,   t_2904,   t_2905;
/* u2_995 Output nets */
wire t_2906,   t_2907,   t_2908;
/* u2_996 Output nets */
wire t_2909,   t_2910,   t_2911;
/* u2_997 Output nets */
wire t_2912,   t_2913,   t_2914;
/* u2_998 Output nets */
wire t_2915,   t_2916,   t_2917;
/* u2_999 Output nets */
wire t_2918,   t_2919,   t_2920;
/* u2_1000 Output nets */
wire t_2921,   t_2922,   t_2923;
/* u2_1001 Output nets */
wire t_2924,   t_2925,   t_2926;
/* u2_1002 Output nets */
wire t_2927,   t_2928,   t_2929;
/* u2_1003 Output nets */
wire t_2930,   t_2931,   t_2932;
/* u2_1004 Output nets */
wire t_2933,   t_2934,   t_2935;
/* u2_1005 Output nets */
wire t_2936,   t_2937,   t_2938;
/* u2_1006 Output nets */
wire t_2939,   t_2940,   t_2941;
/* u1_1007 Output nets */
wire t_2942,   t_2943;
/* u2_1008 Output nets */
wire t_2944,   t_2945,   t_2946;
/* u2_1009 Output nets */
wire t_2947,   t_2948,   t_2949;
/* u2_1010 Output nets */
wire t_2950,   t_2951,   t_2952;
/* u2_1011 Output nets */
wire t_2953,   t_2954,   t_2955;
/* u2_1012 Output nets */
wire t_2956,   t_2957,   t_2958;
/* u2_1013 Output nets */
wire t_2959,   t_2960,   t_2961;
/* u2_1014 Output nets */
wire t_2962,   t_2963,   t_2964;
/* u2_1015 Output nets */
wire t_2965,   t_2966,   t_2967;
/* u2_1016 Output nets */
wire t_2968,   t_2969,   t_2970;
/* u2_1017 Output nets */
wire t_2971,   t_2972,   t_2973;
/* u2_1018 Output nets */
wire t_2974,   t_2975,   t_2976;
/* u2_1019 Output nets */
wire t_2977,   t_2978,   t_2979;
/* u2_1020 Output nets */
wire t_2980,   t_2981,   t_2982;
/* u2_1021 Output nets */
wire t_2983,   t_2984,   t_2985;
/* u2_1022 Output nets */
wire t_2986,   t_2987,   t_2988;
/* u1_1023 Output nets */
wire t_2989,   t_2990;
/* u2_1024 Output nets */
wire t_2991,   t_2992,   t_2993;
/* u2_1025 Output nets */
wire t_2994,   t_2995,   t_2996;
/* u2_1026 Output nets */
wire t_2997,   t_2998,   t_2999;
/* u2_1027 Output nets */
wire t_3000,   t_3001,   t_3002;
/* u2_1028 Output nets */
wire t_3003,   t_3004,   t_3005;
/* u2_1029 Output nets */
wire t_3006,   t_3007,   t_3008;
/* u2_1030 Output nets */
wire t_3009,   t_3010,   t_3011;
/* u2_1031 Output nets */
wire t_3012,   t_3013,   t_3014;
/* u2_1032 Output nets */
wire t_3015,   t_3016,   t_3017;
/* u2_1033 Output nets */
wire t_3018,   t_3019,   t_3020;
/* u2_1034 Output nets */
wire t_3021,   t_3022,   t_3023;
/* u2_1035 Output nets */
wire t_3024,   t_3025,   t_3026;
/* u2_1036 Output nets */
wire t_3027,   t_3028,   t_3029;
/* u2_1037 Output nets */
wire t_3030,   t_3031,   t_3032;
/* u2_1038 Output nets */
wire t_3033,   t_3034,   t_3035;
/* u2_1039 Output nets */
wire t_3036,   t_3037,   t_3038;
/* u2_1040 Output nets */
wire t_3039,   t_3040,   t_3041;
/* u2_1041 Output nets */
wire t_3042,   t_3043,   t_3044;
/* u2_1042 Output nets */
wire t_3045,   t_3046,   t_3047;
/* u2_1043 Output nets */
wire t_3048,   t_3049,   t_3050;
/* u2_1044 Output nets */
wire t_3051,   t_3052,   t_3053;
/* u2_1045 Output nets */
wire t_3054,   t_3055,   t_3056;
/* u2_1046 Output nets */
wire t_3057,   t_3058,   t_3059;
/* u2_1047 Output nets */
wire t_3060,   t_3061,   t_3062;
/* u2_1048 Output nets */
wire t_3063,   t_3064,   t_3065;
/* u2_1049 Output nets */
wire t_3066,   t_3067,   t_3068;
/* u2_1050 Output nets */
wire t_3069,   t_3070,   t_3071;
/* u2_1051 Output nets */
wire t_3072,   t_3073,   t_3074;
/* u2_1052 Output nets */
wire t_3075,   t_3076,   t_3077;
/* u2_1053 Output nets */
wire t_3078,   t_3079,   t_3080;
/* u2_1054 Output nets */
wire t_3081,   t_3082,   t_3083;
/* u1_1055 Output nets */
wire t_3084,   t_3085;
/* u2_1056 Output nets */
wire t_3086,   t_3087,   t_3088;
/* u2_1057 Output nets */
wire t_3089,   t_3090,   t_3091;
/* u2_1058 Output nets */
wire t_3092,   t_3093,   t_3094;
/* u2_1059 Output nets */
wire t_3095,   t_3096,   t_3097;
/* u2_1060 Output nets */
wire t_3098,   t_3099,   t_3100;
/* u2_1061 Output nets */
wire t_3101,   t_3102,   t_3103;
/* u2_1062 Output nets */
wire t_3104,   t_3105,   t_3106;
/* u2_1063 Output nets */
wire t_3107,   t_3108,   t_3109;
/* u2_1064 Output nets */
wire t_3110,   t_3111,   t_3112;
/* u2_1065 Output nets */
wire t_3113,   t_3114,   t_3115;
/* u2_1066 Output nets */
wire t_3116,   t_3117,   t_3118;
/* u2_1067 Output nets */
wire t_3119,   t_3120,   t_3121;
/* u2_1068 Output nets */
wire t_3122,   t_3123,   t_3124;
/* u2_1069 Output nets */
wire t_3125,   t_3126,   t_3127;
/* u2_1070 Output nets */
wire t_3128,   t_3129,   t_3130;
/* u2_1071 Output nets */
wire t_3131,   t_3132,   t_3133;
/* u2_1072 Output nets */
wire t_3134,   t_3135,   t_3136;
/* u2_1073 Output nets */
wire t_3137,   t_3138,   t_3139;
/* u2_1074 Output nets */
wire t_3140,   t_3141,   t_3142;
/* u2_1075 Output nets */
wire t_3143,   t_3144,   t_3145;
/* u2_1076 Output nets */
wire t_3146,   t_3147,   t_3148;
/* u2_1077 Output nets */
wire t_3149,   t_3150,   t_3151;
/* u2_1078 Output nets */
wire t_3152,   t_3153,   t_3154;
/* u2_1079 Output nets */
wire t_3155,   t_3156,   t_3157;
/* u2_1080 Output nets */
wire t_3158,   t_3159,   t_3160;
/* u2_1081 Output nets */
wire t_3161,   t_3162,   t_3163;
/* u2_1082 Output nets */
wire t_3164,   t_3165,   t_3166;
/* u2_1083 Output nets */
wire t_3167,   t_3168,   t_3169;
/* u2_1084 Output nets */
wire t_3170,   t_3171,   t_3172;
/* u2_1085 Output nets */
wire t_3173,   t_3174,   t_3175;
/* u2_1086 Output nets */
wire t_3176,   t_3177,   t_3178;
/* u2_1087 Output nets */
wire t_3179,   t_3180,   t_3181;
/* u2_1088 Output nets */
wire t_3182,   t_3183,   t_3184;
/* u2_1089 Output nets */
wire t_3185,   t_3186,   t_3187;
/* u2_1090 Output nets */
wire t_3188,   t_3189,   t_3190;
/* u2_1091 Output nets */
wire t_3191,   t_3192,   t_3193;
/* u2_1092 Output nets */
wire t_3194,   t_3195,   t_3196;
/* u2_1093 Output nets */
wire t_3197,   t_3198,   t_3199;
/* u2_1094 Output nets */
wire t_3200,   t_3201,   t_3202;
/* u2_1095 Output nets */
wire t_3203,   t_3204,   t_3205;
/* u2_1096 Output nets */
wire t_3206,   t_3207,   t_3208;
/* u2_1097 Output nets */
wire t_3209,   t_3210,   t_3211;
/* u2_1098 Output nets */
wire t_3212,   t_3213,   t_3214;
/* u2_1099 Output nets */
wire t_3215,   t_3216,   t_3217;
/* u2_1100 Output nets */
wire t_3218,   t_3219,   t_3220;
/* u2_1101 Output nets */
wire t_3221,   t_3222,   t_3223;
/* u2_1102 Output nets */
wire t_3224,   t_3225,   t_3226;
/* u2_1103 Output nets */
wire t_3227,   t_3228,   t_3229;
/* u2_1104 Output nets */
wire t_3230,   t_3231,   t_3232;
/* u2_1105 Output nets */
wire t_3233,   t_3234,   t_3235;
/* u2_1106 Output nets */
wire t_3236,   t_3237,   t_3238;
/* u2_1107 Output nets */
wire t_3239,   t_3240,   t_3241;
/* u2_1108 Output nets */
wire t_3242,   t_3243,   t_3244;
/* u2_1109 Output nets */
wire t_3245,   t_3246,   t_3247;
/* u2_1110 Output nets */
wire t_3248,   t_3249,   t_3250;
/* u2_1111 Output nets */
wire t_3251,   t_3252,   t_3253;
/* u2_1112 Output nets */
wire t_3254,   t_3255,   t_3256;
/* u2_1113 Output nets */
wire t_3257,   t_3258,   t_3259;
/* u2_1114 Output nets */
wire t_3260,   t_3261,   t_3262;
/* u2_1115 Output nets */
wire t_3263,   t_3264,   t_3265;
/* u2_1116 Output nets */
wire t_3266,   t_3267,   t_3268;
/* u2_1117 Output nets */
wire t_3269,   t_3270,   t_3271;
/* u2_1118 Output nets */
wire t_3272,   t_3273,   t_3274;
/* u2_1119 Output nets */
wire t_3275,   t_3276,   t_3277;
/* u2_1120 Output nets */
wire t_3278,   t_3279,   t_3280;
/* u2_1121 Output nets */
wire t_3281,   t_3282,   t_3283;
/* u2_1122 Output nets */
wire t_3284,   t_3285,   t_3286;
/* u2_1123 Output nets */
wire t_3287,   t_3288,   t_3289;
/* u2_1124 Output nets */
wire t_3290,   t_3291,   t_3292;
/* u2_1125 Output nets */
wire t_3293,   t_3294,   t_3295;
/* u2_1126 Output nets */
wire t_3296,   t_3297,   t_3298;
/* u2_1127 Output nets */
wire t_3299,   t_3300,   t_3301;
/* u2_1128 Output nets */
wire t_3302,   t_3303,   t_3304;
/* u2_1129 Output nets */
wire t_3305,   t_3306,   t_3307;
/* u2_1130 Output nets */
wire t_3308,   t_3309,   t_3310;
/* u2_1131 Output nets */
wire t_3311,   t_3312,   t_3313;
/* u2_1132 Output nets */
wire t_3314,   t_3315,   t_3316;
/* u2_1133 Output nets */
wire t_3317,   t_3318,   t_3319;
/* u2_1134 Output nets */
wire t_3320,   t_3321,   t_3322;
/* u2_1135 Output nets */
wire t_3323,   t_3324,   t_3325;
/* u2_1136 Output nets */
wire t_3326,   t_3327,   t_3328;
/* u2_1137 Output nets */
wire t_3329,   t_3330,   t_3331;
/* u2_1138 Output nets */
wire t_3332,   t_3333,   t_3334;
/* u2_1139 Output nets */
wire t_3335,   t_3336,   t_3337;
/* u2_1140 Output nets */
wire t_3338,   t_3339,   t_3340;
/* u2_1141 Output nets */
wire t_3341,   t_3342,   t_3343;
/* u2_1142 Output nets */
wire t_3344,   t_3345,   t_3346;
/* u2_1143 Output nets */
wire t_3347,   t_3348,   t_3349;
/* u2_1144 Output nets */
wire t_3350,   t_3351,   t_3352;
/* u2_1145 Output nets */
wire t_3353,   t_3354,   t_3355;
/* u2_1146 Output nets */
wire t_3356,   t_3357,   t_3358;
/* u2_1147 Output nets */
wire t_3359,   t_3360,   t_3361;
/* u2_1148 Output nets */
wire t_3362,   t_3363,   t_3364;
/* u2_1149 Output nets */
wire t_3365,   t_3366,   t_3367;
/* u2_1150 Output nets */
wire t_3368,   t_3369,   t_3370;
/* u2_1151 Output nets */
wire t_3371,   t_3372,   t_3373;
/* u2_1152 Output nets */
wire t_3374,   t_3375,   t_3376;
/* u2_1153 Output nets */
wire t_3377,   t_3378,   t_3379;
/* u2_1154 Output nets */
wire t_3380,   t_3381,   t_3382;
/* u2_1155 Output nets */
wire t_3383,   t_3384,   t_3385;
/* u2_1156 Output nets */
wire t_3386,   t_3387,   t_3388;
/* u2_1157 Output nets */
wire t_3389,   t_3390,   t_3391;
/* u2_1158 Output nets */
wire t_3392,   t_3393,   t_3394;
/* u2_1159 Output nets */
wire t_3395,   t_3396,   t_3397;
/* u2_1160 Output nets */
wire t_3398,   t_3399,   t_3400;
/* u2_1161 Output nets */
wire t_3401,   t_3402,   t_3403;
/* u2_1162 Output nets */
wire t_3404,   t_3405,   t_3406;
/* u2_1163 Output nets */
wire t_3407,   t_3408,   t_3409;
/* u2_1164 Output nets */
wire t_3410,   t_3411,   t_3412;
/* u2_1165 Output nets */
wire t_3413,   t_3414,   t_3415;
/* u2_1166 Output nets */
wire t_3416,   t_3417,   t_3418;
/* u1_1167 Output nets */
wire t_3419,   t_3420;
/* u2_1168 Output nets */
wire t_3421,   t_3422,   t_3423;
/* u2_1169 Output nets */
wire t_3424,   t_3425,   t_3426;
/* u2_1170 Output nets */
wire t_3427,   t_3428,   t_3429;
/* u2_1171 Output nets */
wire t_3430,   t_3431,   t_3432;
/* u2_1172 Output nets */
wire t_3433,   t_3434,   t_3435;
/* u2_1173 Output nets */
wire t_3436,   t_3437,   t_3438;
/* u2_1174 Output nets */
wire t_3439,   t_3440,   t_3441;
/* u2_1175 Output nets */
wire t_3442,   t_3443,   t_3444;
/* u2_1176 Output nets */
wire t_3445,   t_3446,   t_3447;
/* u2_1177 Output nets */
wire t_3448,   t_3449,   t_3450;
/* u2_1178 Output nets */
wire t_3451,   t_3452,   t_3453;
/* u2_1179 Output nets */
wire t_3454,   t_3455,   t_3456;
/* u2_1180 Output nets */
wire t_3457,   t_3458,   t_3459;
/* u2_1181 Output nets */
wire t_3460,   t_3461,   t_3462;
/* u2_1182 Output nets */
wire t_3463,   t_3464,   t_3465;
/* u1_1183 Output nets */
wire t_3466,   t_3467;
/* u2_1184 Output nets */
wire t_3468,   t_3469,   t_3470;
/* u2_1185 Output nets */
wire t_3471,   t_3472,   t_3473;
/* u2_1186 Output nets */
wire t_3474,   t_3475,   t_3476;
/* u2_1187 Output nets */
wire t_3477,   t_3478,   t_3479;
/* u2_1188 Output nets */
wire t_3480,   t_3481,   t_3482;
/* u2_1189 Output nets */
wire t_3483,   t_3484,   t_3485;
/* u2_1190 Output nets */
wire t_3486,   t_3487,   t_3488;
/* u2_1191 Output nets */
wire t_3489,   t_3490,   t_3491;
/* u2_1192 Output nets */
wire t_3492,   t_3493,   t_3494;
/* u2_1193 Output nets */
wire t_3495,   t_3496,   t_3497;
/* u2_1194 Output nets */
wire t_3498,   t_3499,   t_3500;
/* u2_1195 Output nets */
wire t_3501,   t_3502,   t_3503;
/* u2_1196 Output nets */
wire t_3504,   t_3505,   t_3506;
/* u2_1197 Output nets */
wire t_3507,   t_3508,   t_3509;
/* u2_1198 Output nets */
wire t_3510,   t_3511,   t_3512;
/* u1_1199 Output nets */
wire t_3513,   t_3514;
/* u2_1200 Output nets */
wire t_3515,   t_3516,   t_3517;
/* u2_1201 Output nets */
wire t_3518,   t_3519,   t_3520;
/* u2_1202 Output nets */
wire t_3521,   t_3522,   t_3523;
/* u2_1203 Output nets */
wire t_3524,   t_3525,   t_3526;
/* u2_1204 Output nets */
wire t_3527,   t_3528,   t_3529;
/* u2_1205 Output nets */
wire t_3530,   t_3531,   t_3532;
/* u2_1206 Output nets */
wire t_3533,   t_3534,   t_3535;
/* u2_1207 Output nets */
wire t_3536,   t_3537,   t_3538;
/* u2_1208 Output nets */
wire t_3539,   t_3540,   t_3541;
/* u2_1209 Output nets */
wire t_3542,   t_3543,   t_3544;
/* u2_1210 Output nets */
wire t_3545,   t_3546,   t_3547;
/* u2_1211 Output nets */
wire t_3548,   t_3549,   t_3550;
/* u2_1212 Output nets */
wire t_3551,   t_3552,   t_3553;
/* u2_1213 Output nets */
wire t_3554,   t_3555,   t_3556;
/* u2_1214 Output nets */
wire t_3557,   t_3558,   t_3559;
/* u1_1215 Output nets */
wire t_3560,   t_3561;
/* u2_1216 Output nets */
wire t_3562,   t_3563,   t_3564;
/* u2_1217 Output nets */
wire t_3565,   t_3566,   t_3567;
/* u2_1218 Output nets */
wire t_3568,   t_3569,   t_3570;
/* u2_1219 Output nets */
wire t_3571,   t_3572,   t_3573;
/* u2_1220 Output nets */
wire t_3574,   t_3575,   t_3576;
/* u2_1221 Output nets */
wire t_3577,   t_3578,   t_3579;
/* u2_1222 Output nets */
wire t_3580,   t_3581,   t_3582;
/* u2_1223 Output nets */
wire t_3583,   t_3584,   t_3585;
/* u2_1224 Output nets */
wire t_3586,   t_3587,   t_3588;
/* u2_1225 Output nets */
wire t_3589,   t_3590,   t_3591;
/* u2_1226 Output nets */
wire t_3592,   t_3593,   t_3594;
/* u2_1227 Output nets */
wire t_3595,   t_3596,   t_3597;
/* u2_1228 Output nets */
wire t_3598,   t_3599,   t_3600;
/* u2_1229 Output nets */
wire t_3601,   t_3602,   t_3603;
/* u2_1230 Output nets */
wire t_3604,   t_3605,   t_3606;
/* u0_1231 Output nets */
wire t_3607,   t_3608;
/* u2_1232 Output nets */
wire t_3609,   t_3610,   t_3611;
/* u2_1233 Output nets */
wire t_3612,   t_3613,   t_3614;
/* u2_1234 Output nets */
wire t_3615,   t_3616,   t_3617;
/* u2_1235 Output nets */
wire t_3618,   t_3619,   t_3620;
/* u2_1236 Output nets */
wire t_3621,   t_3622,   t_3623;
/* u2_1237 Output nets */
wire t_3624,   t_3625,   t_3626;
/* u2_1238 Output nets */
wire t_3627,   t_3628,   t_3629;
/* u2_1239 Output nets */
wire t_3630,   t_3631,   t_3632;
/* u2_1240 Output nets */
wire t_3633,   t_3634,   t_3635;
/* u2_1241 Output nets */
wire t_3636,   t_3637,   t_3638;
/* u2_1242 Output nets */
wire t_3639,   t_3640,   t_3641;
/* u2_1243 Output nets */
wire t_3642,   t_3643,   t_3644;
/* u2_1244 Output nets */
wire t_3645,   t_3646,   t_3647;
/* u2_1245 Output nets */
wire t_3648,   t_3649,   t_3650;
/* u2_1246 Output nets */
wire t_3651,   t_3652,   t_3653;
/* u0_1247 Output nets */
wire t_3654,   t_3655;
/* u2_1248 Output nets */
wire t_3656,   t_3657,   t_3658;
/* u2_1249 Output nets */
wire t_3659,   t_3660,   t_3661;
/* u2_1250 Output nets */
wire t_3662,   t_3663,   t_3664;
/* u2_1251 Output nets */
wire t_3665,   t_3666,   t_3667;
/* u2_1252 Output nets */
wire t_3668,   t_3669,   t_3670;
/* u2_1253 Output nets */
wire t_3671,   t_3672,   t_3673;
/* u2_1254 Output nets */
wire t_3674,   t_3675,   t_3676;
/* u2_1255 Output nets */
wire t_3677,   t_3678,   t_3679;
/* u2_1256 Output nets */
wire t_3680,   t_3681,   t_3682;
/* u2_1257 Output nets */
wire t_3683,   t_3684,   t_3685;
/* u2_1258 Output nets */
wire t_3686,   t_3687,   t_3688;
/* u2_1259 Output nets */
wire t_3689,   t_3690,   t_3691;
/* u2_1260 Output nets */
wire t_3692,   t_3693,   t_3694;
/* u2_1261 Output nets */
wire t_3695,   t_3696,   t_3697;
/* u2_1262 Output nets */
wire t_3698,   t_3699,   t_3700;
/* u2_1263 Output nets */
wire t_3701,   t_3702,   t_3703;
/* u2_1264 Output nets */
wire t_3704,   t_3705,   t_3706;
/* u2_1265 Output nets */
wire t_3707,   t_3708,   t_3709;
/* u2_1266 Output nets */
wire t_3710,   t_3711,   t_3712;
/* u2_1267 Output nets */
wire t_3713,   t_3714,   t_3715;
/* u2_1268 Output nets */
wire t_3716,   t_3717,   t_3718;
/* u2_1269 Output nets */
wire t_3719,   t_3720,   t_3721;
/* u2_1270 Output nets */
wire t_3722,   t_3723,   t_3724;
/* u2_1271 Output nets */
wire t_3725,   t_3726,   t_3727;
/* u2_1272 Output nets */
wire t_3728,   t_3729,   t_3730;
/* u2_1273 Output nets */
wire t_3731,   t_3732,   t_3733;
/* u2_1274 Output nets */
wire t_3734,   t_3735,   t_3736;
/* u2_1275 Output nets */
wire t_3737,   t_3738,   t_3739;
/* u2_1276 Output nets */
wire t_3740,   t_3741,   t_3742;
/* u2_1277 Output nets */
wire t_3743,   t_3744,   t_3745;
/* u2_1278 Output nets */
wire t_3746,   t_3747,   t_3748;
/* u2_1279 Output nets */
wire t_3749,   t_3750,   t_3751;
/* u2_1280 Output nets */
wire t_3752,   t_3753,   t_3754;
/* u2_1281 Output nets */
wire t_3755,   t_3756,   t_3757;
/* u2_1282 Output nets */
wire t_3758,   t_3759,   t_3760;
/* u2_1283 Output nets */
wire t_3761,   t_3762,   t_3763;
/* u2_1284 Output nets */
wire t_3764,   t_3765,   t_3766;
/* u2_1285 Output nets */
wire t_3767,   t_3768,   t_3769;
/* u2_1286 Output nets */
wire t_3770,   t_3771,   t_3772;
/* u2_1287 Output nets */
wire t_3773,   t_3774,   t_3775;
/* u2_1288 Output nets */
wire t_3776,   t_3777,   t_3778;
/* u2_1289 Output nets */
wire t_3779,   t_3780,   t_3781;
/* u2_1290 Output nets */
wire t_3782,   t_3783,   t_3784;
/* u2_1291 Output nets */
wire t_3785,   t_3786,   t_3787;
/* u1_1292 Output nets */
wire t_3788,   t_3789;
/* u2_1293 Output nets */
wire t_3790,   t_3791,   t_3792;
/* u2_1294 Output nets */
wire t_3793,   t_3794,   t_3795;
/* u2_1295 Output nets */
wire t_3796,   t_3797,   t_3798;
/* u2_1296 Output nets */
wire t_3799,   t_3800,   t_3801;
/* u2_1297 Output nets */
wire t_3802,   t_3803,   t_3804;
/* u2_1298 Output nets */
wire t_3805,   t_3806,   t_3807;
/* u2_1299 Output nets */
wire t_3808,   t_3809,   t_3810;
/* u2_1300 Output nets */
wire t_3811,   t_3812,   t_3813;
/* u2_1301 Output nets */
wire t_3814,   t_3815,   t_3816;
/* u2_1302 Output nets */
wire t_3817,   t_3818,   t_3819;
/* u2_1303 Output nets */
wire t_3820,   t_3821,   t_3822;
/* u2_1304 Output nets */
wire t_3823,   t_3824,   t_3825;
/* u2_1305 Output nets */
wire t_3826,   t_3827,   t_3828;
/* u2_1306 Output nets */
wire t_3829,   t_3830,   t_3831;
/* u1_1307 Output nets */
wire t_3832,   t_3833;
/* u2_1308 Output nets */
wire t_3834,   t_3835,   t_3836;
/* u2_1309 Output nets */
wire t_3837,   t_3838,   t_3839;
/* u2_1310 Output nets */
wire t_3840,   t_3841,   t_3842;
/* u2_1311 Output nets */
wire t_3843,   t_3844,   t_3845;
/* u2_1312 Output nets */
wire t_3846,   t_3847,   t_3848;
/* u2_1313 Output nets */
wire t_3849,   t_3850,   t_3851;
/* u2_1314 Output nets */
wire t_3852,   t_3853,   t_3854;
/* u2_1315 Output nets */
wire t_3855,   t_3856,   t_3857;
/* u2_1316 Output nets */
wire t_3858,   t_3859,   t_3860;
/* u2_1317 Output nets */
wire t_3861,   t_3862,   t_3863;
/* u2_1318 Output nets */
wire t_3864,   t_3865,   t_3866;
/* u2_1319 Output nets */
wire t_3867,   t_3868,   t_3869;
/* u2_1320 Output nets */
wire t_3870,   t_3871,   t_3872;
/* u2_1321 Output nets */
wire t_3873,   t_3874,   t_3875;
/* u1_1322 Output nets */
wire t_3876,   t_3877;
/* u2_1323 Output nets */
wire t_3878,   t_3879,   t_3880;
/* u2_1324 Output nets */
wire t_3881,   t_3882,   t_3883;
/* u2_1325 Output nets */
wire t_3884,   t_3885,   t_3886;
/* u2_1326 Output nets */
wire t_3887,   t_3888,   t_3889;
/* u2_1327 Output nets */
wire t_3890,   t_3891,   t_3892;
/* u2_1328 Output nets */
wire t_3893,   t_3894,   t_3895;
/* u2_1329 Output nets */
wire t_3896,   t_3897,   t_3898;
/* u2_1330 Output nets */
wire t_3899,   t_3900,   t_3901;
/* u2_1331 Output nets */
wire t_3902,   t_3903,   t_3904;
/* u2_1332 Output nets */
wire t_3905,   t_3906,   t_3907;
/* u2_1333 Output nets */
wire t_3908,   t_3909,   t_3910;
/* u2_1334 Output nets */
wire t_3911,   t_3912,   t_3913;
/* u2_1335 Output nets */
wire t_3914,   t_3915,   t_3916;
/* u2_1336 Output nets */
wire t_3917,   t_3918,   t_3919;
/* u1_1337 Output nets */
wire t_3920,   t_3921;
/* u2_1338 Output nets */
wire t_3922,   t_3923,   t_3924;
/* u2_1339 Output nets */
wire t_3925,   t_3926,   t_3927;
/* u2_1340 Output nets */
wire t_3928,   t_3929,   t_3930;
/* u2_1341 Output nets */
wire t_3931,   t_3932,   t_3933;
/* u2_1342 Output nets */
wire t_3934,   t_3935,   t_3936;
/* u2_1343 Output nets */
wire t_3937,   t_3938,   t_3939;
/* u2_1344 Output nets */
wire t_3940,   t_3941,   t_3942;
/* u2_1345 Output nets */
wire t_3943,   t_3944,   t_3945;
/* u2_1346 Output nets */
wire t_3946,   t_3947,   t_3948;
/* u2_1347 Output nets */
wire t_3949,   t_3950,   t_3951;
/* u2_1348 Output nets */
wire t_3952,   t_3953,   t_3954;
/* u2_1349 Output nets */
wire t_3955,   t_3956,   t_3957;
/* u2_1350 Output nets */
wire t_3958,   t_3959,   t_3960;
/* u2_1351 Output nets */
wire t_3961,   t_3962,   t_3963;
/* u0_1352 Output nets */
wire t_3964,   t_3965;
/* u2_1353 Output nets */
wire t_3966,   t_3967,   t_3968;
/* u2_1354 Output nets */
wire t_3969,   t_3970,   t_3971;
/* u2_1355 Output nets */
wire t_3972,   t_3973,   t_3974;
/* u2_1356 Output nets */
wire t_3975,   t_3976,   t_3977;
/* u2_1357 Output nets */
wire t_3978,   t_3979,   t_3980;
/* u2_1358 Output nets */
wire t_3981,   t_3982,   t_3983;
/* u2_1359 Output nets */
wire t_3984,   t_3985,   t_3986;
/* u2_1360 Output nets */
wire t_3987,   t_3988,   t_3989;
/* u2_1361 Output nets */
wire t_3990,   t_3991,   t_3992;
/* u2_1362 Output nets */
wire t_3993,   t_3994,   t_3995;
/* u2_1363 Output nets */
wire t_3996,   t_3997,   t_3998;
/* u2_1364 Output nets */
wire t_3999,   t_4000,   t_4001;
/* u2_1365 Output nets */
wire t_4002,   t_4003,   t_4004;
/* u2_1366 Output nets */
wire t_4005,   t_4006,   t_4007;
/* u0_1367 Output nets */
wire t_4008,   t_4009;
/* u2_1368 Output nets */
wire t_4010,   t_4011,   t_4012;
/* u2_1369 Output nets */
wire t_4013,   t_4014,   t_4015;
/* u2_1370 Output nets */
wire t_4016,   t_4017,   t_4018;
/* u2_1371 Output nets */
wire t_4019,   t_4020,   t_4021;
/* u2_1372 Output nets */
wire t_4022,   t_4023,   t_4024;
/* u2_1373 Output nets */
wire t_4025,   t_4026,   t_4027;
/* u2_1374 Output nets */
wire t_4028,   t_4029,   t_4030;
/* u2_1375 Output nets */
wire t_4031,   t_4032,   t_4033;
/* u2_1376 Output nets */
wire t_4034,   t_4035,   t_4036;
/* u2_1377 Output nets */
wire t_4037,   t_4038,   t_4039;
/* u2_1378 Output nets */
wire t_4040,   t_4041,   t_4042;
/* u2_1379 Output nets */
wire t_4043,   t_4044,   t_4045;
/* u2_1380 Output nets */
wire t_4046,   t_4047,   t_4048;
/* u2_1381 Output nets */
wire t_4049,   t_4050,   t_4051;
/* u2_1382 Output nets */
wire t_4052,   t_4053,   t_4054;
/* u2_1383 Output nets */
wire t_4055,   t_4056,   t_4057;
/* u2_1384 Output nets */
wire t_4058,   t_4059,   t_4060;
/* u2_1385 Output nets */
wire t_4061,   t_4062,   t_4063;
/* u2_1386 Output nets */
wire t_4064,   t_4065,   t_4066;
/* u2_1387 Output nets */
wire t_4067,   t_4068,   t_4069;
/* u2_1388 Output nets */
wire t_4070,   t_4071,   t_4072;
/* u2_1389 Output nets */
wire t_4073,   t_4074,   t_4075;
/* u2_1390 Output nets */
wire t_4076,   t_4077,   t_4078;
/* u2_1391 Output nets */
wire t_4079,   t_4080,   t_4081;
/* u2_1392 Output nets */
wire t_4082,   t_4083,   t_4084;
/* u2_1393 Output nets */
wire t_4085,   t_4086,   t_4087;
/* u2_1394 Output nets */
wire t_4088,   t_4089,   t_4090;
/* u2_1395 Output nets */
wire t_4091,   t_4092,   t_4093;
/* u2_1396 Output nets */
wire t_4094,   t_4095,   t_4096;
/* u2_1397 Output nets */
wire t_4097,   t_4098,   t_4099;
/* u2_1398 Output nets */
wire t_4100,   t_4101,   t_4102;
/* u2_1399 Output nets */
wire t_4103,   t_4104,   t_4105;
/* u2_1400 Output nets */
wire t_4106,   t_4107,   t_4108;
/* u2_1401 Output nets */
wire t_4109,   t_4110,   t_4111;
/* u2_1402 Output nets */
wire t_4112,   t_4113,   t_4114;
/* u2_1403 Output nets */
wire t_4115,   t_4116,   t_4117;
/* u2_1404 Output nets */
wire t_4118,   t_4119,   t_4120;
/* u2_1405 Output nets */
wire t_4121,   t_4122,   t_4123;
/* u2_1406 Output nets */
wire t_4124,   t_4125,   t_4126;
/* u2_1407 Output nets */
wire t_4127,   t_4128,   t_4129;
/* u2_1408 Output nets */
wire t_4130,   t_4131,   t_4132;
/* u1_1409 Output nets */
wire t_4133,   t_4134;
/* u2_1410 Output nets */
wire t_4135,   t_4136,   t_4137;
/* u2_1411 Output nets */
wire t_4138,   t_4139,   t_4140;
/* u2_1412 Output nets */
wire t_4141,   t_4142,   t_4143;
/* u2_1413 Output nets */
wire t_4144,   t_4145,   t_4146;
/* u2_1414 Output nets */
wire t_4147,   t_4148,   t_4149;
/* u2_1415 Output nets */
wire t_4150,   t_4151,   t_4152;
/* u2_1416 Output nets */
wire t_4153,   t_4154,   t_4155;
/* u2_1417 Output nets */
wire t_4156,   t_4157,   t_4158;
/* u2_1418 Output nets */
wire t_4159,   t_4160,   t_4161;
/* u2_1419 Output nets */
wire t_4162,   t_4163,   t_4164;
/* u2_1420 Output nets */
wire t_4165,   t_4166,   t_4167;
/* u2_1421 Output nets */
wire t_4168,   t_4169,   t_4170;
/* u2_1422 Output nets */
wire t_4171,   t_4172,   t_4173;
/* u1_1423 Output nets */
wire t_4174,   t_4175;
/* u2_1424 Output nets */
wire t_4176,   t_4177,   t_4178;
/* u2_1425 Output nets */
wire t_4179,   t_4180,   t_4181;
/* u2_1426 Output nets */
wire t_4182,   t_4183,   t_4184;
/* u2_1427 Output nets */
wire t_4185,   t_4186,   t_4187;
/* u2_1428 Output nets */
wire t_4188,   t_4189,   t_4190;
/* u2_1429 Output nets */
wire t_4191,   t_4192,   t_4193;
/* u2_1430 Output nets */
wire t_4194,   t_4195,   t_4196;
/* u2_1431 Output nets */
wire t_4197,   t_4198,   t_4199;
/* u2_1432 Output nets */
wire t_4200,   t_4201,   t_4202;
/* u2_1433 Output nets */
wire t_4203,   t_4204,   t_4205;
/* u2_1434 Output nets */
wire t_4206,   t_4207,   t_4208;
/* u2_1435 Output nets */
wire t_4209,   t_4210,   t_4211;
/* u2_1436 Output nets */
wire t_4212,   t_4213,   t_4214;
/* u1_1437 Output nets */
wire t_4215,   t_4216;
/* u2_1438 Output nets */
wire t_4217,   t_4218,   t_4219;
/* u2_1439 Output nets */
wire t_4220,   t_4221,   t_4222;
/* u2_1440 Output nets */
wire t_4223,   t_4224,   t_4225;
/* u2_1441 Output nets */
wire t_4226,   t_4227,   t_4228;
/* u2_1442 Output nets */
wire t_4229,   t_4230,   t_4231;
/* u2_1443 Output nets */
wire t_4232,   t_4233,   t_4234;
/* u2_1444 Output nets */
wire t_4235,   t_4236,   t_4237;
/* u2_1445 Output nets */
wire t_4238,   t_4239,   t_4240;
/* u2_1446 Output nets */
wire t_4241,   t_4242,   t_4243;
/* u2_1447 Output nets */
wire t_4244,   t_4245,   t_4246;
/* u2_1448 Output nets */
wire t_4247,   t_4248,   t_4249;
/* u2_1449 Output nets */
wire t_4250,   t_4251,   t_4252;
/* u2_1450 Output nets */
wire t_4253,   t_4254,   t_4255;
/* u1_1451 Output nets */
wire t_4256,   t_4257;
/* u2_1452 Output nets */
wire t_4258,   t_4259,   t_4260;
/* u2_1453 Output nets */
wire t_4261,   t_4262,   t_4263;
/* u2_1454 Output nets */
wire t_4264,   t_4265,   t_4266;
/* u2_1455 Output nets */
wire t_4267,   t_4268,   t_4269;
/* u2_1456 Output nets */
wire t_4270,   t_4271,   t_4272;
/* u2_1457 Output nets */
wire t_4273,   t_4274,   t_4275;
/* u2_1458 Output nets */
wire t_4276,   t_4277,   t_4278;
/* u2_1459 Output nets */
wire t_4279,   t_4280,   t_4281;
/* u2_1460 Output nets */
wire t_4282,   t_4283,   t_4284;
/* u2_1461 Output nets */
wire t_4285,   t_4286,   t_4287;
/* u2_1462 Output nets */
wire t_4288,   t_4289,   t_4290;
/* u2_1463 Output nets */
wire t_4291,   t_4292,   t_4293;
/* u2_1464 Output nets */
wire t_4294,   t_4295,   t_4296;
/* u0_1465 Output nets */
wire t_4297,   t_4298;
/* u2_1466 Output nets */
wire t_4299,   t_4300,   t_4301;
/* u2_1467 Output nets */
wire t_4302,   t_4303,   t_4304;
/* u2_1468 Output nets */
wire t_4305,   t_4306,   t_4307;
/* u2_1469 Output nets */
wire t_4308,   t_4309,   t_4310;
/* u2_1470 Output nets */
wire t_4311,   t_4312,   t_4313;
/* u2_1471 Output nets */
wire t_4314,   t_4315,   t_4316;
/* u2_1472 Output nets */
wire t_4317,   t_4318,   t_4319;
/* u2_1473 Output nets */
wire t_4320,   t_4321,   t_4322;
/* u2_1474 Output nets */
wire t_4323,   t_4324,   t_4325;
/* u2_1475 Output nets */
wire t_4326,   t_4327,   t_4328;
/* u2_1476 Output nets */
wire t_4329,   t_4330,   t_4331;
/* u2_1477 Output nets */
wire t_4332,   t_4333,   t_4334;
/* u2_1478 Output nets */
wire t_4335,   t_4336,   t_4337;
/* u0_1479 Output nets */
wire t_4338,   t_4339;
/* u2_1480 Output nets */
wire t_4340,   t_4341,   t_4342;
/* u2_1481 Output nets */
wire t_4343,   t_4344,   t_4345;
/* u2_1482 Output nets */
wire t_4346,   t_4347,   t_4348;
/* u2_1483 Output nets */
wire t_4349,   t_4350,   t_4351;
/* u2_1484 Output nets */
wire t_4352,   t_4353,   t_4354;
/* u2_1485 Output nets */
wire t_4355,   t_4356,   t_4357;
/* u2_1486 Output nets */
wire t_4358,   t_4359,   t_4360;
/* u2_1487 Output nets */
wire t_4361,   t_4362,   t_4363;
/* u2_1488 Output nets */
wire t_4364,   t_4365,   t_4366;
/* u2_1489 Output nets */
wire t_4367,   t_4368,   t_4369;
/* u2_1490 Output nets */
wire t_4370,   t_4371,   t_4372;
/* u2_1491 Output nets */
wire t_4373,   t_4374,   t_4375;
/* u2_1492 Output nets */
wire t_4376,   t_4377,   t_4378;
/* u2_1493 Output nets */
wire t_4379,   t_4380,   t_4381;
/* u2_1494 Output nets */
wire t_4382,   t_4383,   t_4384;
/* u2_1495 Output nets */
wire t_4385,   t_4386,   t_4387;
/* u2_1496 Output nets */
wire t_4388,   t_4389,   t_4390;
/* u2_1497 Output nets */
wire t_4391,   t_4392,   t_4393;
/* u2_1498 Output nets */
wire t_4394,   t_4395,   t_4396;
/* u2_1499 Output nets */
wire t_4397,   t_4398,   t_4399;
/* u2_1500 Output nets */
wire t_4400,   t_4401,   t_4402;
/* u2_1501 Output nets */
wire t_4403,   t_4404,   t_4405;
/* u2_1502 Output nets */
wire t_4406,   t_4407,   t_4408;
/* u2_1503 Output nets */
wire t_4409,   t_4410,   t_4411;
/* u2_1504 Output nets */
wire t_4412,   t_4413,   t_4414;
/* u2_1505 Output nets */
wire t_4415,   t_4416,   t_4417;
/* u2_1506 Output nets */
wire t_4418,   t_4419,   t_4420;
/* u2_1507 Output nets */
wire t_4421,   t_4422,   t_4423;
/* u2_1508 Output nets */
wire t_4424,   t_4425,   t_4426;
/* u2_1509 Output nets */
wire t_4427,   t_4428,   t_4429;
/* u2_1510 Output nets */
wire t_4430,   t_4431,   t_4432;
/* u2_1511 Output nets */
wire t_4433,   t_4434,   t_4435;
/* u2_1512 Output nets */
wire t_4436,   t_4437,   t_4438;
/* u2_1513 Output nets */
wire t_4439,   t_4440,   t_4441;
/* u2_1514 Output nets */
wire t_4442,   t_4443,   t_4444;
/* u2_1515 Output nets */
wire t_4445,   t_4446,   t_4447;
/* u2_1516 Output nets */
wire t_4448,   t_4449,   t_4450;
/* u2_1517 Output nets */
wire t_4451,   t_4452,   t_4453;
/* u1_1518 Output nets */
wire t_4454,   t_4455;
/* u2_1519 Output nets */
wire t_4456,   t_4457,   t_4458;
/* u2_1520 Output nets */
wire t_4459,   t_4460,   t_4461;
/* u2_1521 Output nets */
wire t_4462,   t_4463,   t_4464;
/* u2_1522 Output nets */
wire t_4465,   t_4466,   t_4467;
/* u2_1523 Output nets */
wire t_4468,   t_4469,   t_4470;
/* u2_1524 Output nets */
wire t_4471,   t_4472,   t_4473;
/* u2_1525 Output nets */
wire t_4474,   t_4475,   t_4476;
/* u2_1526 Output nets */
wire t_4477,   t_4478,   t_4479;
/* u2_1527 Output nets */
wire t_4480,   t_4481,   t_4482;
/* u2_1528 Output nets */
wire t_4483,   t_4484,   t_4485;
/* u2_1529 Output nets */
wire t_4486,   t_4487,   t_4488;
/* u2_1530 Output nets */
wire t_4489,   t_4490,   t_4491;
/* u1_1531 Output nets */
wire t_4492,   t_4493;
/* u2_1532 Output nets */
wire t_4494,   t_4495,   t_4496;
/* u2_1533 Output nets */
wire t_4497,   t_4498,   t_4499;
/* u2_1534 Output nets */
wire t_4500,   t_4501,   t_4502;
/* u2_1535 Output nets */
wire t_4503,   t_4504,   t_4505;
/* u2_1536 Output nets */
wire t_4506,   t_4507,   t_4508;
/* u2_1537 Output nets */
wire t_4509,   t_4510,   t_4511;
/* u2_1538 Output nets */
wire t_4512,   t_4513,   t_4514;
/* u2_1539 Output nets */
wire t_4515,   t_4516,   t_4517;
/* u2_1540 Output nets */
wire t_4518,   t_4519,   t_4520;
/* u2_1541 Output nets */
wire t_4521,   t_4522,   t_4523;
/* u2_1542 Output nets */
wire t_4524,   t_4525,   t_4526;
/* u2_1543 Output nets */
wire t_4527,   t_4528,   t_4529;
/* u1_1544 Output nets */
wire t_4530,   t_4531;
/* u2_1545 Output nets */
wire t_4532,   t_4533,   t_4534;
/* u2_1546 Output nets */
wire t_4535,   t_4536,   t_4537;
/* u2_1547 Output nets */
wire t_4538,   t_4539,   t_4540;
/* u2_1548 Output nets */
wire t_4541,   t_4542,   t_4543;
/* u2_1549 Output nets */
wire t_4544,   t_4545,   t_4546;
/* u2_1550 Output nets */
wire t_4547,   t_4548,   t_4549;
/* u2_1551 Output nets */
wire t_4550,   t_4551,   t_4552;
/* u2_1552 Output nets */
wire t_4553,   t_4554,   t_4555;
/* u2_1553 Output nets */
wire t_4556,   t_4557,   t_4558;
/* u2_1554 Output nets */
wire t_4559,   t_4560,   t_4561;
/* u2_1555 Output nets */
wire t_4562,   t_4563,   t_4564;
/* u2_1556 Output nets */
wire t_4565,   t_4566,   t_4567;
/* u1_1557 Output nets */
wire t_4568,   t_4569;
/* u2_1558 Output nets */
wire t_4570,   t_4571,   t_4572;
/* u2_1559 Output nets */
wire t_4573,   t_4574,   t_4575;
/* u2_1560 Output nets */
wire t_4576,   t_4577,   t_4578;
/* u2_1561 Output nets */
wire t_4579,   t_4580,   t_4581;
/* u2_1562 Output nets */
wire t_4582,   t_4583,   t_4584;
/* u2_1563 Output nets */
wire t_4585,   t_4586,   t_4587;
/* u2_1564 Output nets */
wire t_4588,   t_4589,   t_4590;
/* u2_1565 Output nets */
wire t_4591,   t_4592,   t_4593;
/* u2_1566 Output nets */
wire t_4594,   t_4595,   t_4596;
/* u2_1567 Output nets */
wire t_4597,   t_4598,   t_4599;
/* u2_1568 Output nets */
wire t_4600,   t_4601,   t_4602;
/* u2_1569 Output nets */
wire t_4603,   t_4604,   t_4605;
/* u0_1570 Output nets */
wire t_4606,   t_4607;
/* u2_1571 Output nets */
wire t_4608,   t_4609,   t_4610;
/* u2_1572 Output nets */
wire t_4611,   t_4612,   t_4613;
/* u2_1573 Output nets */
wire t_4614,   t_4615,   t_4616;
/* u2_1574 Output nets */
wire t_4617,   t_4618,   t_4619;
/* u2_1575 Output nets */
wire t_4620,   t_4621,   t_4622;
/* u2_1576 Output nets */
wire t_4623,   t_4624,   t_4625;
/* u2_1577 Output nets */
wire t_4626,   t_4627,   t_4628;
/* u2_1578 Output nets */
wire t_4629,   t_4630,   t_4631;
/* u2_1579 Output nets */
wire t_4632,   t_4633,   t_4634;
/* u2_1580 Output nets */
wire t_4635,   t_4636,   t_4637;
/* u2_1581 Output nets */
wire t_4638,   t_4639,   t_4640;
/* u2_1582 Output nets */
wire t_4641,   t_4642,   t_4643;
/* u0_1583 Output nets */
wire t_4644,   t_4645;
/* u2_1584 Output nets */
wire t_4646,   t_4647,   t_4648;
/* u2_1585 Output nets */
wire t_4649,   t_4650,   t_4651;
/* u2_1586 Output nets */
wire t_4652,   t_4653,   t_4654;
/* u2_1587 Output nets */
wire t_4655,   t_4656,   t_4657;
/* u2_1588 Output nets */
wire t_4658,   t_4659,   t_4660;
/* u2_1589 Output nets */
wire t_4661,   t_4662,   t_4663;
/* u2_1590 Output nets */
wire t_4664,   t_4665,   t_4666;
/* u2_1591 Output nets */
wire t_4667,   t_4668,   t_4669;
/* u2_1592 Output nets */
wire t_4670,   t_4671,   t_4672;
/* u2_1593 Output nets */
wire t_4673,   t_4674,   t_4675;
/* u2_1594 Output nets */
wire t_4676,   t_4677,   t_4678;
/* u2_1595 Output nets */
wire t_4679,   t_4680,   t_4681;
/* u2_1596 Output nets */
wire t_4682,   t_4683,   t_4684;
/* u2_1597 Output nets */
wire t_4685,   t_4686,   t_4687;
/* u2_1598 Output nets */
wire t_4688,   t_4689,   t_4690;
/* u2_1599 Output nets */
wire t_4691,   t_4692,   t_4693;
/* u2_1600 Output nets */
wire t_4694,   t_4695,   t_4696;
/* u2_1601 Output nets */
wire t_4697,   t_4698,   t_4699;
/* u2_1602 Output nets */
wire t_4700,   t_4701,   t_4702;
/* u2_1603 Output nets */
wire t_4703,   t_4704,   t_4705;
/* u2_1604 Output nets */
wire t_4706,   t_4707,   t_4708;
/* u2_1605 Output nets */
wire t_4709,   t_4710,   t_4711;
/* u2_1606 Output nets */
wire t_4712,   t_4713,   t_4714;
/* u2_1607 Output nets */
wire t_4715,   t_4716,   t_4717;
/* u2_1608 Output nets */
wire t_4718,   t_4719,   t_4720;
/* u2_1609 Output nets */
wire t_4721,   t_4722,   t_4723;
/* u2_1610 Output nets */
wire t_4724,   t_4725,   t_4726;
/* u2_1611 Output nets */
wire t_4727,   t_4728,   t_4729;
/* u2_1612 Output nets */
wire t_4730,   t_4731,   t_4732;
/* u2_1613 Output nets */
wire t_4733,   t_4734,   t_4735;
/* u2_1614 Output nets */
wire t_4736,   t_4737,   t_4738;
/* u2_1615 Output nets */
wire t_4739,   t_4740,   t_4741;
/* u2_1616 Output nets */
wire t_4742,   t_4743,   t_4744;
/* u2_1617 Output nets */
wire t_4745,   t_4746,   t_4747;
/* u2_1618 Output nets */
wire t_4748,   t_4749,   t_4750;
/* u1_1619 Output nets */
wire t_4751,   t_4752;
/* u2_1620 Output nets */
wire t_4753,   t_4754,   t_4755;
/* u2_1621 Output nets */
wire t_4756,   t_4757,   t_4758;
/* u2_1622 Output nets */
wire t_4759,   t_4760,   t_4761;
/* u2_1623 Output nets */
wire t_4762,   t_4763,   t_4764;
/* u2_1624 Output nets */
wire t_4765,   t_4766,   t_4767;
/* u2_1625 Output nets */
wire t_4768,   t_4769,   t_4770;
/* u2_1626 Output nets */
wire t_4771,   t_4772,   t_4773;
/* u2_1627 Output nets */
wire t_4774,   t_4775,   t_4776;
/* u2_1628 Output nets */
wire t_4777,   t_4778,   t_4779;
/* u2_1629 Output nets */
wire t_4780,   t_4781,   t_4782;
/* u2_1630 Output nets */
wire t_4783,   t_4784,   t_4785;
/* u1_1631 Output nets */
wire t_4786,   t_4787;
/* u2_1632 Output nets */
wire t_4788,   t_4789,   t_4790;
/* u2_1633 Output nets */
wire t_4791,   t_4792,   t_4793;
/* u2_1634 Output nets */
wire t_4794,   t_4795,   t_4796;
/* u2_1635 Output nets */
wire t_4797,   t_4798,   t_4799;
/* u2_1636 Output nets */
wire t_4800,   t_4801,   t_4802;
/* u2_1637 Output nets */
wire t_4803,   t_4804,   t_4805;
/* u2_1638 Output nets */
wire t_4806,   t_4807,   t_4808;
/* u2_1639 Output nets */
wire t_4809,   t_4810,   t_4811;
/* u2_1640 Output nets */
wire t_4812,   t_4813,   t_4814;
/* u2_1641 Output nets */
wire t_4815,   t_4816,   t_4817;
/* u2_1642 Output nets */
wire t_4818,   t_4819,   t_4820;
/* u1_1643 Output nets */
wire t_4821,   t_4822;
/* u2_1644 Output nets */
wire t_4823,   t_4824,   t_4825;
/* u2_1645 Output nets */
wire t_4826,   t_4827,   t_4828;
/* u2_1646 Output nets */
wire t_4829,   t_4830,   t_4831;
/* u2_1647 Output nets */
wire t_4832,   t_4833,   t_4834;
/* u2_1648 Output nets */
wire t_4835,   t_4836,   t_4837;
/* u2_1649 Output nets */
wire t_4838,   t_4839,   t_4840;
/* u2_1650 Output nets */
wire t_4841,   t_4842,   t_4843;
/* u2_1651 Output nets */
wire t_4844,   t_4845,   t_4846;
/* u2_1652 Output nets */
wire t_4847,   t_4848,   t_4849;
/* u2_1653 Output nets */
wire t_4850,   t_4851,   t_4852;
/* u2_1654 Output nets */
wire t_4853,   t_4854,   t_4855;
/* u1_1655 Output nets */
wire t_4856,   t_4857;
/* u2_1656 Output nets */
wire t_4858,   t_4859,   t_4860;
/* u2_1657 Output nets */
wire t_4861,   t_4862,   t_4863;
/* u2_1658 Output nets */
wire t_4864,   t_4865,   t_4866;
/* u2_1659 Output nets */
wire t_4867,   t_4868,   t_4869;
/* u2_1660 Output nets */
wire t_4870,   t_4871,   t_4872;
/* u2_1661 Output nets */
wire t_4873,   t_4874,   t_4875;
/* u2_1662 Output nets */
wire t_4876,   t_4877,   t_4878;
/* u2_1663 Output nets */
wire t_4879,   t_4880,   t_4881;
/* u2_1664 Output nets */
wire t_4882,   t_4883,   t_4884;
/* u2_1665 Output nets */
wire t_4885,   t_4886,   t_4887;
/* u2_1666 Output nets */
wire t_4888,   t_4889,   t_4890;
/* u0_1667 Output nets */
wire t_4891,   t_4892;
/* u2_1668 Output nets */
wire t_4893,   t_4894,   t_4895;
/* u2_1669 Output nets */
wire t_4896,   t_4897,   t_4898;
/* u2_1670 Output nets */
wire t_4899,   t_4900,   t_4901;
/* u2_1671 Output nets */
wire t_4902,   t_4903,   t_4904;
/* u2_1672 Output nets */
wire t_4905,   t_4906,   t_4907;
/* u2_1673 Output nets */
wire t_4908,   t_4909,   t_4910;
/* u2_1674 Output nets */
wire t_4911,   t_4912,   t_4913;
/* u2_1675 Output nets */
wire t_4914,   t_4915,   t_4916;
/* u2_1676 Output nets */
wire t_4917,   t_4918,   t_4919;
/* u2_1677 Output nets */
wire t_4920,   t_4921,   t_4922;
/* u2_1678 Output nets */
wire t_4923,   t_4924,   t_4925;
/* u0_1679 Output nets */
wire t_4926,   t_4927;
/* u2_1680 Output nets */
wire t_4928,   t_4929,   t_4930;
/* u2_1681 Output nets */
wire t_4931,   t_4932,   t_4933;
/* u2_1682 Output nets */
wire t_4934,   t_4935,   t_4936;
/* u2_1683 Output nets */
wire t_4937,   t_4938,   t_4939;
/* u2_1684 Output nets */
wire t_4940,   t_4941,   t_4942;
/* u2_1685 Output nets */
wire t_4943,   t_4944,   t_4945;
/* u2_1686 Output nets */
wire t_4946,   t_4947,   t_4948;
/* u2_1687 Output nets */
wire t_4949,   t_4950,   t_4951;
/* u2_1688 Output nets */
wire t_4952,   t_4953,   t_4954;
/* u2_1689 Output nets */
wire t_4955,   t_4956,   t_4957;
/* u2_1690 Output nets */
wire t_4958,   t_4959,   t_4960;
/* u2_1691 Output nets */
wire t_4961,   t_4962,   t_4963;
/* u2_1692 Output nets */
wire t_4964,   t_4965,   t_4966;
/* u2_1693 Output nets */
wire t_4967,   t_4968,   t_4969;
/* u2_1694 Output nets */
wire t_4970,   t_4971,   t_4972;
/* u2_1695 Output nets */
wire t_4973,   t_4974,   t_4975;
/* u2_1696 Output nets */
wire t_4976,   t_4977,   t_4978;
/* u2_1697 Output nets */
wire t_4979,   t_4980,   t_4981;
/* u2_1698 Output nets */
wire t_4982,   t_4983,   t_4984;
/* u2_1699 Output nets */
wire t_4985,   t_4986,   t_4987;
/* u2_1700 Output nets */
wire t_4988,   t_4989,   t_4990;
/* u2_1701 Output nets */
wire t_4991,   t_4992,   t_4993;
/* u2_1702 Output nets */
wire t_4994,   t_4995,   t_4996;
/* u2_1703 Output nets */
wire t_4997,   t_4998,   t_4999;
/* u2_1704 Output nets */
wire t_5000,   t_5001,   t_5002;
/* u2_1705 Output nets */
wire t_5003,   t_5004,   t_5005;
/* u2_1706 Output nets */
wire t_5006,   t_5007,   t_5008;
/* u2_1707 Output nets */
wire t_5009,   t_5010,   t_5011;
/* u2_1708 Output nets */
wire t_5012,   t_5013,   t_5014;
/* u2_1709 Output nets */
wire t_5015,   t_5016,   t_5017;
/* u2_1710 Output nets */
wire t_5018,   t_5019,   t_5020;
/* u2_1711 Output nets */
wire t_5021,   t_5022,   t_5023;
/* u1_1712 Output nets */
wire t_5024,   t_5025;
/* u2_1713 Output nets */
wire t_5026,   t_5027,   t_5028;
/* u2_1714 Output nets */
wire t_5029,   t_5030,   t_5031;
/* u2_1715 Output nets */
wire t_5032,   t_5033,   t_5034;
/* u2_1716 Output nets */
wire t_5035,   t_5036,   t_5037;
/* u2_1717 Output nets */
wire t_5038,   t_5039,   t_5040;
/* u2_1718 Output nets */
wire t_5041,   t_5042,   t_5043;
/* u2_1719 Output nets */
wire t_5044,   t_5045,   t_5046;
/* u2_1720 Output nets */
wire t_5047,   t_5048,   t_5049;
/* u2_1721 Output nets */
wire t_5050,   t_5051,   t_5052;
/* u2_1722 Output nets */
wire t_5053,   t_5054,   t_5055;
/* u1_1723 Output nets */
wire t_5056,   t_5057;
/* u2_1724 Output nets */
wire t_5058,   t_5059,   t_5060;
/* u2_1725 Output nets */
wire t_5061,   t_5062,   t_5063;
/* u2_1726 Output nets */
wire t_5064,   t_5065,   t_5066;
/* u2_1727 Output nets */
wire t_5067,   t_5068,   t_5069;
/* u2_1728 Output nets */
wire t_5070,   t_5071,   t_5072;
/* u2_1729 Output nets */
wire t_5073,   t_5074,   t_5075;
/* u2_1730 Output nets */
wire t_5076,   t_5077,   t_5078;
/* u2_1731 Output nets */
wire t_5079,   t_5080,   t_5081;
/* u2_1732 Output nets */
wire t_5082,   t_5083,   t_5084;
/* u2_1733 Output nets */
wire t_5085,   t_5086,   t_5087;
/* u1_1734 Output nets */
wire t_5088,   t_5089;
/* u2_1735 Output nets */
wire t_5090,   t_5091,   t_5092;
/* u2_1736 Output nets */
wire t_5093,   t_5094,   t_5095;
/* u2_1737 Output nets */
wire t_5096,   t_5097,   t_5098;
/* u2_1738 Output nets */
wire t_5099,   t_5100,   t_5101;
/* u2_1739 Output nets */
wire t_5102,   t_5103,   t_5104;
/* u2_1740 Output nets */
wire t_5105,   t_5106,   t_5107;
/* u2_1741 Output nets */
wire t_5108,   t_5109,   t_5110;
/* u2_1742 Output nets */
wire t_5111,   t_5112,   t_5113;
/* u2_1743 Output nets */
wire t_5114,   t_5115,   t_5116;
/* u2_1744 Output nets */
wire t_5117,   t_5118,   t_5119;
/* u1_1745 Output nets */
wire t_5120,   t_5121;
/* u2_1746 Output nets */
wire t_5122,   t_5123,   t_5124;
/* u2_1747 Output nets */
wire t_5125,   t_5126,   t_5127;
/* u2_1748 Output nets */
wire t_5128,   t_5129,   t_5130;
/* u2_1749 Output nets */
wire t_5131,   t_5132,   t_5133;
/* u2_1750 Output nets */
wire t_5134,   t_5135,   t_5136;
/* u2_1751 Output nets */
wire t_5137,   t_5138,   t_5139;
/* u2_1752 Output nets */
wire t_5140,   t_5141,   t_5142;
/* u2_1753 Output nets */
wire t_5143,   t_5144,   t_5145;
/* u2_1754 Output nets */
wire t_5146,   t_5147,   t_5148;
/* u2_1755 Output nets */
wire t_5149,   t_5150,   t_5151;
/* u0_1756 Output nets */
wire t_5152,   t_5153;
/* u2_1757 Output nets */
wire t_5154,   t_5155,   t_5156;
/* u2_1758 Output nets */
wire t_5157,   t_5158,   t_5159;
/* u2_1759 Output nets */
wire t_5160,   t_5161,   t_5162;
/* u2_1760 Output nets */
wire t_5163,   t_5164,   t_5165;
/* u2_1761 Output nets */
wire t_5166,   t_5167,   t_5168;
/* u2_1762 Output nets */
wire t_5169,   t_5170,   t_5171;
/* u2_1763 Output nets */
wire t_5172,   t_5173,   t_5174;
/* u2_1764 Output nets */
wire t_5175,   t_5176,   t_5177;
/* u2_1765 Output nets */
wire t_5178,   t_5179,   t_5180;
/* u2_1766 Output nets */
wire t_5181,   t_5182,   t_5183;
/* u0_1767 Output nets */
wire t_5184,   t_5185;
/* u2_1768 Output nets */
wire t_5186,   t_5187,   t_5188;
/* u2_1769 Output nets */
wire t_5189,   t_5190,   t_5191;
/* u2_1770 Output nets */
wire t_5192,   t_5193,   t_5194;
/* u2_1771 Output nets */
wire t_5195,   t_5196,   t_5197;
/* u2_1772 Output nets */
wire t_5198,   t_5199,   t_5200;
/* u2_1773 Output nets */
wire t_5201,   t_5202,   t_5203;
/* u2_1774 Output nets */
wire t_5204,   t_5205,   t_5206;
/* u2_1775 Output nets */
wire t_5207,   t_5208,   t_5209;
/* u2_1776 Output nets */
wire t_5210,   t_5211,   t_5212;
/* u2_1777 Output nets */
wire t_5213,   t_5214,   t_5215;
/* u2_1778 Output nets */
wire t_5216,   t_5217,   t_5218;
/* u2_1779 Output nets */
wire t_5219,   t_5220,   t_5221;
/* u2_1780 Output nets */
wire t_5222,   t_5223,   t_5224;
/* u2_1781 Output nets */
wire t_5225,   t_5226,   t_5227;
/* u2_1782 Output nets */
wire t_5228,   t_5229,   t_5230;
/* u2_1783 Output nets */
wire t_5231,   t_5232,   t_5233;
/* u2_1784 Output nets */
wire t_5234,   t_5235,   t_5236;
/* u2_1785 Output nets */
wire t_5237,   t_5238,   t_5239;
/* u2_1786 Output nets */
wire t_5240,   t_5241,   t_5242;
/* u2_1787 Output nets */
wire t_5243,   t_5244,   t_5245;
/* u2_1788 Output nets */
wire t_5246,   t_5247,   t_5248;
/* u2_1789 Output nets */
wire t_5249,   t_5250,   t_5251;
/* u2_1790 Output nets */
wire t_5252,   t_5253,   t_5254;
/* u2_1791 Output nets */
wire t_5255,   t_5256,   t_5257;
/* u2_1792 Output nets */
wire t_5258,   t_5259,   t_5260;
/* u2_1793 Output nets */
wire t_5261,   t_5262,   t_5263;
/* u2_1794 Output nets */
wire t_5264,   t_5265,   t_5266;
/* u2_1795 Output nets */
wire t_5267,   t_5268,   t_5269;
/* u2_1796 Output nets */
wire t_5270,   t_5271,   t_5272;
/* u1_1797 Output nets */
wire t_5273,   t_5274;
/* u2_1798 Output nets */
wire t_5275,   t_5276,   t_5277;
/* u2_1799 Output nets */
wire t_5278,   t_5279,   t_5280;
/* u2_1800 Output nets */
wire t_5281,   t_5282,   t_5283;
/* u2_1801 Output nets */
wire t_5284,   t_5285,   t_5286;
/* u2_1802 Output nets */
wire t_5287,   t_5288,   t_5289;
/* u2_1803 Output nets */
wire t_5290,   t_5291,   t_5292;
/* u2_1804 Output nets */
wire t_5293,   t_5294,   t_5295;
/* u2_1805 Output nets */
wire t_5296,   t_5297,   t_5298;
/* u2_1806 Output nets */
wire t_5299,   t_5300,   t_5301;
/* u1_1807 Output nets */
wire t_5302,   t_5303;
/* u2_1808 Output nets */
wire t_5304,   t_5305,   t_5306;
/* u2_1809 Output nets */
wire t_5307,   t_5308,   t_5309;
/* u2_1810 Output nets */
wire t_5310,   t_5311,   t_5312;
/* u2_1811 Output nets */
wire t_5313,   t_5314,   t_5315;
/* u2_1812 Output nets */
wire t_5316,   t_5317,   t_5318;
/* u2_1813 Output nets */
wire t_5319,   t_5320,   t_5321;
/* u2_1814 Output nets */
wire t_5322,   t_5323,   t_5324;
/* u2_1815 Output nets */
wire t_5325,   t_5326,   t_5327;
/* u2_1816 Output nets */
wire t_5328,   t_5329,   t_5330;
/* u1_1817 Output nets */
wire t_5331,   t_5332;
/* u2_1818 Output nets */
wire t_5333,   t_5334,   t_5335;
/* u2_1819 Output nets */
wire t_5336,   t_5337,   t_5338;
/* u2_1820 Output nets */
wire t_5339,   t_5340,   t_5341;
/* u2_1821 Output nets */
wire t_5342,   t_5343,   t_5344;
/* u2_1822 Output nets */
wire t_5345,   t_5346,   t_5347;
/* u2_1823 Output nets */
wire t_5348,   t_5349,   t_5350;
/* u2_1824 Output nets */
wire t_5351,   t_5352,   t_5353;
/* u2_1825 Output nets */
wire t_5354,   t_5355,   t_5356;
/* u2_1826 Output nets */
wire t_5357,   t_5358,   t_5359;
/* u1_1827 Output nets */
wire t_5360,   t_5361;
/* u2_1828 Output nets */
wire t_5362,   t_5363,   t_5364;
/* u2_1829 Output nets */
wire t_5365,   t_5366,   t_5367;
/* u2_1830 Output nets */
wire t_5368,   t_5369,   t_5370;
/* u2_1831 Output nets */
wire t_5371,   t_5372,   t_5373;
/* u2_1832 Output nets */
wire t_5374,   t_5375,   t_5376;
/* u2_1833 Output nets */
wire t_5377,   t_5378,   t_5379;
/* u2_1834 Output nets */
wire t_5380,   t_5381,   t_5382;
/* u2_1835 Output nets */
wire t_5383,   t_5384,   t_5385;
/* u2_1836 Output nets */
wire t_5386,   t_5387,   t_5388;
/* u0_1837 Output nets */
wire t_5389,   t_5390;
/* u2_1838 Output nets */
wire t_5391,   t_5392,   t_5393;
/* u2_1839 Output nets */
wire t_5394,   t_5395,   t_5396;
/* u2_1840 Output nets */
wire t_5397,   t_5398,   t_5399;
/* u2_1841 Output nets */
wire t_5400,   t_5401,   t_5402;
/* u2_1842 Output nets */
wire t_5403,   t_5404,   t_5405;
/* u2_1843 Output nets */
wire t_5406,   t_5407,   t_5408;
/* u2_1844 Output nets */
wire t_5409,   t_5410,   t_5411;
/* u2_1845 Output nets */
wire t_5412,   t_5413,   t_5414;
/* u2_1846 Output nets */
wire t_5415,   t_5416,   t_5417;
/* u0_1847 Output nets */
wire t_5418,   t_5419;
/* u2_1848 Output nets */
wire t_5420,   t_5421,   t_5422;
/* u2_1849 Output nets */
wire t_5423,   t_5424,   t_5425;
/* u2_1850 Output nets */
wire t_5426,   t_5427,   t_5428;
/* u2_1851 Output nets */
wire t_5429,   t_5430,   t_5431;
/* u2_1852 Output nets */
wire t_5432,   t_5433,   t_5434;
/* u2_1853 Output nets */
wire t_5435,   t_5436,   t_5437;
/* u2_1854 Output nets */
wire t_5438,   t_5439,   t_5440;
/* u2_1855 Output nets */
wire t_5441,   t_5442,   t_5443;
/* u2_1856 Output nets */
wire t_5444,   t_5445,   t_5446;
/* u2_1857 Output nets */
wire t_5447,   t_5448,   t_5449;
/* u2_1858 Output nets */
wire t_5450,   t_5451,   t_5452;
/* u2_1859 Output nets */
wire t_5453,   t_5454,   t_5455;
/* u2_1860 Output nets */
wire t_5456,   t_5457,   t_5458;
/* u2_1861 Output nets */
wire t_5459,   t_5460,   t_5461;
/* u2_1862 Output nets */
wire t_5462,   t_5463,   t_5464;
/* u2_1863 Output nets */
wire t_5465,   t_5466,   t_5467;
/* u2_1864 Output nets */
wire t_5468,   t_5469,   t_5470;
/* u2_1865 Output nets */
wire t_5471,   t_5472,   t_5473;
/* u2_1866 Output nets */
wire t_5474,   t_5475,   t_5476;
/* u2_1867 Output nets */
wire t_5477,   t_5478,   t_5479;
/* u2_1868 Output nets */
wire t_5480,   t_5481,   t_5482;
/* u2_1869 Output nets */
wire t_5483,   t_5484,   t_5485;
/* u2_1870 Output nets */
wire t_5486,   t_5487,   t_5488;
/* u2_1871 Output nets */
wire t_5489,   t_5490,   t_5491;
/* u2_1872 Output nets */
wire t_5492,   t_5493,   t_5494;
/* u2_1873 Output nets */
wire t_5495,   t_5496,   t_5497;
/* u1_1874 Output nets */
wire t_5498,   t_5499;
/* u2_1875 Output nets */
wire t_5500,   t_5501,   t_5502;
/* u2_1876 Output nets */
wire t_5503,   t_5504,   t_5505;
/* u2_1877 Output nets */
wire t_5506,   t_5507,   t_5508;
/* u2_1878 Output nets */
wire t_5509,   t_5510,   t_5511;
/* u2_1879 Output nets */
wire t_5512,   t_5513,   t_5514;
/* u2_1880 Output nets */
wire t_5515,   t_5516,   t_5517;
/* u2_1881 Output nets */
wire t_5518,   t_5519,   t_5520;
/* u2_1882 Output nets */
wire t_5521,   t_5522,   t_5523;
/* u1_1883 Output nets */
wire t_5524,   t_5525;
/* u2_1884 Output nets */
wire t_5526,   t_5527,   t_5528;
/* u2_1885 Output nets */
wire t_5529,   t_5530,   t_5531;
/* u2_1886 Output nets */
wire t_5532,   t_5533,   t_5534;
/* u2_1887 Output nets */
wire t_5535,   t_5536,   t_5537;
/* u2_1888 Output nets */
wire t_5538,   t_5539,   t_5540;
/* u2_1889 Output nets */
wire t_5541,   t_5542,   t_5543;
/* u2_1890 Output nets */
wire t_5544,   t_5545,   t_5546;
/* u2_1891 Output nets */
wire t_5547,   t_5548,   t_5549;
/* u1_1892 Output nets */
wire t_5550,   t_5551;
/* u2_1893 Output nets */
wire t_5552,   t_5553,   t_5554;
/* u2_1894 Output nets */
wire t_5555,   t_5556,   t_5557;
/* u2_1895 Output nets */
wire t_5558,   t_5559,   t_5560;
/* u2_1896 Output nets */
wire t_5561,   t_5562,   t_5563;
/* u2_1897 Output nets */
wire t_5564,   t_5565,   t_5566;
/* u2_1898 Output nets */
wire t_5567,   t_5568,   t_5569;
/* u2_1899 Output nets */
wire t_5570,   t_5571,   t_5572;
/* u2_1900 Output nets */
wire t_5573,   t_5574,   t_5575;
/* u1_1901 Output nets */
wire t_5576,   t_5577;
/* u2_1902 Output nets */
wire t_5578,   t_5579,   t_5580;
/* u2_1903 Output nets */
wire t_5581,   t_5582,   t_5583;
/* u2_1904 Output nets */
wire t_5584,   t_5585,   t_5586;
/* u2_1905 Output nets */
wire t_5587,   t_5588,   t_5589;
/* u2_1906 Output nets */
wire t_5590,   t_5591,   t_5592;
/* u2_1907 Output nets */
wire t_5593,   t_5594,   t_5595;
/* u2_1908 Output nets */
wire t_5596,   t_5597,   t_5598;
/* u2_1909 Output nets */
wire t_5599,   t_5600,   t_5601;
/* u0_1910 Output nets */
wire t_5602,   t_5603;
/* u2_1911 Output nets */
wire t_5604,   t_5605,   t_5606;
/* u2_1912 Output nets */
wire t_5607,   t_5608,   t_5609;
/* u2_1913 Output nets */
wire t_5610,   t_5611,   t_5612;
/* u2_1914 Output nets */
wire t_5613,   t_5614,   t_5615;
/* u2_1915 Output nets */
wire t_5616,   t_5617,   t_5618;
/* u2_1916 Output nets */
wire t_5619,   t_5620,   t_5621;
/* u2_1917 Output nets */
wire t_5622,   t_5623,   t_5624;
/* u2_1918 Output nets */
wire t_5625,   t_5626,   t_5627;
/* u0_1919 Output nets */
wire t_5628,   t_5629;
/* u2_1920 Output nets */
wire t_5630,   t_5631,   t_5632;
/* u2_1921 Output nets */
wire t_5633,   t_5634,   t_5635;
/* u2_1922 Output nets */
wire t_5636,   t_5637,   t_5638;
/* u2_1923 Output nets */
wire t_5639,   t_5640,   t_5641;
/* u2_1924 Output nets */
wire t_5642,   t_5643,   t_5644;
/* u2_1925 Output nets */
wire t_5645,   t_5646,   t_5647;
/* u2_1926 Output nets */
wire t_5648,   t_5649,   t_5650;
/* u2_1927 Output nets */
wire t_5651,   t_5652,   t_5653;
/* u2_1928 Output nets */
wire t_5654,   t_5655,   t_5656;
/* u2_1929 Output nets */
wire t_5657,   t_5658,   t_5659;
/* u2_1930 Output nets */
wire t_5660,   t_5661,   t_5662;
/* u2_1931 Output nets */
wire t_5663,   t_5664,   t_5665;
/* u2_1932 Output nets */
wire t_5666,   t_5667,   t_5668;
/* u2_1933 Output nets */
wire t_5669,   t_5670,   t_5671;
/* u2_1934 Output nets */
wire t_5672,   t_5673,   t_5674;
/* u2_1935 Output nets */
wire t_5675,   t_5676,   t_5677;
/* u2_1936 Output nets */
wire t_5678,   t_5679,   t_5680;
/* u2_1937 Output nets */
wire t_5681,   t_5682,   t_5683;
/* u2_1938 Output nets */
wire t_5684,   t_5685,   t_5686;
/* u2_1939 Output nets */
wire t_5687,   t_5688,   t_5689;
/* u2_1940 Output nets */
wire t_5690,   t_5691,   t_5692;
/* u2_1941 Output nets */
wire t_5693,   t_5694,   t_5695;
/* u2_1942 Output nets */
wire t_5696,   t_5697,   t_5698;
/* u1_1943 Output nets */
wire t_5699,   t_5700;
/* u2_1944 Output nets */
wire t_5701,   t_5702,   t_5703;
/* u2_1945 Output nets */
wire t_5704,   t_5705,   t_5706;
/* u2_1946 Output nets */
wire t_5707,   t_5708,   t_5709;
/* u2_1947 Output nets */
wire t_5710,   t_5711,   t_5712;
/* u2_1948 Output nets */
wire t_5713,   t_5714,   t_5715;
/* u2_1949 Output nets */
wire t_5716,   t_5717,   t_5718;
/* u2_1950 Output nets */
wire t_5719,   t_5720,   t_5721;
/* u1_1951 Output nets */
wire t_5722,   t_5723;
/* u2_1952 Output nets */
wire t_5724,   t_5725,   t_5726;
/* u2_1953 Output nets */
wire t_5727,   t_5728,   t_5729;
/* u2_1954 Output nets */
wire t_5730,   t_5731,   t_5732;
/* u2_1955 Output nets */
wire t_5733,   t_5734,   t_5735;
/* u2_1956 Output nets */
wire t_5736,   t_5737,   t_5738;
/* u2_1957 Output nets */
wire t_5739,   t_5740,   t_5741;
/* u2_1958 Output nets */
wire t_5742,   t_5743,   t_5744;
/* u1_1959 Output nets */
wire t_5745,   t_5746;
/* u2_1960 Output nets */
wire t_5747,   t_5748,   t_5749;
/* u2_1961 Output nets */
wire t_5750,   t_5751,   t_5752;
/* u2_1962 Output nets */
wire t_5753,   t_5754,   t_5755;
/* u2_1963 Output nets */
wire t_5756,   t_5757,   t_5758;
/* u2_1964 Output nets */
wire t_5759,   t_5760,   t_5761;
/* u2_1965 Output nets */
wire t_5762,   t_5763,   t_5764;
/* u2_1966 Output nets */
wire t_5765,   t_5766,   t_5767;
/* u1_1967 Output nets */
wire t_5768,   t_5769;
/* u2_1968 Output nets */
wire t_5770,   t_5771,   t_5772;
/* u2_1969 Output nets */
wire t_5773,   t_5774,   t_5775;
/* u2_1970 Output nets */
wire t_5776,   t_5777,   t_5778;
/* u2_1971 Output nets */
wire t_5779,   t_5780,   t_5781;
/* u2_1972 Output nets */
wire t_5782,   t_5783,   t_5784;
/* u2_1973 Output nets */
wire t_5785,   t_5786,   t_5787;
/* u2_1974 Output nets */
wire t_5788,   t_5789,   t_5790;
/* u0_1975 Output nets */
wire t_5791,   t_5792;
/* u2_1976 Output nets */
wire t_5793,   t_5794,   t_5795;
/* u2_1977 Output nets */
wire t_5796,   t_5797,   t_5798;
/* u2_1978 Output nets */
wire t_5799,   t_5800,   t_5801;
/* u2_1979 Output nets */
wire t_5802,   t_5803,   t_5804;
/* u2_1980 Output nets */
wire t_5805,   t_5806,   t_5807;
/* u2_1981 Output nets */
wire t_5808,   t_5809,   t_5810;
/* u2_1982 Output nets */
wire t_5811,   t_5812,   t_5813;
/* u0_1983 Output nets */
wire t_5814,   t_5815;
/* u2_1984 Output nets */
wire t_5816,   t_5817,   t_5818;
/* u2_1985 Output nets */
wire t_5819,   t_5820,   t_5821;
/* u2_1986 Output nets */
wire t_5822,   t_5823,   t_5824;
/* u2_1987 Output nets */
wire t_5825,   t_5826,   t_5827;
/* u2_1988 Output nets */
wire t_5828,   t_5829,   t_5830;
/* u2_1989 Output nets */
wire t_5831,   t_5832,   t_5833;
/* u2_1990 Output nets */
wire t_5834,   t_5835,   t_5836;
/* u2_1991 Output nets */
wire t_5837,   t_5838,   t_5839;
/* u2_1992 Output nets */
wire t_5840,   t_5841,   t_5842;
/* u2_1993 Output nets */
wire t_5843,   t_5844,   t_5845;
/* u2_1994 Output nets */
wire t_5846,   t_5847,   t_5848;
/* u2_1995 Output nets */
wire t_5849,   t_5850,   t_5851;
/* u2_1996 Output nets */
wire t_5852,   t_5853,   t_5854;
/* u2_1997 Output nets */
wire t_5855,   t_5856,   t_5857;
/* u2_1998 Output nets */
wire t_5858,   t_5859,   t_5860;
/* u2_1999 Output nets */
wire t_5861,   t_5862,   t_5863;
/* u2_2000 Output nets */
wire t_5864,   t_5865,   t_5866;
/* u2_2001 Output nets */
wire t_5867,   t_5868,   t_5869;
/* u2_2002 Output nets */
wire t_5870,   t_5871,   t_5872;
/* u2_2003 Output nets */
wire t_5873,   t_5874,   t_5875;
/* u1_2004 Output nets */
wire t_5876,   t_5877;
/* u2_2005 Output nets */
wire t_5878,   t_5879,   t_5880;
/* u2_2006 Output nets */
wire t_5881,   t_5882,   t_5883;
/* u2_2007 Output nets */
wire t_5884,   t_5885,   t_5886;
/* u2_2008 Output nets */
wire t_5887,   t_5888,   t_5889;
/* u2_2009 Output nets */
wire t_5890,   t_5891,   t_5892;
/* u2_2010 Output nets */
wire t_5893,   t_5894,   t_5895;
/* u1_2011 Output nets */
wire t_5896,   t_5897;
/* u2_2012 Output nets */
wire t_5898,   t_5899,   t_5900;
/* u2_2013 Output nets */
wire t_5901,   t_5902,   t_5903;
/* u2_2014 Output nets */
wire t_5904,   t_5905,   t_5906;
/* u2_2015 Output nets */
wire t_5907,   t_5908,   t_5909;
/* u2_2016 Output nets */
wire t_5910,   t_5911,   t_5912;
/* u2_2017 Output nets */
wire t_5913,   t_5914,   t_5915;
/* u1_2018 Output nets */
wire t_5916,   t_5917;
/* u2_2019 Output nets */
wire t_5918,   t_5919,   t_5920;
/* u2_2020 Output nets */
wire t_5921,   t_5922,   t_5923;
/* u2_2021 Output nets */
wire t_5924,   t_5925,   t_5926;
/* u2_2022 Output nets */
wire t_5927,   t_5928,   t_5929;
/* u2_2023 Output nets */
wire t_5930,   t_5931,   t_5932;
/* u2_2024 Output nets */
wire t_5933,   t_5934,   t_5935;
/* u1_2025 Output nets */
wire t_5936,   t_5937;
/* u2_2026 Output nets */
wire t_5938,   t_5939,   t_5940;
/* u2_2027 Output nets */
wire t_5941,   t_5942,   t_5943;
/* u2_2028 Output nets */
wire t_5944,   t_5945,   t_5946;
/* u2_2029 Output nets */
wire t_5947,   t_5948,   t_5949;
/* u2_2030 Output nets */
wire t_5950,   t_5951,   t_5952;
/* u2_2031 Output nets */
wire t_5953,   t_5954,   t_5955;
/* u0_2032 Output nets */
wire t_5956,   t_5957;
/* u2_2033 Output nets */
wire t_5958,   t_5959,   t_5960;
/* u2_2034 Output nets */
wire t_5961,   t_5962,   t_5963;
/* u2_2035 Output nets */
wire t_5964,   t_5965,   t_5966;
/* u2_2036 Output nets */
wire t_5967,   t_5968,   t_5969;
/* u2_2037 Output nets */
wire t_5970,   t_5971,   t_5972;
/* u2_2038 Output nets */
wire t_5973,   t_5974,   t_5975;
/* u0_2039 Output nets */
wire t_5976,   t_5977;
/* u2_2040 Output nets */
wire t_5978,   t_5979,   t_5980;
/* u2_2041 Output nets */
wire t_5981,   t_5982,   t_5983;
/* u2_2042 Output nets */
wire t_5984,   t_5985,   t_5986;
/* u2_2043 Output nets */
wire t_5987,   t_5988,   t_5989;
/* u2_2044 Output nets */
wire t_5990,   t_5991,   t_5992;
/* u2_2045 Output nets */
wire t_5993,   t_5994,   t_5995;
/* u2_2046 Output nets */
wire t_5996,   t_5997,   t_5998;
/* u2_2047 Output nets */
wire t_5999,   t_6000,   t_6001;
/* u2_2048 Output nets */
wire t_6002,   t_6003,   t_6004;
/* u2_2049 Output nets */
wire t_6005,   t_6006,   t_6007;
/* u2_2050 Output nets */
wire t_6008,   t_6009,   t_6010;
/* u2_2051 Output nets */
wire t_6011,   t_6012,   t_6013;
/* u2_2052 Output nets */
wire t_6014,   t_6015,   t_6016;
/* u2_2053 Output nets */
wire t_6017,   t_6018,   t_6019;
/* u2_2054 Output nets */
wire t_6020,   t_6021,   t_6022;
/* u2_2055 Output nets */
wire t_6023,   t_6024,   t_6025;
/* u2_2056 Output nets */
wire t_6026,   t_6027,   t_6028;
/* u1_2057 Output nets */
wire t_6029,   t_6030;
/* u2_2058 Output nets */
wire t_6031,   t_6032,   t_6033;
/* u2_2059 Output nets */
wire t_6034,   t_6035,   t_6036;
/* u2_2060 Output nets */
wire t_6037,   t_6038,   t_6039;
/* u2_2061 Output nets */
wire t_6040,   t_6041,   t_6042;
/* u2_2062 Output nets */
wire t_6043,   t_6044,   t_6045;
/* u1_2063 Output nets */
wire t_6046,   t_6047;
/* u2_2064 Output nets */
wire t_6048,   t_6049,   t_6050;
/* u2_2065 Output nets */
wire t_6051,   t_6052,   t_6053;
/* u2_2066 Output nets */
wire t_6054,   t_6055,   t_6056;
/* u2_2067 Output nets */
wire t_6057,   t_6058,   t_6059;
/* u2_2068 Output nets */
wire t_6060,   t_6061,   t_6062;
/* u1_2069 Output nets */
wire t_6063,   t_6064;
/* u2_2070 Output nets */
wire t_6065,   t_6066,   t_6067;
/* u2_2071 Output nets */
wire t_6068,   t_6069,   t_6070;
/* u2_2072 Output nets */
wire t_6071,   t_6072,   t_6073;
/* u2_2073 Output nets */
wire t_6074,   t_6075,   t_6076;
/* u2_2074 Output nets */
wire t_6077,   t_6078,   t_6079;
/* u1_2075 Output nets */
wire t_6080,   t_6081;
/* u2_2076 Output nets */
wire t_6082,   t_6083,   t_6084;
/* u2_2077 Output nets */
wire t_6085,   t_6086,   t_6087;
/* u2_2078 Output nets */
wire t_6088,   t_6089,   t_6090;
/* u2_2079 Output nets */
wire t_6091,   t_6092,   t_6093;
/* u2_2080 Output nets */
wire t_6094,   t_6095,   t_6096;
/* u0_2081 Output nets */
wire t_6097,   t_6098;
/* u2_2082 Output nets */
wire t_6099,   t_6100,   t_6101;
/* u2_2083 Output nets */
wire t_6102,   t_6103,   t_6104;
/* u2_2084 Output nets */
wire t_6105,   t_6106,   t_6107;
/* u2_2085 Output nets */
wire t_6108,   t_6109,   t_6110;
/* u2_2086 Output nets */
wire t_6111,   t_6112,   t_6113;
/* u0_2087 Output nets */
wire t_6114,   t_6115;
/* u2_2088 Output nets */
wire t_6116,   t_6117,   t_6118;
/* u2_2089 Output nets */
wire t_6119,   t_6120,   t_6121;
/* u2_2090 Output nets */
wire t_6122,   t_6123,   t_6124;
/* u2_2091 Output nets */
wire t_6125,   t_6126,   t_6127;
/* u2_2092 Output nets */
wire t_6128,   t_6129,   t_6130;
/* u2_2093 Output nets */
wire t_6131,   t_6132,   t_6133;
/* u2_2094 Output nets */
wire t_6134,   t_6135,   t_6136;
/* u2_2095 Output nets */
wire t_6137,   t_6138,   t_6139;
/* u2_2096 Output nets */
wire t_6140,   t_6141,   t_6142;
/* u2_2097 Output nets */
wire t_6143,   t_6144,   t_6145;
/* u2_2098 Output nets */
wire t_6146,   t_6147,   t_6148;
/* u2_2099 Output nets */
wire t_6149,   t_6150,   t_6151;
/* u2_2100 Output nets */
wire t_6152,   t_6153,   t_6154;
/* u2_2101 Output nets */
wire t_6155,   t_6156,   t_6157;
/* u1_2102 Output nets */
wire t_6158,   t_6159;
/* u2_2103 Output nets */
wire t_6160,   t_6161,   t_6162;
/* u2_2104 Output nets */
wire t_6163,   t_6164,   t_6165;
/* u2_2105 Output nets */
wire t_6166,   t_6167,   t_6168;
/* u2_2106 Output nets */
wire t_6169,   t_6170,   t_6171;
/* u1_2107 Output nets */
wire t_6172,   t_6173;
/* u2_2108 Output nets */
wire t_6174,   t_6175,   t_6176;
/* u2_2109 Output nets */
wire t_6177,   t_6178,   t_6179;
/* u2_2110 Output nets */
wire t_6180,   t_6181,   t_6182;
/* u2_2111 Output nets */
wire t_6183,   t_6184,   t_6185;
/* u1_2112 Output nets */
wire t_6186,   t_6187;
/* u2_2113 Output nets */
wire t_6188,   t_6189,   t_6190;
/* u2_2114 Output nets */
wire t_6191,   t_6192,   t_6193;
/* u2_2115 Output nets */
wire t_6194,   t_6195,   t_6196;
/* u2_2116 Output nets */
wire t_6197,   t_6198,   t_6199;
/* u1_2117 Output nets */
wire t_6200,   t_6201;
/* u2_2118 Output nets */
wire t_6202,   t_6203,   t_6204;
/* u2_2119 Output nets */
wire t_6205,   t_6206,   t_6207;
/* u2_2120 Output nets */
wire t_6208,   t_6209,   t_6210;
/* u2_2121 Output nets */
wire t_6211,   t_6212,   t_6213;
/* u0_2122 Output nets */
wire t_6214,   t_6215;
/* u2_2123 Output nets */
wire t_6216,   t_6217,   t_6218;
/* u2_2124 Output nets */
wire t_6219,   t_6220,   t_6221;
/* u2_2125 Output nets */
wire t_6222,   t_6223,   t_6224;
/* u2_2126 Output nets */
wire t_6225,   t_6226,   t_6227;
/* u0_2127 Output nets */
wire t_6228,   t_6229;
/* u2_2128 Output nets */
wire t_6230,   t_6231,   t_6232;
/* u2_2129 Output nets */
wire t_6233,   t_6234,   t_6235;
/* u2_2130 Output nets */
wire t_6236,   t_6237,   t_6238;
/* u2_2131 Output nets */
wire t_6239,   t_6240,   t_6241;
/* u2_2132 Output nets */
wire t_6242,   t_6243,   t_6244;
/* u2_2133 Output nets */
wire t_6245,   t_6246,   t_6247;
/* u2_2134 Output nets */
wire t_6248,   t_6249,   t_6250;
/* u2_2135 Output nets */
wire t_6251,   t_6252,   t_6253;
/* u2_2136 Output nets */
wire t_6254,   t_6255,   t_6256;
/* u2_2137 Output nets */
wire t_6257,   t_6258,   t_6259;
/* u2_2138 Output nets */
wire t_6260,   t_6261,   t_6262;
/* u1_2139 Output nets */
wire t_6263,   t_6264;
/* u2_2140 Output nets */
wire t_6265,   t_6266,   t_6267;
/* u2_2141 Output nets */
wire t_6268,   t_6269,   t_6270;
/* u2_2142 Output nets */
wire t_6271,   t_6272,   t_6273;
/* u1_2143 Output nets */
wire t_6274,   t_6275;
/* u2_2144 Output nets */
wire t_6276,   t_6277,   t_6278;
/* u2_2145 Output nets */
wire t_6279,   t_6280,   t_6281;
/* u2_2146 Output nets */
wire t_6282,   t_6283,   t_6284;
/* u1_2147 Output nets */
wire t_6285,   t_6286;
/* u2_2148 Output nets */
wire t_6287,   t_6288,   t_6289;
/* u2_2149 Output nets */
wire t_6290,   t_6291,   t_6292;
/* u2_2150 Output nets */
wire t_6293,   t_6294,   t_6295;
/* u1_2151 Output nets */
wire t_6296,   t_6297;
/* u2_2152 Output nets */
wire t_6298,   t_6299,   t_6300;
/* u2_2153 Output nets */
wire t_6301,   t_6302,   t_6303;
/* u2_2154 Output nets */
wire t_6304,   t_6305,   t_6306;
/* u0_2155 Output nets */
wire t_6307,   t_6308;
/* u2_2156 Output nets */
wire t_6309,   t_6310,   t_6311;
/* u2_2157 Output nets */
wire t_6312,   t_6313,   t_6314;
/* u2_2158 Output nets */
wire t_6315,   t_6316,   t_6317;
/* u0_2159 Output nets */
wire t_6318,   t_6319;
/* u2_2160 Output nets */
wire t_6320,   t_6321,   t_6322;
/* u2_2161 Output nets */
wire t_6323,   t_6324,   t_6325;
/* u2_2162 Output nets */
wire t_6326,   t_6327,   t_6328;
/* u2_2163 Output nets */
wire t_6329,   t_6330,   t_6331;
/* u2_2164 Output nets */
wire t_6332,   t_6333,   t_6334;
/* u2_2165 Output nets */
wire t_6335,   t_6336,   t_6337;
/* u2_2166 Output nets */
wire t_6338,   t_6339,   t_6340;
/* u2_2167 Output nets */
wire t_6341,   t_6342,   t_6343;
/* u1_2168 Output nets */
wire t_6344,   t_6345;
/* u2_2169 Output nets */
wire t_6346,   t_6347,   t_6348;
/* u2_2170 Output nets */
wire t_6349,   t_6350,   t_6351;
/* u1_2171 Output nets */
wire t_6352,   t_6353;
/* u2_2172 Output nets */
wire t_6354,   t_6355,   t_6356;
/* u2_2173 Output nets */
wire t_6357,   t_6358,   t_6359;
/* u1_2174 Output nets */
wire t_6360,   t_6361;
/* u2_2175 Output nets */
wire t_6362,   t_6363,   t_6364;
/* u2_2176 Output nets */
wire t_6365,   t_6366,   t_6367;
/* u1_2177 Output nets */
wire t_6368,   t_6369;
/* u2_2178 Output nets */
wire t_6370,   t_6371,   t_6372;
/* u2_2179 Output nets */
wire t_6373,   t_6374,   t_6375;
/* u0_2180 Output nets */
wire t_6376,   t_6377;
/* u2_2181 Output nets */
wire t_6378,   t_6379,   t_6380;
/* u2_2182 Output nets */
wire t_6381,   t_6382,   t_6383;
/* u0_2183 Output nets */
wire t_6384,   t_6385;
/* u2_2184 Output nets */
wire t_6386,   t_6387,   t_6388;
/* u2_2185 Output nets */
wire t_6389,   t_6390,   t_6391;
/* u2_2186 Output nets */
wire t_6392,   t_6393,   t_6394;
/* u2_2187 Output nets */
wire t_6395,   t_6396,   t_6397;
/* u2_2188 Output nets */
wire t_6398,   t_6399,   t_6400;
/* u1_2189 Output nets */
wire t_6401,   t_6402;
/* u2_2190 Output nets */
wire t_6403,   t_6404,   t_6405;
/* u1_2191 Output nets */
wire t_6406,   t_6407;
/* u2_2192 Output nets */
wire t_6408,   t_6409,   t_6410;
/* u1_2193 Output nets */
wire t_6411,   t_6412;
/* u2_2194 Output nets */
wire t_6413,   t_6414,   t_6415;
/* u1_2195 Output nets */
wire t_6416,   t_6417;
/* u2_2196 Output nets */
wire t_6418,   t_6419,   t_6420;
/* u0_2197 Output nets */
wire t_6421,   t_6422;
/* u2_2198 Output nets */
wire t_6423,   t_6424,   t_6425;
/* u0_2199 Output nets */
wire t_6426,   t_6427;
/* u2_2200 Output nets */
wire t_6428,   t_6429,   t_6430;
/* u2_2201 Output nets */
wire t_6431,   t_6432,   t_6433;
/* u1_2202 Output nets */
wire t_6434,   t_6435;
/* u1_2203 Output nets */
wire t_6436,   t_6437;
/* u0_2204 Output nets */
wire t_6438,   t_6439;
/* u0_2205 Output nets */
wire t_6440;

/* compress stage 1 */
half_adder u0_1(.a(s_0_1), .b(s_0_0), .o(t_0), .cout(t_1));
compressor_3_2 u1_2(.a(s_2_2), .b(s_2_1), .cin(s_2_0), .o(t_2), .cout(t_3));
half_adder u0_3(.a(s_3_1), .b(s_3_0), .o(t_4), .cout(t_5));
compressor_4_2 u2_4(.a(s_4_3), .b(s_4_2), .c(s_4_1), .d(s_4_0), .cin(t_5), .o(t_6), .co(t_7), .cout(t_8));
compressor_3_2 u1_5(.a(s_5_1), .b(s_5_0), .cin(t_8), .o(t_9), .cout(t_10));
compressor_4_2 u2_6(.a(s_6_4), .b(s_6_3), .c(s_6_2), .d(s_6_1), .cin(s_6_0), .o(t_11), .co(t_12), .cout(t_13));
compressor_4_2 u2_7(.a(s_7_3), .b(s_7_2), .c(s_7_1), .d(s_7_0), .cin(t_13), .o(t_14), .co(t_15), .cout(t_16));
compressor_4_2 u2_8(.a(s_8_3), .b(s_8_2), .c(s_8_1), .d(s_8_0), .cin(t_16), .o(t_17), .co(t_18), .cout(t_19));
half_adder u0_9(.a(s_8_5), .b(s_8_4), .o(t_20), .cout(t_21));
compressor_4_2 u2_10(.a(s_9_2), .b(s_9_1), .c(s_9_0), .d(t_19), .cin(t_21), .o(t_22), .co(t_23), .cout(t_24));
half_adder u0_11(.a(s_9_4), .b(s_9_3), .o(t_25), .cout(t_26));
compressor_4_2 u2_12(.a(s_10_2), .b(s_10_1), .c(s_10_0), .d(t_24), .cin(t_26), .o(t_27), .co(t_28), .cout(t_29));
compressor_3_2 u1_13(.a(s_10_5), .b(s_10_4), .cin(s_10_3), .o(t_30), .cout(t_31));
compressor_4_2 u2_14(.a(s_11_2), .b(s_11_1), .c(s_11_0), .d(t_29), .cin(t_31), .o(t_32), .co(t_33), .cout(t_34));
compressor_3_2 u1_15(.a(s_11_5), .b(s_11_4), .cin(s_11_3), .o(t_35), .cout(t_36));
compressor_4_2 u2_16(.a(s_12_2), .b(s_12_1), .c(s_12_0), .d(t_34), .cin(t_36), .o(t_37), .co(t_38), .cout(t_39));
compressor_4_2 u2_17(.a(s_12_7), .b(s_12_6), .c(s_12_5), .d(s_12_4), .cin(s_12_3), .o(t_40), .co(t_41), .cout(t_42));
compressor_4_2 u2_18(.a(s_13_2), .b(s_13_1), .c(s_13_0), .d(t_39), .cin(t_42), .o(t_43), .co(t_44), .cout(t_45));
compressor_3_2 u1_19(.a(s_13_5), .b(s_13_4), .cin(s_13_3), .o(t_46), .cout(t_47));
compressor_4_2 u2_20(.a(s_14_2), .b(s_14_1), .c(s_14_0), .d(t_45), .cin(t_47), .o(t_48), .co(t_49), .cout(t_50));
compressor_4_2 u2_21(.a(s_14_7), .b(s_14_6), .c(s_14_5), .d(s_14_4), .cin(s_14_3), .o(t_51), .co(t_52), .cout(t_53));
compressor_4_2 u2_22(.a(s_15_2), .b(s_15_1), .c(s_15_0), .d(t_50), .cin(t_53), .o(t_54), .co(t_55), .cout(t_56));
compressor_4_2 u2_23(.a(s_15_7), .b(s_15_6), .c(s_15_5), .d(s_15_4), .cin(s_15_3), .o(t_57), .co(t_58), .cout(t_59));
compressor_4_2 u2_24(.a(s_16_2), .b(s_16_1), .c(s_16_0), .d(t_56), .cin(t_59), .o(t_60), .co(t_61), .cout(t_62));
compressor_4_2 u2_25(.a(s_16_7), .b(s_16_6), .c(s_16_5), .d(s_16_4), .cin(s_16_3), .o(t_63), .co(t_64), .cout(t_65));
half_adder u0_26(.a(s_16_9), .b(s_16_8), .o(t_66), .cout(t_67));
compressor_4_2 u2_27(.a(s_17_2), .b(s_17_1), .c(s_17_0), .d(t_62), .cin(t_65), .o(t_68), .co(t_69), .cout(t_70));
compressor_4_2 u2_28(.a(s_17_6), .b(s_17_5), .c(s_17_4), .d(s_17_3), .cin(t_67), .o(t_71), .co(t_72), .cout(t_73));
half_adder u0_29(.a(s_17_8), .b(s_17_7), .o(t_74), .cout(t_75));
compressor_4_2 u2_30(.a(s_18_2), .b(s_18_1), .c(s_18_0), .d(t_70), .cin(t_73), .o(t_76), .co(t_77), .cout(t_78));
compressor_4_2 u2_31(.a(s_18_6), .b(s_18_5), .c(s_18_4), .d(s_18_3), .cin(t_75), .o(t_79), .co(t_80), .cout(t_81));
compressor_3_2 u1_32(.a(s_18_9), .b(s_18_8), .cin(s_18_7), .o(t_82), .cout(t_83));
compressor_4_2 u2_33(.a(s_19_2), .b(s_19_1), .c(s_19_0), .d(t_78), .cin(t_81), .o(t_84), .co(t_85), .cout(t_86));
compressor_4_2 u2_34(.a(s_19_6), .b(s_19_5), .c(s_19_4), .d(s_19_3), .cin(t_83), .o(t_87), .co(t_88), .cout(t_89));
compressor_3_2 u1_35(.a(s_19_9), .b(s_19_8), .cin(s_19_7), .o(t_90), .cout(t_91));
compressor_4_2 u2_36(.a(s_20_2), .b(s_20_1), .c(s_20_0), .d(t_86), .cin(t_89), .o(t_92), .co(t_93), .cout(t_94));
compressor_4_2 u2_37(.a(s_20_6), .b(s_20_5), .c(s_20_4), .d(s_20_3), .cin(t_91), .o(t_95), .co(t_96), .cout(t_97));
compressor_4_2 u2_38(.a(s_20_11), .b(s_20_10), .c(s_20_9), .d(s_20_8), .cin(s_20_7), .o(t_98), .co(t_99), .cout(t_100));
compressor_4_2 u2_39(.a(s_21_2), .b(s_21_1), .c(s_21_0), .d(t_94), .cin(t_97), .o(t_101), .co(t_102), .cout(t_103));
compressor_4_2 u2_40(.a(s_21_6), .b(s_21_5), .c(s_21_4), .d(s_21_3), .cin(t_100), .o(t_104), .co(t_105), .cout(t_106));
compressor_3_2 u1_41(.a(s_21_9), .b(s_21_8), .cin(s_21_7), .o(t_107), .cout(t_108));
compressor_4_2 u2_42(.a(s_22_2), .b(s_22_1), .c(s_22_0), .d(t_103), .cin(t_106), .o(t_109), .co(t_110), .cout(t_111));
compressor_4_2 u2_43(.a(s_22_6), .b(s_22_5), .c(s_22_4), .d(s_22_3), .cin(t_108), .o(t_112), .co(t_113), .cout(t_114));
compressor_4_2 u2_44(.a(s_22_11), .b(s_22_10), .c(s_22_9), .d(s_22_8), .cin(s_22_7), .o(t_115), .co(t_116), .cout(t_117));
compressor_4_2 u2_45(.a(s_23_2), .b(s_23_1), .c(s_23_0), .d(t_111), .cin(t_114), .o(t_118), .co(t_119), .cout(t_120));
compressor_4_2 u2_46(.a(s_23_6), .b(s_23_5), .c(s_23_4), .d(s_23_3), .cin(t_117), .o(t_121), .co(t_122), .cout(t_123));
compressor_4_2 u2_47(.a(s_23_11), .b(s_23_10), .c(s_23_9), .d(s_23_8), .cin(s_23_7), .o(t_124), .co(t_125), .cout(t_126));
compressor_4_2 u2_48(.a(s_24_2), .b(s_24_1), .c(s_24_0), .d(t_120), .cin(t_123), .o(t_127), .co(t_128), .cout(t_129));
compressor_4_2 u2_49(.a(s_24_6), .b(s_24_5), .c(s_24_4), .d(s_24_3), .cin(t_126), .o(t_130), .co(t_131), .cout(t_132));
compressor_4_2 u2_50(.a(s_24_11), .b(s_24_10), .c(s_24_9), .d(s_24_8), .cin(s_24_7), .o(t_133), .co(t_134), .cout(t_135));
half_adder u0_51(.a(s_24_13), .b(s_24_12), .o(t_136), .cout(t_137));
compressor_4_2 u2_52(.a(s_25_2), .b(s_25_1), .c(s_25_0), .d(t_129), .cin(t_132), .o(t_138), .co(t_139), .cout(t_140));
compressor_4_2 u2_53(.a(s_25_5), .b(s_25_4), .c(s_25_3), .d(t_135), .cin(t_137), .o(t_141), .co(t_142), .cout(t_143));
compressor_4_2 u2_54(.a(s_25_10), .b(s_25_9), .c(s_25_8), .d(s_25_7), .cin(s_25_6), .o(t_144), .co(t_145), .cout(t_146));
half_adder u0_55(.a(s_25_12), .b(s_25_11), .o(t_147), .cout(t_148));
compressor_4_2 u2_56(.a(s_26_2), .b(s_26_1), .c(s_26_0), .d(t_140), .cin(t_143), .o(t_149), .co(t_150), .cout(t_151));
compressor_4_2 u2_57(.a(s_26_5), .b(s_26_4), .c(s_26_3), .d(t_146), .cin(t_148), .o(t_152), .co(t_153), .cout(t_154));
compressor_4_2 u2_58(.a(s_26_10), .b(s_26_9), .c(s_26_8), .d(s_26_7), .cin(s_26_6), .o(t_155), .co(t_156), .cout(t_157));
compressor_3_2 u1_59(.a(s_26_13), .b(s_26_12), .cin(s_26_11), .o(t_158), .cout(t_159));
compressor_4_2 u2_60(.a(s_27_2), .b(s_27_1), .c(s_27_0), .d(t_151), .cin(t_154), .o(t_160), .co(t_161), .cout(t_162));
compressor_4_2 u2_61(.a(s_27_5), .b(s_27_4), .c(s_27_3), .d(t_157), .cin(t_159), .o(t_163), .co(t_164), .cout(t_165));
compressor_4_2 u2_62(.a(s_27_10), .b(s_27_9), .c(s_27_8), .d(s_27_7), .cin(s_27_6), .o(t_166), .co(t_167), .cout(t_168));
compressor_3_2 u1_63(.a(s_27_13), .b(s_27_12), .cin(s_27_11), .o(t_169), .cout(t_170));
compressor_4_2 u2_64(.a(s_28_2), .b(s_28_1), .c(s_28_0), .d(t_162), .cin(t_165), .o(t_171), .co(t_172), .cout(t_173));
compressor_4_2 u2_65(.a(s_28_5), .b(s_28_4), .c(s_28_3), .d(t_168), .cin(t_170), .o(t_174), .co(t_175), .cout(t_176));
compressor_4_2 u2_66(.a(s_28_10), .b(s_28_9), .c(s_28_8), .d(s_28_7), .cin(s_28_6), .o(t_177), .co(t_178), .cout(t_179));
compressor_4_2 u2_67(.a(s_28_15), .b(s_28_14), .c(s_28_13), .d(s_28_12), .cin(s_28_11), .o(t_180), .co(t_181), .cout(t_182));
compressor_4_2 u2_68(.a(s_29_2), .b(s_29_1), .c(s_29_0), .d(t_173), .cin(t_176), .o(t_183), .co(t_184), .cout(t_185));
compressor_4_2 u2_69(.a(s_29_5), .b(s_29_4), .c(s_29_3), .d(t_179), .cin(t_182), .o(t_186), .co(t_187), .cout(t_188));
compressor_4_2 u2_70(.a(s_29_10), .b(s_29_9), .c(s_29_8), .d(s_29_7), .cin(s_29_6), .o(t_189), .co(t_190), .cout(t_191));
compressor_3_2 u1_71(.a(s_29_13), .b(s_29_12), .cin(s_29_11), .o(t_192), .cout(t_193));
compressor_4_2 u2_72(.a(s_30_2), .b(s_30_1), .c(s_30_0), .d(t_185), .cin(t_188), .o(t_194), .co(t_195), .cout(t_196));
compressor_4_2 u2_73(.a(s_30_5), .b(s_30_4), .c(s_30_3), .d(t_191), .cin(t_193), .o(t_197), .co(t_198), .cout(t_199));
compressor_4_2 u2_74(.a(s_30_10), .b(s_30_9), .c(s_30_8), .d(s_30_7), .cin(s_30_6), .o(t_200), .co(t_201), .cout(t_202));
compressor_4_2 u2_75(.a(s_30_15), .b(s_30_14), .c(s_30_13), .d(s_30_12), .cin(s_30_11), .o(t_203), .co(t_204), .cout(t_205));
compressor_4_2 u2_76(.a(s_31_2), .b(s_31_1), .c(s_31_0), .d(t_196), .cin(t_199), .o(t_206), .co(t_207), .cout(t_208));
compressor_4_2 u2_77(.a(s_31_5), .b(s_31_4), .c(s_31_3), .d(t_202), .cin(t_205), .o(t_209), .co(t_210), .cout(t_211));
compressor_4_2 u2_78(.a(s_31_10), .b(s_31_9), .c(s_31_8), .d(s_31_7), .cin(s_31_6), .o(t_212), .co(t_213), .cout(t_214));
compressor_4_2 u2_79(.a(s_31_15), .b(s_31_14), .c(s_31_13), .d(s_31_12), .cin(s_31_11), .o(t_215), .co(t_216), .cout(t_217));
compressor_4_2 u2_80(.a(s_32_2), .b(s_32_1), .c(s_32_0), .d(t_208), .cin(t_211), .o(t_218), .co(t_219), .cout(t_220));
compressor_4_2 u2_81(.a(s_32_5), .b(s_32_4), .c(s_32_3), .d(t_214), .cin(t_217), .o(t_221), .co(t_222), .cout(t_223));
compressor_4_2 u2_82(.a(s_32_10), .b(s_32_9), .c(s_32_8), .d(s_32_7), .cin(s_32_6), .o(t_224), .co(t_225), .cout(t_226));
compressor_4_2 u2_83(.a(s_32_15), .b(s_32_14), .c(s_32_13), .d(s_32_12), .cin(s_32_11), .o(t_227), .co(t_228), .cout(t_229));
half_adder u0_84(.a(s_32_17), .b(s_32_16), .o(t_230), .cout(t_231));
compressor_4_2 u2_85(.a(s_33_2), .b(s_33_1), .c(s_33_0), .d(t_220), .cin(t_223), .o(t_232), .co(t_233), .cout(t_234));
compressor_4_2 u2_86(.a(s_33_5), .b(s_33_4), .c(s_33_3), .d(t_226), .cin(t_229), .o(t_235), .co(t_236), .cout(t_237));
compressor_4_2 u2_87(.a(s_33_9), .b(s_33_8), .c(s_33_7), .d(s_33_6), .cin(t_231), .o(t_238), .co(t_239), .cout(t_240));
compressor_4_2 u2_88(.a(s_33_14), .b(s_33_13), .c(s_33_12), .d(s_33_11), .cin(s_33_10), .o(t_241), .co(t_242), .cout(t_243));
half_adder u0_89(.a(s_33_16), .b(s_33_15), .o(t_244), .cout(t_245));
compressor_4_2 u2_90(.a(s_34_2), .b(s_34_1), .c(s_34_0), .d(t_234), .cin(t_237), .o(t_246), .co(t_247), .cout(t_248));
compressor_4_2 u2_91(.a(s_34_5), .b(s_34_4), .c(s_34_3), .d(t_240), .cin(t_243), .o(t_249), .co(t_250), .cout(t_251));
compressor_4_2 u2_92(.a(s_34_9), .b(s_34_8), .c(s_34_7), .d(s_34_6), .cin(t_245), .o(t_252), .co(t_253), .cout(t_254));
compressor_4_2 u2_93(.a(s_34_14), .b(s_34_13), .c(s_34_12), .d(s_34_11), .cin(s_34_10), .o(t_255), .co(t_256), .cout(t_257));
compressor_3_2 u1_94(.a(s_34_17), .b(s_34_16), .cin(s_34_15), .o(t_258), .cout(t_259));
compressor_4_2 u2_95(.a(s_35_2), .b(s_35_1), .c(s_35_0), .d(t_248), .cin(t_251), .o(t_260), .co(t_261), .cout(t_262));
compressor_4_2 u2_96(.a(s_35_5), .b(s_35_4), .c(s_35_3), .d(t_254), .cin(t_257), .o(t_263), .co(t_264), .cout(t_265));
compressor_4_2 u2_97(.a(s_35_9), .b(s_35_8), .c(s_35_7), .d(s_35_6), .cin(t_259), .o(t_266), .co(t_267), .cout(t_268));
compressor_4_2 u2_98(.a(s_35_14), .b(s_35_13), .c(s_35_12), .d(s_35_11), .cin(s_35_10), .o(t_269), .co(t_270), .cout(t_271));
compressor_3_2 u1_99(.a(s_35_17), .b(s_35_16), .cin(s_35_15), .o(t_272), .cout(t_273));
compressor_4_2 u2_100(.a(s_36_2), .b(s_36_1), .c(s_36_0), .d(t_262), .cin(t_265), .o(t_274), .co(t_275), .cout(t_276));
compressor_4_2 u2_101(.a(s_36_5), .b(s_36_4), .c(s_36_3), .d(t_268), .cin(t_271), .o(t_277), .co(t_278), .cout(t_279));
compressor_4_2 u2_102(.a(s_36_9), .b(s_36_8), .c(s_36_7), .d(s_36_6), .cin(t_273), .o(t_280), .co(t_281), .cout(t_282));
compressor_4_2 u2_103(.a(s_36_14), .b(s_36_13), .c(s_36_12), .d(s_36_11), .cin(s_36_10), .o(t_283), .co(t_284), .cout(t_285));
compressor_4_2 u2_104(.a(s_36_19), .b(s_36_18), .c(s_36_17), .d(s_36_16), .cin(s_36_15), .o(t_286), .co(t_287), .cout(t_288));
compressor_4_2 u2_105(.a(s_37_2), .b(s_37_1), .c(s_37_0), .d(t_276), .cin(t_279), .o(t_289), .co(t_290), .cout(t_291));
compressor_4_2 u2_106(.a(s_37_5), .b(s_37_4), .c(s_37_3), .d(t_282), .cin(t_285), .o(t_292), .co(t_293), .cout(t_294));
compressor_4_2 u2_107(.a(s_37_9), .b(s_37_8), .c(s_37_7), .d(s_37_6), .cin(t_288), .o(t_295), .co(t_296), .cout(t_297));
compressor_4_2 u2_108(.a(s_37_14), .b(s_37_13), .c(s_37_12), .d(s_37_11), .cin(s_37_10), .o(t_298), .co(t_299), .cout(t_300));
compressor_3_2 u1_109(.a(s_37_17), .b(s_37_16), .cin(s_37_15), .o(t_301), .cout(t_302));
compressor_4_2 u2_110(.a(s_38_2), .b(s_38_1), .c(s_38_0), .d(t_291), .cin(t_294), .o(t_303), .co(t_304), .cout(t_305));
compressor_4_2 u2_111(.a(s_38_5), .b(s_38_4), .c(s_38_3), .d(t_297), .cin(t_300), .o(t_306), .co(t_307), .cout(t_308));
compressor_4_2 u2_112(.a(s_38_9), .b(s_38_8), .c(s_38_7), .d(s_38_6), .cin(t_302), .o(t_309), .co(t_310), .cout(t_311));
compressor_4_2 u2_113(.a(s_38_14), .b(s_38_13), .c(s_38_12), .d(s_38_11), .cin(s_38_10), .o(t_312), .co(t_313), .cout(t_314));
compressor_4_2 u2_114(.a(s_38_19), .b(s_38_18), .c(s_38_17), .d(s_38_16), .cin(s_38_15), .o(t_315), .co(t_316), .cout(t_317));
compressor_4_2 u2_115(.a(s_39_2), .b(s_39_1), .c(s_39_0), .d(t_305), .cin(t_308), .o(t_318), .co(t_319), .cout(t_320));
compressor_4_2 u2_116(.a(s_39_5), .b(s_39_4), .c(s_39_3), .d(t_311), .cin(t_314), .o(t_321), .co(t_322), .cout(t_323));
compressor_4_2 u2_117(.a(s_39_9), .b(s_39_8), .c(s_39_7), .d(s_39_6), .cin(t_317), .o(t_324), .co(t_325), .cout(t_326));
compressor_4_2 u2_118(.a(s_39_14), .b(s_39_13), .c(s_39_12), .d(s_39_11), .cin(s_39_10), .o(t_327), .co(t_328), .cout(t_329));
compressor_4_2 u2_119(.a(s_39_19), .b(s_39_18), .c(s_39_17), .d(s_39_16), .cin(s_39_15), .o(t_330), .co(t_331), .cout(t_332));
compressor_4_2 u2_120(.a(s_40_2), .b(s_40_1), .c(s_40_0), .d(t_320), .cin(t_323), .o(t_333), .co(t_334), .cout(t_335));
compressor_4_2 u2_121(.a(s_40_5), .b(s_40_4), .c(s_40_3), .d(t_326), .cin(t_329), .o(t_336), .co(t_337), .cout(t_338));
compressor_4_2 u2_122(.a(s_40_9), .b(s_40_8), .c(s_40_7), .d(s_40_6), .cin(t_332), .o(t_339), .co(t_340), .cout(t_341));
compressor_4_2 u2_123(.a(s_40_14), .b(s_40_13), .c(s_40_12), .d(s_40_11), .cin(s_40_10), .o(t_342), .co(t_343), .cout(t_344));
compressor_4_2 u2_124(.a(s_40_19), .b(s_40_18), .c(s_40_17), .d(s_40_16), .cin(s_40_15), .o(t_345), .co(t_346), .cout(t_347));
half_adder u0_125(.a(s_40_21), .b(s_40_20), .o(t_348), .cout(t_349));
compressor_4_2 u2_126(.a(s_41_2), .b(s_41_1), .c(s_41_0), .d(t_335), .cin(t_338), .o(t_350), .co(t_351), .cout(t_352));
compressor_4_2 u2_127(.a(s_41_5), .b(s_41_4), .c(s_41_3), .d(t_341), .cin(t_344), .o(t_353), .co(t_354), .cout(t_355));
compressor_4_2 u2_128(.a(s_41_8), .b(s_41_7), .c(s_41_6), .d(t_347), .cin(t_349), .o(t_356), .co(t_357), .cout(t_358));
compressor_4_2 u2_129(.a(s_41_13), .b(s_41_12), .c(s_41_11), .d(s_41_10), .cin(s_41_9), .o(t_359), .co(t_360), .cout(t_361));
compressor_4_2 u2_130(.a(s_41_18), .b(s_41_17), .c(s_41_16), .d(s_41_15), .cin(s_41_14), .o(t_362), .co(t_363), .cout(t_364));
half_adder u0_131(.a(s_41_20), .b(s_41_19), .o(t_365), .cout(t_366));
compressor_4_2 u2_132(.a(s_42_2), .b(s_42_1), .c(s_42_0), .d(t_352), .cin(t_355), .o(t_367), .co(t_368), .cout(t_369));
compressor_4_2 u2_133(.a(s_42_5), .b(s_42_4), .c(s_42_3), .d(t_358), .cin(t_361), .o(t_370), .co(t_371), .cout(t_372));
compressor_4_2 u2_134(.a(s_42_8), .b(s_42_7), .c(s_42_6), .d(t_364), .cin(t_366), .o(t_373), .co(t_374), .cout(t_375));
compressor_4_2 u2_135(.a(s_42_13), .b(s_42_12), .c(s_42_11), .d(s_42_10), .cin(s_42_9), .o(t_376), .co(t_377), .cout(t_378));
compressor_4_2 u2_136(.a(s_42_18), .b(s_42_17), .c(s_42_16), .d(s_42_15), .cin(s_42_14), .o(t_379), .co(t_380), .cout(t_381));
compressor_3_2 u1_137(.a(s_42_21), .b(s_42_20), .cin(s_42_19), .o(t_382), .cout(t_383));
compressor_4_2 u2_138(.a(s_43_2), .b(s_43_1), .c(s_43_0), .d(t_369), .cin(t_372), .o(t_384), .co(t_385), .cout(t_386));
compressor_4_2 u2_139(.a(s_43_5), .b(s_43_4), .c(s_43_3), .d(t_375), .cin(t_378), .o(t_387), .co(t_388), .cout(t_389));
compressor_4_2 u2_140(.a(s_43_8), .b(s_43_7), .c(s_43_6), .d(t_381), .cin(t_383), .o(t_390), .co(t_391), .cout(t_392));
compressor_4_2 u2_141(.a(s_43_13), .b(s_43_12), .c(s_43_11), .d(s_43_10), .cin(s_43_9), .o(t_393), .co(t_394), .cout(t_395));
compressor_4_2 u2_142(.a(s_43_18), .b(s_43_17), .c(s_43_16), .d(s_43_15), .cin(s_43_14), .o(t_396), .co(t_397), .cout(t_398));
compressor_3_2 u1_143(.a(s_43_21), .b(s_43_20), .cin(s_43_19), .o(t_399), .cout(t_400));
compressor_4_2 u2_144(.a(s_44_2), .b(s_44_1), .c(s_44_0), .d(t_386), .cin(t_389), .o(t_401), .co(t_402), .cout(t_403));
compressor_4_2 u2_145(.a(s_44_5), .b(s_44_4), .c(s_44_3), .d(t_392), .cin(t_395), .o(t_404), .co(t_405), .cout(t_406));
compressor_4_2 u2_146(.a(s_44_8), .b(s_44_7), .c(s_44_6), .d(t_398), .cin(t_400), .o(t_407), .co(t_408), .cout(t_409));
compressor_4_2 u2_147(.a(s_44_13), .b(s_44_12), .c(s_44_11), .d(s_44_10), .cin(s_44_9), .o(t_410), .co(t_411), .cout(t_412));
compressor_4_2 u2_148(.a(s_44_18), .b(s_44_17), .c(s_44_16), .d(s_44_15), .cin(s_44_14), .o(t_413), .co(t_414), .cout(t_415));
compressor_4_2 u2_149(.a(s_44_23), .b(s_44_22), .c(s_44_21), .d(s_44_20), .cin(s_44_19), .o(t_416), .co(t_417), .cout(t_418));
compressor_4_2 u2_150(.a(s_45_2), .b(s_45_1), .c(s_45_0), .d(t_403), .cin(t_406), .o(t_419), .co(t_420), .cout(t_421));
compressor_4_2 u2_151(.a(s_45_5), .b(s_45_4), .c(s_45_3), .d(t_409), .cin(t_412), .o(t_422), .co(t_423), .cout(t_424));
compressor_4_2 u2_152(.a(s_45_8), .b(s_45_7), .c(s_45_6), .d(t_415), .cin(t_418), .o(t_425), .co(t_426), .cout(t_427));
compressor_4_2 u2_153(.a(s_45_13), .b(s_45_12), .c(s_45_11), .d(s_45_10), .cin(s_45_9), .o(t_428), .co(t_429), .cout(t_430));
compressor_4_2 u2_154(.a(s_45_18), .b(s_45_17), .c(s_45_16), .d(s_45_15), .cin(s_45_14), .o(t_431), .co(t_432), .cout(t_433));
compressor_3_2 u1_155(.a(s_45_21), .b(s_45_20), .cin(s_45_19), .o(t_434), .cout(t_435));
compressor_4_2 u2_156(.a(s_46_2), .b(s_46_1), .c(s_46_0), .d(t_421), .cin(t_424), .o(t_436), .co(t_437), .cout(t_438));
compressor_4_2 u2_157(.a(s_46_5), .b(s_46_4), .c(s_46_3), .d(t_427), .cin(t_430), .o(t_439), .co(t_440), .cout(t_441));
compressor_4_2 u2_158(.a(s_46_8), .b(s_46_7), .c(s_46_6), .d(t_433), .cin(t_435), .o(t_442), .co(t_443), .cout(t_444));
compressor_4_2 u2_159(.a(s_46_13), .b(s_46_12), .c(s_46_11), .d(s_46_10), .cin(s_46_9), .o(t_445), .co(t_446), .cout(t_447));
compressor_4_2 u2_160(.a(s_46_18), .b(s_46_17), .c(s_46_16), .d(s_46_15), .cin(s_46_14), .o(t_448), .co(t_449), .cout(t_450));
compressor_4_2 u2_161(.a(s_46_23), .b(s_46_22), .c(s_46_21), .d(s_46_20), .cin(s_46_19), .o(t_451), .co(t_452), .cout(t_453));
compressor_4_2 u2_162(.a(s_47_2), .b(s_47_1), .c(s_47_0), .d(t_438), .cin(t_441), .o(t_454), .co(t_455), .cout(t_456));
compressor_4_2 u2_163(.a(s_47_5), .b(s_47_4), .c(s_47_3), .d(t_444), .cin(t_447), .o(t_457), .co(t_458), .cout(t_459));
compressor_4_2 u2_164(.a(s_47_8), .b(s_47_7), .c(s_47_6), .d(t_450), .cin(t_453), .o(t_460), .co(t_461), .cout(t_462));
compressor_4_2 u2_165(.a(s_47_13), .b(s_47_12), .c(s_47_11), .d(s_47_10), .cin(s_47_9), .o(t_463), .co(t_464), .cout(t_465));
compressor_4_2 u2_166(.a(s_47_18), .b(s_47_17), .c(s_47_16), .d(s_47_15), .cin(s_47_14), .o(t_466), .co(t_467), .cout(t_468));
compressor_4_2 u2_167(.a(s_47_23), .b(s_47_22), .c(s_47_21), .d(s_47_20), .cin(s_47_19), .o(t_469), .co(t_470), .cout(t_471));
compressor_4_2 u2_168(.a(s_48_2), .b(s_48_1), .c(s_48_0), .d(t_456), .cin(t_459), .o(t_472), .co(t_473), .cout(t_474));
compressor_4_2 u2_169(.a(s_48_5), .b(s_48_4), .c(s_48_3), .d(t_462), .cin(t_465), .o(t_475), .co(t_476), .cout(t_477));
compressor_4_2 u2_170(.a(s_48_8), .b(s_48_7), .c(s_48_6), .d(t_468), .cin(t_471), .o(t_478), .co(t_479), .cout(t_480));
compressor_4_2 u2_171(.a(s_48_13), .b(s_48_12), .c(s_48_11), .d(s_48_10), .cin(s_48_9), .o(t_481), .co(t_482), .cout(t_483));
compressor_4_2 u2_172(.a(s_48_18), .b(s_48_17), .c(s_48_16), .d(s_48_15), .cin(s_48_14), .o(t_484), .co(t_485), .cout(t_486));
compressor_4_2 u2_173(.a(s_48_23), .b(s_48_22), .c(s_48_21), .d(s_48_20), .cin(s_48_19), .o(t_487), .co(t_488), .cout(t_489));
half_adder u0_174(.a(s_48_25), .b(s_48_24), .o(t_490), .cout(t_491));
compressor_4_2 u2_175(.a(s_49_2), .b(s_49_1), .c(s_49_0), .d(t_474), .cin(t_477), .o(t_492), .co(t_493), .cout(t_494));
compressor_4_2 u2_176(.a(s_49_5), .b(s_49_4), .c(s_49_3), .d(t_480), .cin(t_483), .o(t_495), .co(t_496), .cout(t_497));
compressor_4_2 u2_177(.a(s_49_8), .b(s_49_7), .c(s_49_6), .d(t_486), .cin(t_489), .o(t_498), .co(t_499), .cout(t_500));
compressor_4_2 u2_178(.a(s_49_12), .b(s_49_11), .c(s_49_10), .d(s_49_9), .cin(t_491), .o(t_501), .co(t_502), .cout(t_503));
compressor_4_2 u2_179(.a(s_49_17), .b(s_49_16), .c(s_49_15), .d(s_49_14), .cin(s_49_13), .o(t_504), .co(t_505), .cout(t_506));
compressor_4_2 u2_180(.a(s_49_22), .b(s_49_21), .c(s_49_20), .d(s_49_19), .cin(s_49_18), .o(t_507), .co(t_508), .cout(t_509));
half_adder u0_181(.a(s_49_24), .b(s_49_23), .o(t_510), .cout(t_511));
compressor_4_2 u2_182(.a(s_50_2), .b(s_50_1), .c(s_50_0), .d(t_494), .cin(t_497), .o(t_512), .co(t_513), .cout(t_514));
compressor_4_2 u2_183(.a(s_50_5), .b(s_50_4), .c(s_50_3), .d(t_500), .cin(t_503), .o(t_515), .co(t_516), .cout(t_517));
compressor_4_2 u2_184(.a(s_50_8), .b(s_50_7), .c(s_50_6), .d(t_506), .cin(t_509), .o(t_518), .co(t_519), .cout(t_520));
compressor_4_2 u2_185(.a(s_50_12), .b(s_50_11), .c(s_50_10), .d(s_50_9), .cin(t_511), .o(t_521), .co(t_522), .cout(t_523));
compressor_4_2 u2_186(.a(s_50_17), .b(s_50_16), .c(s_50_15), .d(s_50_14), .cin(s_50_13), .o(t_524), .co(t_525), .cout(t_526));
compressor_4_2 u2_187(.a(s_50_22), .b(s_50_21), .c(s_50_20), .d(s_50_19), .cin(s_50_18), .o(t_527), .co(t_528), .cout(t_529));
compressor_3_2 u1_188(.a(s_50_25), .b(s_50_24), .cin(s_50_23), .o(t_530), .cout(t_531));
compressor_4_2 u2_189(.a(s_51_2), .b(s_51_1), .c(s_51_0), .d(t_514), .cin(t_517), .o(t_532), .co(t_533), .cout(t_534));
compressor_4_2 u2_190(.a(s_51_5), .b(s_51_4), .c(s_51_3), .d(t_520), .cin(t_523), .o(t_535), .co(t_536), .cout(t_537));
compressor_4_2 u2_191(.a(s_51_8), .b(s_51_7), .c(s_51_6), .d(t_526), .cin(t_529), .o(t_538), .co(t_539), .cout(t_540));
compressor_4_2 u2_192(.a(s_51_12), .b(s_51_11), .c(s_51_10), .d(s_51_9), .cin(t_531), .o(t_541), .co(t_542), .cout(t_543));
compressor_4_2 u2_193(.a(s_51_17), .b(s_51_16), .c(s_51_15), .d(s_51_14), .cin(s_51_13), .o(t_544), .co(t_545), .cout(t_546));
compressor_4_2 u2_194(.a(s_51_22), .b(s_51_21), .c(s_51_20), .d(s_51_19), .cin(s_51_18), .o(t_547), .co(t_548), .cout(t_549));
compressor_3_2 u1_195(.a(s_51_25), .b(s_51_24), .cin(s_51_23), .o(t_550), .cout(t_551));
compressor_4_2 u2_196(.a(s_52_2), .b(s_52_1), .c(s_52_0), .d(t_534), .cin(t_537), .o(t_552), .co(t_553), .cout(t_554));
compressor_4_2 u2_197(.a(s_52_5), .b(s_52_4), .c(s_52_3), .d(t_540), .cin(t_543), .o(t_555), .co(t_556), .cout(t_557));
compressor_4_2 u2_198(.a(s_52_8), .b(s_52_7), .c(s_52_6), .d(t_546), .cin(t_549), .o(t_558), .co(t_559), .cout(t_560));
compressor_4_2 u2_199(.a(s_52_12), .b(s_52_11), .c(s_52_10), .d(s_52_9), .cin(t_551), .o(t_561), .co(t_562), .cout(t_563));
compressor_4_2 u2_200(.a(s_52_17), .b(s_52_16), .c(s_52_15), .d(s_52_14), .cin(s_52_13), .o(t_564), .co(t_565), .cout(t_566));
compressor_4_2 u2_201(.a(s_52_22), .b(s_52_21), .c(s_52_20), .d(s_52_19), .cin(s_52_18), .o(t_567), .co(t_568), .cout(t_569));
compressor_4_2 u2_202(.a(s_52_27), .b(s_52_26), .c(s_52_25), .d(s_52_24), .cin(s_52_23), .o(t_570), .co(t_571), .cout(t_572));
compressor_4_2 u2_203(.a(s_53_2), .b(s_53_1), .c(s_53_0), .d(t_554), .cin(t_557), .o(t_573), .co(t_574), .cout(t_575));
compressor_4_2 u2_204(.a(s_53_5), .b(s_53_4), .c(s_53_3), .d(t_560), .cin(t_563), .o(t_576), .co(t_577), .cout(t_578));
compressor_4_2 u2_205(.a(s_53_8), .b(s_53_7), .c(s_53_6), .d(t_566), .cin(t_569), .o(t_579), .co(t_580), .cout(t_581));
compressor_4_2 u2_206(.a(s_53_12), .b(s_53_11), .c(s_53_10), .d(s_53_9), .cin(t_572), .o(t_582), .co(t_583), .cout(t_584));
compressor_4_2 u2_207(.a(s_53_17), .b(s_53_16), .c(s_53_15), .d(s_53_14), .cin(s_53_13), .o(t_585), .co(t_586), .cout(t_587));
compressor_4_2 u2_208(.a(s_53_22), .b(s_53_21), .c(s_53_20), .d(s_53_19), .cin(s_53_18), .o(t_588), .co(t_589), .cout(t_590));
compressor_3_2 u1_209(.a(s_53_25), .b(s_53_24), .cin(s_53_23), .o(t_591), .cout(t_592));
compressor_4_2 u2_210(.a(s_54_2), .b(s_54_1), .c(s_54_0), .d(t_575), .cin(t_578), .o(t_593), .co(t_594), .cout(t_595));
compressor_4_2 u2_211(.a(s_54_5), .b(s_54_4), .c(s_54_3), .d(t_581), .cin(t_584), .o(t_596), .co(t_597), .cout(t_598));
compressor_4_2 u2_212(.a(s_54_8), .b(s_54_7), .c(s_54_6), .d(t_587), .cin(t_590), .o(t_599), .co(t_600), .cout(t_601));
compressor_4_2 u2_213(.a(s_54_12), .b(s_54_11), .c(s_54_10), .d(s_54_9), .cin(t_592), .o(t_602), .co(t_603), .cout(t_604));
compressor_4_2 u2_214(.a(s_54_17), .b(s_54_16), .c(s_54_15), .d(s_54_14), .cin(s_54_13), .o(t_605), .co(t_606), .cout(t_607));
compressor_4_2 u2_215(.a(s_54_22), .b(s_54_21), .c(s_54_20), .d(s_54_19), .cin(s_54_18), .o(t_608), .co(t_609), .cout(t_610));
compressor_4_2 u2_216(.a(s_54_27), .b(s_54_26), .c(s_54_25), .d(s_54_24), .cin(s_54_23), .o(t_611), .co(t_612), .cout(t_613));
compressor_4_2 u2_217(.a(s_55_2), .b(s_55_1), .c(s_55_0), .d(t_595), .cin(t_598), .o(t_614), .co(t_615), .cout(t_616));
compressor_4_2 u2_218(.a(s_55_5), .b(s_55_4), .c(s_55_3), .d(t_601), .cin(t_604), .o(t_617), .co(t_618), .cout(t_619));
compressor_4_2 u2_219(.a(s_55_8), .b(s_55_7), .c(s_55_6), .d(t_607), .cin(t_610), .o(t_620), .co(t_621), .cout(t_622));
compressor_4_2 u2_220(.a(s_55_12), .b(s_55_11), .c(s_55_10), .d(s_55_9), .cin(t_613), .o(t_623), .co(t_624), .cout(t_625));
compressor_4_2 u2_221(.a(s_55_17), .b(s_55_16), .c(s_55_15), .d(s_55_14), .cin(s_55_13), .o(t_626), .co(t_627), .cout(t_628));
compressor_4_2 u2_222(.a(s_55_22), .b(s_55_21), .c(s_55_20), .d(s_55_19), .cin(s_55_18), .o(t_629), .co(t_630), .cout(t_631));
compressor_4_2 u2_223(.a(s_55_27), .b(s_55_26), .c(s_55_25), .d(s_55_24), .cin(s_55_23), .o(t_632), .co(t_633), .cout(t_634));
compressor_4_2 u2_224(.a(s_56_2), .b(s_56_1), .c(s_56_0), .d(t_616), .cin(t_619), .o(t_635), .co(t_636), .cout(t_637));
compressor_4_2 u2_225(.a(s_56_5), .b(s_56_4), .c(s_56_3), .d(t_622), .cin(t_625), .o(t_638), .co(t_639), .cout(t_640));
compressor_4_2 u2_226(.a(s_56_8), .b(s_56_7), .c(s_56_6), .d(t_628), .cin(t_631), .o(t_641), .co(t_642), .cout(t_643));
compressor_4_2 u2_227(.a(s_56_12), .b(s_56_11), .c(s_56_10), .d(s_56_9), .cin(t_634), .o(t_644), .co(t_645), .cout(t_646));
compressor_4_2 u2_228(.a(s_56_17), .b(s_56_16), .c(s_56_15), .d(s_56_14), .cin(s_56_13), .o(t_647), .co(t_648), .cout(t_649));
compressor_4_2 u2_229(.a(s_56_22), .b(s_56_21), .c(s_56_20), .d(s_56_19), .cin(s_56_18), .o(t_650), .co(t_651), .cout(t_652));
compressor_4_2 u2_230(.a(s_56_27), .b(s_56_26), .c(s_56_25), .d(s_56_24), .cin(s_56_23), .o(t_653), .co(t_654), .cout(t_655));
half_adder u0_231(.a(s_56_29), .b(s_56_28), .o(t_656), .cout(t_657));
compressor_4_2 u2_232(.a(s_57_2), .b(s_57_1), .c(s_57_0), .d(t_637), .cin(t_640), .o(t_658), .co(t_659), .cout(t_660));
compressor_4_2 u2_233(.a(s_57_5), .b(s_57_4), .c(s_57_3), .d(t_643), .cin(t_646), .o(t_661), .co(t_662), .cout(t_663));
compressor_4_2 u2_234(.a(s_57_8), .b(s_57_7), .c(s_57_6), .d(t_649), .cin(t_652), .o(t_664), .co(t_665), .cout(t_666));
compressor_4_2 u2_235(.a(s_57_11), .b(s_57_10), .c(s_57_9), .d(t_655), .cin(t_657), .o(t_667), .co(t_668), .cout(t_669));
compressor_4_2 u2_236(.a(s_57_16), .b(s_57_15), .c(s_57_14), .d(s_57_13), .cin(s_57_12), .o(t_670), .co(t_671), .cout(t_672));
compressor_4_2 u2_237(.a(s_57_21), .b(s_57_20), .c(s_57_19), .d(s_57_18), .cin(s_57_17), .o(t_673), .co(t_674), .cout(t_675));
compressor_4_2 u2_238(.a(s_57_26), .b(s_57_25), .c(s_57_24), .d(s_57_23), .cin(s_57_22), .o(t_676), .co(t_677), .cout(t_678));
half_adder u0_239(.a(s_57_28), .b(s_57_27), .o(t_679), .cout(t_680));
compressor_4_2 u2_240(.a(s_58_2), .b(s_58_1), .c(s_58_0), .d(t_660), .cin(t_663), .o(t_681), .co(t_682), .cout(t_683));
compressor_4_2 u2_241(.a(s_58_5), .b(s_58_4), .c(s_58_3), .d(t_666), .cin(t_669), .o(t_684), .co(t_685), .cout(t_686));
compressor_4_2 u2_242(.a(s_58_8), .b(s_58_7), .c(s_58_6), .d(t_672), .cin(t_675), .o(t_687), .co(t_688), .cout(t_689));
compressor_4_2 u2_243(.a(s_58_11), .b(s_58_10), .c(s_58_9), .d(t_678), .cin(t_680), .o(t_690), .co(t_691), .cout(t_692));
compressor_4_2 u2_244(.a(s_58_16), .b(s_58_15), .c(s_58_14), .d(s_58_13), .cin(s_58_12), .o(t_693), .co(t_694), .cout(t_695));
compressor_4_2 u2_245(.a(s_58_21), .b(s_58_20), .c(s_58_19), .d(s_58_18), .cin(s_58_17), .o(t_696), .co(t_697), .cout(t_698));
compressor_4_2 u2_246(.a(s_58_26), .b(s_58_25), .c(s_58_24), .d(s_58_23), .cin(s_58_22), .o(t_699), .co(t_700), .cout(t_701));
compressor_3_2 u1_247(.a(s_58_29), .b(s_58_28), .cin(s_58_27), .o(t_702), .cout(t_703));
compressor_4_2 u2_248(.a(s_59_2), .b(s_59_1), .c(s_59_0), .d(t_683), .cin(t_686), .o(t_704), .co(t_705), .cout(t_706));
compressor_4_2 u2_249(.a(s_59_5), .b(s_59_4), .c(s_59_3), .d(t_689), .cin(t_692), .o(t_707), .co(t_708), .cout(t_709));
compressor_4_2 u2_250(.a(s_59_8), .b(s_59_7), .c(s_59_6), .d(t_695), .cin(t_698), .o(t_710), .co(t_711), .cout(t_712));
compressor_4_2 u2_251(.a(s_59_11), .b(s_59_10), .c(s_59_9), .d(t_701), .cin(t_703), .o(t_713), .co(t_714), .cout(t_715));
compressor_4_2 u2_252(.a(s_59_16), .b(s_59_15), .c(s_59_14), .d(s_59_13), .cin(s_59_12), .o(t_716), .co(t_717), .cout(t_718));
compressor_4_2 u2_253(.a(s_59_21), .b(s_59_20), .c(s_59_19), .d(s_59_18), .cin(s_59_17), .o(t_719), .co(t_720), .cout(t_721));
compressor_4_2 u2_254(.a(s_59_26), .b(s_59_25), .c(s_59_24), .d(s_59_23), .cin(s_59_22), .o(t_722), .co(t_723), .cout(t_724));
compressor_3_2 u1_255(.a(s_59_29), .b(s_59_28), .cin(s_59_27), .o(t_725), .cout(t_726));
compressor_4_2 u2_256(.a(s_60_2), .b(s_60_1), .c(s_60_0), .d(t_706), .cin(t_709), .o(t_727), .co(t_728), .cout(t_729));
compressor_4_2 u2_257(.a(s_60_5), .b(s_60_4), .c(s_60_3), .d(t_712), .cin(t_715), .o(t_730), .co(t_731), .cout(t_732));
compressor_4_2 u2_258(.a(s_60_8), .b(s_60_7), .c(s_60_6), .d(t_718), .cin(t_721), .o(t_733), .co(t_734), .cout(t_735));
compressor_4_2 u2_259(.a(s_60_11), .b(s_60_10), .c(s_60_9), .d(t_724), .cin(t_726), .o(t_736), .co(t_737), .cout(t_738));
compressor_4_2 u2_260(.a(s_60_16), .b(s_60_15), .c(s_60_14), .d(s_60_13), .cin(s_60_12), .o(t_739), .co(t_740), .cout(t_741));
compressor_4_2 u2_261(.a(s_60_21), .b(s_60_20), .c(s_60_19), .d(s_60_18), .cin(s_60_17), .o(t_742), .co(t_743), .cout(t_744));
compressor_4_2 u2_262(.a(s_60_26), .b(s_60_25), .c(s_60_24), .d(s_60_23), .cin(s_60_22), .o(t_745), .co(t_746), .cout(t_747));
compressor_4_2 u2_263(.a(s_60_31), .b(s_60_30), .c(s_60_29), .d(s_60_28), .cin(s_60_27), .o(t_748), .co(t_749), .cout(t_750));
compressor_4_2 u2_264(.a(s_61_2), .b(s_61_1), .c(s_61_0), .d(t_729), .cin(t_732), .o(t_751), .co(t_752), .cout(t_753));
compressor_4_2 u2_265(.a(s_61_5), .b(s_61_4), .c(s_61_3), .d(t_735), .cin(t_738), .o(t_754), .co(t_755), .cout(t_756));
compressor_4_2 u2_266(.a(s_61_8), .b(s_61_7), .c(s_61_6), .d(t_741), .cin(t_744), .o(t_757), .co(t_758), .cout(t_759));
compressor_4_2 u2_267(.a(s_61_11), .b(s_61_10), .c(s_61_9), .d(t_747), .cin(t_750), .o(t_760), .co(t_761), .cout(t_762));
compressor_4_2 u2_268(.a(s_61_16), .b(s_61_15), .c(s_61_14), .d(s_61_13), .cin(s_61_12), .o(t_763), .co(t_764), .cout(t_765));
compressor_4_2 u2_269(.a(s_61_21), .b(s_61_20), .c(s_61_19), .d(s_61_18), .cin(s_61_17), .o(t_766), .co(t_767), .cout(t_768));
compressor_4_2 u2_270(.a(s_61_26), .b(s_61_25), .c(s_61_24), .d(s_61_23), .cin(s_61_22), .o(t_769), .co(t_770), .cout(t_771));
compressor_3_2 u1_271(.a(s_61_29), .b(s_61_28), .cin(s_61_27), .o(t_772), .cout(t_773));
compressor_4_2 u2_272(.a(s_62_2), .b(s_62_1), .c(s_62_0), .d(t_753), .cin(t_756), .o(t_774), .co(t_775), .cout(t_776));
compressor_4_2 u2_273(.a(s_62_5), .b(s_62_4), .c(s_62_3), .d(t_759), .cin(t_762), .o(t_777), .co(t_778), .cout(t_779));
compressor_4_2 u2_274(.a(s_62_8), .b(s_62_7), .c(s_62_6), .d(t_765), .cin(t_768), .o(t_780), .co(t_781), .cout(t_782));
compressor_4_2 u2_275(.a(s_62_11), .b(s_62_10), .c(s_62_9), .d(t_771), .cin(t_773), .o(t_783), .co(t_784), .cout(t_785));
compressor_4_2 u2_276(.a(s_62_16), .b(s_62_15), .c(s_62_14), .d(s_62_13), .cin(s_62_12), .o(t_786), .co(t_787), .cout(t_788));
compressor_4_2 u2_277(.a(s_62_21), .b(s_62_20), .c(s_62_19), .d(s_62_18), .cin(s_62_17), .o(t_789), .co(t_790), .cout(t_791));
compressor_4_2 u2_278(.a(s_62_26), .b(s_62_25), .c(s_62_24), .d(s_62_23), .cin(s_62_22), .o(t_792), .co(t_793), .cout(t_794));
compressor_4_2 u2_279(.a(s_62_31), .b(s_62_30), .c(s_62_29), .d(s_62_28), .cin(s_62_27), .o(t_795), .co(t_796), .cout(t_797));
compressor_4_2 u2_280(.a(s_63_2), .b(s_63_1), .c(s_63_0), .d(t_776), .cin(t_779), .o(t_798), .co(t_799), .cout(t_800));
compressor_4_2 u2_281(.a(s_63_5), .b(s_63_4), .c(s_63_3), .d(t_782), .cin(t_785), .o(t_801), .co(t_802), .cout(t_803));
compressor_4_2 u2_282(.a(s_63_8), .b(s_63_7), .c(s_63_6), .d(t_788), .cin(t_791), .o(t_804), .co(t_805), .cout(t_806));
compressor_4_2 u2_283(.a(s_63_11), .b(s_63_10), .c(s_63_9), .d(t_794), .cin(t_797), .o(t_807), .co(t_808), .cout(t_809));
compressor_4_2 u2_284(.a(s_63_16), .b(s_63_15), .c(s_63_14), .d(s_63_13), .cin(s_63_12), .o(t_810), .co(t_811), .cout(t_812));
compressor_4_2 u2_285(.a(s_63_21), .b(s_63_20), .c(s_63_19), .d(s_63_18), .cin(s_63_17), .o(t_813), .co(t_814), .cout(t_815));
compressor_4_2 u2_286(.a(s_63_26), .b(s_63_25), .c(s_63_24), .d(s_63_23), .cin(s_63_22), .o(t_816), .co(t_817), .cout(t_818));
compressor_4_2 u2_287(.a(s_63_31), .b(s_63_30), .c(s_63_29), .d(s_63_28), .cin(s_63_27), .o(t_819), .co(t_820), .cout(t_821));
compressor_4_2 u2_288(.a(s_64_2), .b(s_64_1), .c(s_64_0), .d(t_800), .cin(t_803), .o(t_822), .co(t_823), .cout(t_824));
compressor_4_2 u2_289(.a(s_64_5), .b(s_64_4), .c(s_64_3), .d(t_806), .cin(t_809), .o(t_825), .co(t_826), .cout(t_827));
compressor_4_2 u2_290(.a(s_64_8), .b(s_64_7), .c(s_64_6), .d(t_812), .cin(t_815), .o(t_828), .co(t_829), .cout(t_830));
compressor_4_2 u2_291(.a(s_64_11), .b(s_64_10), .c(s_64_9), .d(t_818), .cin(t_821), .o(t_831), .co(t_832), .cout(t_833));
compressor_4_2 u2_292(.a(s_64_16), .b(s_64_15), .c(s_64_14), .d(s_64_13), .cin(s_64_12), .o(t_834), .co(t_835), .cout(t_836));
compressor_4_2 u2_293(.a(s_64_21), .b(s_64_20), .c(s_64_19), .d(s_64_18), .cin(s_64_17), .o(t_837), .co(t_838), .cout(t_839));
compressor_4_2 u2_294(.a(s_64_26), .b(s_64_25), .c(s_64_24), .d(s_64_23), .cin(s_64_22), .o(t_840), .co(t_841), .cout(t_842));
compressor_4_2 u2_295(.a(s_64_31), .b(s_64_30), .c(s_64_29), .d(s_64_28), .cin(s_64_27), .o(t_843), .co(t_844), .cout(t_845));
half_adder u0_296(.a(s_64_33), .b(s_64_32), .o(t_846), .cout(t_847));
compressor_4_2 u2_297(.a(s_65_2), .b(s_65_1), .c(s_65_0), .d(t_824), .cin(t_827), .o(t_848), .co(t_849), .cout(t_850));
compressor_4_2 u2_298(.a(s_65_5), .b(s_65_4), .c(s_65_3), .d(t_830), .cin(t_833), .o(t_851), .co(t_852), .cout(t_853));
compressor_4_2 u2_299(.a(s_65_8), .b(s_65_7), .c(s_65_6), .d(t_836), .cin(t_839), .o(t_854), .co(t_855), .cout(t_856));
compressor_4_2 u2_300(.a(s_65_11), .b(s_65_10), .c(s_65_9), .d(t_842), .cin(t_845), .o(t_857), .co(t_858), .cout(t_859));
compressor_4_2 u2_301(.a(s_65_15), .b(s_65_14), .c(s_65_13), .d(s_65_12), .cin(t_847), .o(t_860), .co(t_861), .cout(t_862));
compressor_4_2 u2_302(.a(s_65_20), .b(s_65_19), .c(s_65_18), .d(s_65_17), .cin(s_65_16), .o(t_863), .co(t_864), .cout(t_865));
compressor_4_2 u2_303(.a(s_65_25), .b(s_65_24), .c(s_65_23), .d(s_65_22), .cin(s_65_21), .o(t_866), .co(t_867), .cout(t_868));
compressor_4_2 u2_304(.a(s_65_30), .b(s_65_29), .c(s_65_28), .d(s_65_27), .cin(s_65_26), .o(t_869), .co(t_870), .cout(t_871));
half_adder u0_305(.a(s_65_32), .b(s_65_31), .o(t_872), .cout(t_873));
compressor_4_2 u2_306(.a(s_66_2), .b(s_66_1), .c(s_66_0), .d(t_850), .cin(t_853), .o(t_874), .co(t_875), .cout(t_876));
compressor_4_2 u2_307(.a(s_66_5), .b(s_66_4), .c(s_66_3), .d(t_856), .cin(t_859), .o(t_877), .co(t_878), .cout(t_879));
compressor_4_2 u2_308(.a(s_66_8), .b(s_66_7), .c(s_66_6), .d(t_862), .cin(t_865), .o(t_880), .co(t_881), .cout(t_882));
compressor_4_2 u2_309(.a(s_66_11), .b(s_66_10), .c(s_66_9), .d(t_868), .cin(t_871), .o(t_883), .co(t_884), .cout(t_885));
compressor_4_2 u2_310(.a(s_66_15), .b(s_66_14), .c(s_66_13), .d(s_66_12), .cin(t_873), .o(t_886), .co(t_887), .cout(t_888));
compressor_4_2 u2_311(.a(s_66_20), .b(s_66_19), .c(s_66_18), .d(s_66_17), .cin(s_66_16), .o(t_889), .co(t_890), .cout(t_891));
compressor_4_2 u2_312(.a(s_66_25), .b(s_66_24), .c(s_66_23), .d(s_66_22), .cin(s_66_21), .o(t_892), .co(t_893), .cout(t_894));
compressor_4_2 u2_313(.a(s_66_30), .b(s_66_29), .c(s_66_28), .d(s_66_27), .cin(s_66_26), .o(t_895), .co(t_896), .cout(t_897));
compressor_3_2 u1_314(.a(s_66_33), .b(s_66_32), .cin(s_66_31), .o(t_898), .cout(t_899));
compressor_4_2 u2_315(.a(s_67_2), .b(s_67_1), .c(s_67_0), .d(t_876), .cin(t_879), .o(t_900), .co(t_901), .cout(t_902));
compressor_4_2 u2_316(.a(s_67_5), .b(s_67_4), .c(s_67_3), .d(t_882), .cin(t_885), .o(t_903), .co(t_904), .cout(t_905));
compressor_4_2 u2_317(.a(s_67_8), .b(s_67_7), .c(s_67_6), .d(t_888), .cin(t_891), .o(t_906), .co(t_907), .cout(t_908));
compressor_4_2 u2_318(.a(s_67_11), .b(s_67_10), .c(s_67_9), .d(t_894), .cin(t_897), .o(t_909), .co(t_910), .cout(t_911));
compressor_4_2 u2_319(.a(s_67_15), .b(s_67_14), .c(s_67_13), .d(s_67_12), .cin(t_899), .o(t_912), .co(t_913), .cout(t_914));
compressor_4_2 u2_320(.a(s_67_20), .b(s_67_19), .c(s_67_18), .d(s_67_17), .cin(s_67_16), .o(t_915), .co(t_916), .cout(t_917));
compressor_4_2 u2_321(.a(s_67_25), .b(s_67_24), .c(s_67_23), .d(s_67_22), .cin(s_67_21), .o(t_918), .co(t_919), .cout(t_920));
compressor_4_2 u2_322(.a(s_67_30), .b(s_67_29), .c(s_67_28), .d(s_67_27), .cin(s_67_26), .o(t_921), .co(t_922), .cout(t_923));
compressor_3_2 u1_323(.a(s_67_33), .b(s_67_32), .cin(s_67_31), .o(t_924), .cout(t_925));
compressor_4_2 u2_324(.a(s_68_2), .b(s_68_1), .c(s_68_0), .d(t_902), .cin(t_905), .o(t_926), .co(t_927), .cout(t_928));
compressor_4_2 u2_325(.a(s_68_5), .b(s_68_4), .c(s_68_3), .d(t_908), .cin(t_911), .o(t_929), .co(t_930), .cout(t_931));
compressor_4_2 u2_326(.a(s_68_8), .b(s_68_7), .c(s_68_6), .d(t_914), .cin(t_917), .o(t_932), .co(t_933), .cout(t_934));
compressor_4_2 u2_327(.a(s_68_11), .b(s_68_10), .c(s_68_9), .d(t_920), .cin(t_923), .o(t_935), .co(t_936), .cout(t_937));
compressor_4_2 u2_328(.a(s_68_15), .b(s_68_14), .c(s_68_13), .d(s_68_12), .cin(t_925), .o(t_938), .co(t_939), .cout(t_940));
compressor_4_2 u2_329(.a(s_68_20), .b(s_68_19), .c(s_68_18), .d(s_68_17), .cin(s_68_16), .o(t_941), .co(t_942), .cout(t_943));
compressor_4_2 u2_330(.a(s_68_25), .b(s_68_24), .c(s_68_23), .d(s_68_22), .cin(s_68_21), .o(t_944), .co(t_945), .cout(t_946));
compressor_4_2 u2_331(.a(s_68_30), .b(s_68_29), .c(s_68_28), .d(s_68_27), .cin(s_68_26), .o(t_947), .co(t_948), .cout(t_949));
compressor_4_2 u2_332(.a(s_68_35), .b(s_68_34), .c(s_68_33), .d(s_68_32), .cin(s_68_31), .o(t_950), .co(t_951), .cout(t_952));
compressor_4_2 u2_333(.a(s_69_2), .b(s_69_1), .c(s_69_0), .d(t_928), .cin(t_931), .o(t_953), .co(t_954), .cout(t_955));
compressor_4_2 u2_334(.a(s_69_5), .b(s_69_4), .c(s_69_3), .d(t_934), .cin(t_937), .o(t_956), .co(t_957), .cout(t_958));
compressor_4_2 u2_335(.a(s_69_8), .b(s_69_7), .c(s_69_6), .d(t_940), .cin(t_943), .o(t_959), .co(t_960), .cout(t_961));
compressor_4_2 u2_336(.a(s_69_11), .b(s_69_10), .c(s_69_9), .d(t_946), .cin(t_949), .o(t_962), .co(t_963), .cout(t_964));
compressor_4_2 u2_337(.a(s_69_15), .b(s_69_14), .c(s_69_13), .d(s_69_12), .cin(t_952), .o(t_965), .co(t_966), .cout(t_967));
compressor_4_2 u2_338(.a(s_69_20), .b(s_69_19), .c(s_69_18), .d(s_69_17), .cin(s_69_16), .o(t_968), .co(t_969), .cout(t_970));
compressor_4_2 u2_339(.a(s_69_25), .b(s_69_24), .c(s_69_23), .d(s_69_22), .cin(s_69_21), .o(t_971), .co(t_972), .cout(t_973));
compressor_4_2 u2_340(.a(s_69_30), .b(s_69_29), .c(s_69_28), .d(s_69_27), .cin(s_69_26), .o(t_974), .co(t_975), .cout(t_976));
compressor_3_2 u1_341(.a(s_69_33), .b(s_69_32), .cin(s_69_31), .o(t_977), .cout(t_978));
compressor_4_2 u2_342(.a(s_70_2), .b(s_70_1), .c(s_70_0), .d(t_955), .cin(t_958), .o(t_979), .co(t_980), .cout(t_981));
compressor_4_2 u2_343(.a(s_70_5), .b(s_70_4), .c(s_70_3), .d(t_961), .cin(t_964), .o(t_982), .co(t_983), .cout(t_984));
compressor_4_2 u2_344(.a(s_70_8), .b(s_70_7), .c(s_70_6), .d(t_967), .cin(t_970), .o(t_985), .co(t_986), .cout(t_987));
compressor_4_2 u2_345(.a(s_70_11), .b(s_70_10), .c(s_70_9), .d(t_973), .cin(t_976), .o(t_988), .co(t_989), .cout(t_990));
compressor_4_2 u2_346(.a(s_70_15), .b(s_70_14), .c(s_70_13), .d(s_70_12), .cin(t_978), .o(t_991), .co(t_992), .cout(t_993));
compressor_4_2 u2_347(.a(s_70_20), .b(s_70_19), .c(s_70_18), .d(s_70_17), .cin(s_70_16), .o(t_994), .co(t_995), .cout(t_996));
compressor_4_2 u2_348(.a(s_70_25), .b(s_70_24), .c(s_70_23), .d(s_70_22), .cin(s_70_21), .o(t_997), .co(t_998), .cout(t_999));
compressor_4_2 u2_349(.a(s_70_30), .b(s_70_29), .c(s_70_28), .d(s_70_27), .cin(s_70_26), .o(t_1000), .co(t_1001), .cout(t_1002));
compressor_4_2 u2_350(.a(s_70_35), .b(s_70_34), .c(s_70_33), .d(s_70_32), .cin(s_70_31), .o(t_1003), .co(t_1004), .cout(t_1005));
compressor_4_2 u2_351(.a(s_71_2), .b(s_71_1), .c(s_71_0), .d(t_981), .cin(t_984), .o(t_1006), .co(t_1007), .cout(t_1008));
compressor_4_2 u2_352(.a(s_71_5), .b(s_71_4), .c(s_71_3), .d(t_987), .cin(t_990), .o(t_1009), .co(t_1010), .cout(t_1011));
compressor_4_2 u2_353(.a(s_71_8), .b(s_71_7), .c(s_71_6), .d(t_993), .cin(t_996), .o(t_1012), .co(t_1013), .cout(t_1014));
compressor_4_2 u2_354(.a(s_71_11), .b(s_71_10), .c(s_71_9), .d(t_999), .cin(t_1002), .o(t_1015), .co(t_1016), .cout(t_1017));
compressor_4_2 u2_355(.a(s_71_15), .b(s_71_14), .c(s_71_13), .d(s_71_12), .cin(t_1005), .o(t_1018), .co(t_1019), .cout(t_1020));
compressor_4_2 u2_356(.a(s_71_20), .b(s_71_19), .c(s_71_18), .d(s_71_17), .cin(s_71_16), .o(t_1021), .co(t_1022), .cout(t_1023));
compressor_4_2 u2_357(.a(s_71_25), .b(s_71_24), .c(s_71_23), .d(s_71_22), .cin(s_71_21), .o(t_1024), .co(t_1025), .cout(t_1026));
compressor_4_2 u2_358(.a(s_71_30), .b(s_71_29), .c(s_71_28), .d(s_71_27), .cin(s_71_26), .o(t_1027), .co(t_1028), .cout(t_1029));
compressor_4_2 u2_359(.a(s_71_35), .b(s_71_34), .c(s_71_33), .d(s_71_32), .cin(s_71_31), .o(t_1030), .co(t_1031), .cout(t_1032));
compressor_4_2 u2_360(.a(s_72_2), .b(s_72_1), .c(s_72_0), .d(t_1008), .cin(t_1011), .o(t_1033), .co(t_1034), .cout(t_1035));
compressor_4_2 u2_361(.a(s_72_5), .b(s_72_4), .c(s_72_3), .d(t_1014), .cin(t_1017), .o(t_1036), .co(t_1037), .cout(t_1038));
compressor_4_2 u2_362(.a(s_72_8), .b(s_72_7), .c(s_72_6), .d(t_1020), .cin(t_1023), .o(t_1039), .co(t_1040), .cout(t_1041));
compressor_4_2 u2_363(.a(s_72_11), .b(s_72_10), .c(s_72_9), .d(t_1026), .cin(t_1029), .o(t_1042), .co(t_1043), .cout(t_1044));
compressor_4_2 u2_364(.a(s_72_15), .b(s_72_14), .c(s_72_13), .d(s_72_12), .cin(t_1032), .o(t_1045), .co(t_1046), .cout(t_1047));
compressor_4_2 u2_365(.a(s_72_20), .b(s_72_19), .c(s_72_18), .d(s_72_17), .cin(s_72_16), .o(t_1048), .co(t_1049), .cout(t_1050));
compressor_4_2 u2_366(.a(s_72_25), .b(s_72_24), .c(s_72_23), .d(s_72_22), .cin(s_72_21), .o(t_1051), .co(t_1052), .cout(t_1053));
compressor_4_2 u2_367(.a(s_72_30), .b(s_72_29), .c(s_72_28), .d(s_72_27), .cin(s_72_26), .o(t_1054), .co(t_1055), .cout(t_1056));
compressor_4_2 u2_368(.a(s_72_35), .b(s_72_34), .c(s_72_33), .d(s_72_32), .cin(s_72_31), .o(t_1057), .co(t_1058), .cout(t_1059));
half_adder u0_369(.a(s_72_37), .b(s_72_36), .o(t_1060), .cout(t_1061));
compressor_4_2 u2_370(.a(s_73_2), .b(s_73_1), .c(s_73_0), .d(t_1035), .cin(t_1038), .o(t_1062), .co(t_1063), .cout(t_1064));
compressor_4_2 u2_371(.a(s_73_5), .b(s_73_4), .c(s_73_3), .d(t_1041), .cin(t_1044), .o(t_1065), .co(t_1066), .cout(t_1067));
compressor_4_2 u2_372(.a(s_73_8), .b(s_73_7), .c(s_73_6), .d(t_1047), .cin(t_1050), .o(t_1068), .co(t_1069), .cout(t_1070));
compressor_4_2 u2_373(.a(s_73_11), .b(s_73_10), .c(s_73_9), .d(t_1053), .cin(t_1056), .o(t_1071), .co(t_1072), .cout(t_1073));
compressor_4_2 u2_374(.a(s_73_14), .b(s_73_13), .c(s_73_12), .d(t_1059), .cin(t_1061), .o(t_1074), .co(t_1075), .cout(t_1076));
compressor_4_2 u2_375(.a(s_73_19), .b(s_73_18), .c(s_73_17), .d(s_73_16), .cin(s_73_15), .o(t_1077), .co(t_1078), .cout(t_1079));
compressor_4_2 u2_376(.a(s_73_24), .b(s_73_23), .c(s_73_22), .d(s_73_21), .cin(s_73_20), .o(t_1080), .co(t_1081), .cout(t_1082));
compressor_4_2 u2_377(.a(s_73_29), .b(s_73_28), .c(s_73_27), .d(s_73_26), .cin(s_73_25), .o(t_1083), .co(t_1084), .cout(t_1085));
compressor_4_2 u2_378(.a(s_73_34), .b(s_73_33), .c(s_73_32), .d(s_73_31), .cin(s_73_30), .o(t_1086), .co(t_1087), .cout(t_1088));
half_adder u0_379(.a(s_73_36), .b(s_73_35), .o(t_1089), .cout(t_1090));
compressor_4_2 u2_380(.a(s_74_2), .b(s_74_1), .c(s_74_0), .d(t_1064), .cin(t_1067), .o(t_1091), .co(t_1092), .cout(t_1093));
compressor_4_2 u2_381(.a(s_74_5), .b(s_74_4), .c(s_74_3), .d(t_1070), .cin(t_1073), .o(t_1094), .co(t_1095), .cout(t_1096));
compressor_4_2 u2_382(.a(s_74_8), .b(s_74_7), .c(s_74_6), .d(t_1076), .cin(t_1079), .o(t_1097), .co(t_1098), .cout(t_1099));
compressor_4_2 u2_383(.a(s_74_11), .b(s_74_10), .c(s_74_9), .d(t_1082), .cin(t_1085), .o(t_1100), .co(t_1101), .cout(t_1102));
compressor_4_2 u2_384(.a(s_74_14), .b(s_74_13), .c(s_74_12), .d(t_1088), .cin(t_1090), .o(t_1103), .co(t_1104), .cout(t_1105));
compressor_4_2 u2_385(.a(s_74_19), .b(s_74_18), .c(s_74_17), .d(s_74_16), .cin(s_74_15), .o(t_1106), .co(t_1107), .cout(t_1108));
compressor_4_2 u2_386(.a(s_74_24), .b(s_74_23), .c(s_74_22), .d(s_74_21), .cin(s_74_20), .o(t_1109), .co(t_1110), .cout(t_1111));
compressor_4_2 u2_387(.a(s_74_29), .b(s_74_28), .c(s_74_27), .d(s_74_26), .cin(s_74_25), .o(t_1112), .co(t_1113), .cout(t_1114));
compressor_4_2 u2_388(.a(s_74_34), .b(s_74_33), .c(s_74_32), .d(s_74_31), .cin(s_74_30), .o(t_1115), .co(t_1116), .cout(t_1117));
compressor_3_2 u1_389(.a(s_74_37), .b(s_74_36), .cin(s_74_35), .o(t_1118), .cout(t_1119));
compressor_4_2 u2_390(.a(s_75_2), .b(s_75_1), .c(s_75_0), .d(t_1093), .cin(t_1096), .o(t_1120), .co(t_1121), .cout(t_1122));
compressor_4_2 u2_391(.a(s_75_5), .b(s_75_4), .c(s_75_3), .d(t_1099), .cin(t_1102), .o(t_1123), .co(t_1124), .cout(t_1125));
compressor_4_2 u2_392(.a(s_75_8), .b(s_75_7), .c(s_75_6), .d(t_1105), .cin(t_1108), .o(t_1126), .co(t_1127), .cout(t_1128));
compressor_4_2 u2_393(.a(s_75_11), .b(s_75_10), .c(s_75_9), .d(t_1111), .cin(t_1114), .o(t_1129), .co(t_1130), .cout(t_1131));
compressor_4_2 u2_394(.a(s_75_14), .b(s_75_13), .c(s_75_12), .d(t_1117), .cin(t_1119), .o(t_1132), .co(t_1133), .cout(t_1134));
compressor_4_2 u2_395(.a(s_75_19), .b(s_75_18), .c(s_75_17), .d(s_75_16), .cin(s_75_15), .o(t_1135), .co(t_1136), .cout(t_1137));
compressor_4_2 u2_396(.a(s_75_24), .b(s_75_23), .c(s_75_22), .d(s_75_21), .cin(s_75_20), .o(t_1138), .co(t_1139), .cout(t_1140));
compressor_4_2 u2_397(.a(s_75_29), .b(s_75_28), .c(s_75_27), .d(s_75_26), .cin(s_75_25), .o(t_1141), .co(t_1142), .cout(t_1143));
compressor_4_2 u2_398(.a(s_75_34), .b(s_75_33), .c(s_75_32), .d(s_75_31), .cin(s_75_30), .o(t_1144), .co(t_1145), .cout(t_1146));
compressor_3_2 u1_399(.a(s_75_37), .b(s_75_36), .cin(s_75_35), .o(t_1147), .cout(t_1148));
compressor_4_2 u2_400(.a(s_76_2), .b(s_76_1), .c(s_76_0), .d(t_1122), .cin(t_1125), .o(t_1149), .co(t_1150), .cout(t_1151));
compressor_4_2 u2_401(.a(s_76_5), .b(s_76_4), .c(s_76_3), .d(t_1128), .cin(t_1131), .o(t_1152), .co(t_1153), .cout(t_1154));
compressor_4_2 u2_402(.a(s_76_8), .b(s_76_7), .c(s_76_6), .d(t_1134), .cin(t_1137), .o(t_1155), .co(t_1156), .cout(t_1157));
compressor_4_2 u2_403(.a(s_76_11), .b(s_76_10), .c(s_76_9), .d(t_1140), .cin(t_1143), .o(t_1158), .co(t_1159), .cout(t_1160));
compressor_4_2 u2_404(.a(s_76_14), .b(s_76_13), .c(s_76_12), .d(t_1146), .cin(t_1148), .o(t_1161), .co(t_1162), .cout(t_1163));
compressor_4_2 u2_405(.a(s_76_19), .b(s_76_18), .c(s_76_17), .d(s_76_16), .cin(s_76_15), .o(t_1164), .co(t_1165), .cout(t_1166));
compressor_4_2 u2_406(.a(s_76_24), .b(s_76_23), .c(s_76_22), .d(s_76_21), .cin(s_76_20), .o(t_1167), .co(t_1168), .cout(t_1169));
compressor_4_2 u2_407(.a(s_76_29), .b(s_76_28), .c(s_76_27), .d(s_76_26), .cin(s_76_25), .o(t_1170), .co(t_1171), .cout(t_1172));
compressor_4_2 u2_408(.a(s_76_34), .b(s_76_33), .c(s_76_32), .d(s_76_31), .cin(s_76_30), .o(t_1173), .co(t_1174), .cout(t_1175));
compressor_4_2 u2_409(.a(s_76_39), .b(s_76_38), .c(s_76_37), .d(s_76_36), .cin(s_76_35), .o(t_1176), .co(t_1177), .cout(t_1178));
compressor_4_2 u2_410(.a(s_77_2), .b(s_77_1), .c(s_77_0), .d(t_1151), .cin(t_1154), .o(t_1179), .co(t_1180), .cout(t_1181));
compressor_4_2 u2_411(.a(s_77_5), .b(s_77_4), .c(s_77_3), .d(t_1157), .cin(t_1160), .o(t_1182), .co(t_1183), .cout(t_1184));
compressor_4_2 u2_412(.a(s_77_8), .b(s_77_7), .c(s_77_6), .d(t_1163), .cin(t_1166), .o(t_1185), .co(t_1186), .cout(t_1187));
compressor_4_2 u2_413(.a(s_77_11), .b(s_77_10), .c(s_77_9), .d(t_1169), .cin(t_1172), .o(t_1188), .co(t_1189), .cout(t_1190));
compressor_4_2 u2_414(.a(s_77_14), .b(s_77_13), .c(s_77_12), .d(t_1175), .cin(t_1178), .o(t_1191), .co(t_1192), .cout(t_1193));
compressor_4_2 u2_415(.a(s_77_19), .b(s_77_18), .c(s_77_17), .d(s_77_16), .cin(s_77_15), .o(t_1194), .co(t_1195), .cout(t_1196));
compressor_4_2 u2_416(.a(s_77_24), .b(s_77_23), .c(s_77_22), .d(s_77_21), .cin(s_77_20), .o(t_1197), .co(t_1198), .cout(t_1199));
compressor_4_2 u2_417(.a(s_77_29), .b(s_77_28), .c(s_77_27), .d(s_77_26), .cin(s_77_25), .o(t_1200), .co(t_1201), .cout(t_1202));
compressor_4_2 u2_418(.a(s_77_34), .b(s_77_33), .c(s_77_32), .d(s_77_31), .cin(s_77_30), .o(t_1203), .co(t_1204), .cout(t_1205));
compressor_3_2 u1_419(.a(s_77_37), .b(s_77_36), .cin(s_77_35), .o(t_1206), .cout(t_1207));
compressor_4_2 u2_420(.a(s_78_2), .b(s_78_1), .c(s_78_0), .d(t_1181), .cin(t_1184), .o(t_1208), .co(t_1209), .cout(t_1210));
compressor_4_2 u2_421(.a(s_78_5), .b(s_78_4), .c(s_78_3), .d(t_1187), .cin(t_1190), .o(t_1211), .co(t_1212), .cout(t_1213));
compressor_4_2 u2_422(.a(s_78_8), .b(s_78_7), .c(s_78_6), .d(t_1193), .cin(t_1196), .o(t_1214), .co(t_1215), .cout(t_1216));
compressor_4_2 u2_423(.a(s_78_11), .b(s_78_10), .c(s_78_9), .d(t_1199), .cin(t_1202), .o(t_1217), .co(t_1218), .cout(t_1219));
compressor_4_2 u2_424(.a(s_78_14), .b(s_78_13), .c(s_78_12), .d(t_1205), .cin(t_1207), .o(t_1220), .co(t_1221), .cout(t_1222));
compressor_4_2 u2_425(.a(s_78_19), .b(s_78_18), .c(s_78_17), .d(s_78_16), .cin(s_78_15), .o(t_1223), .co(t_1224), .cout(t_1225));
compressor_4_2 u2_426(.a(s_78_24), .b(s_78_23), .c(s_78_22), .d(s_78_21), .cin(s_78_20), .o(t_1226), .co(t_1227), .cout(t_1228));
compressor_4_2 u2_427(.a(s_78_29), .b(s_78_28), .c(s_78_27), .d(s_78_26), .cin(s_78_25), .o(t_1229), .co(t_1230), .cout(t_1231));
compressor_4_2 u2_428(.a(s_78_34), .b(s_78_33), .c(s_78_32), .d(s_78_31), .cin(s_78_30), .o(t_1232), .co(t_1233), .cout(t_1234));
compressor_4_2 u2_429(.a(s_78_39), .b(s_78_38), .c(s_78_37), .d(s_78_36), .cin(s_78_35), .o(t_1235), .co(t_1236), .cout(t_1237));
compressor_4_2 u2_430(.a(s_79_2), .b(s_79_1), .c(s_79_0), .d(t_1210), .cin(t_1213), .o(t_1238), .co(t_1239), .cout(t_1240));
compressor_4_2 u2_431(.a(s_79_5), .b(s_79_4), .c(s_79_3), .d(t_1216), .cin(t_1219), .o(t_1241), .co(t_1242), .cout(t_1243));
compressor_4_2 u2_432(.a(s_79_8), .b(s_79_7), .c(s_79_6), .d(t_1222), .cin(t_1225), .o(t_1244), .co(t_1245), .cout(t_1246));
compressor_4_2 u2_433(.a(s_79_11), .b(s_79_10), .c(s_79_9), .d(t_1228), .cin(t_1231), .o(t_1247), .co(t_1248), .cout(t_1249));
compressor_4_2 u2_434(.a(s_79_14), .b(s_79_13), .c(s_79_12), .d(t_1234), .cin(t_1237), .o(t_1250), .co(t_1251), .cout(t_1252));
compressor_4_2 u2_435(.a(s_79_19), .b(s_79_18), .c(s_79_17), .d(s_79_16), .cin(s_79_15), .o(t_1253), .co(t_1254), .cout(t_1255));
compressor_4_2 u2_436(.a(s_79_24), .b(s_79_23), .c(s_79_22), .d(s_79_21), .cin(s_79_20), .o(t_1256), .co(t_1257), .cout(t_1258));
compressor_4_2 u2_437(.a(s_79_29), .b(s_79_28), .c(s_79_27), .d(s_79_26), .cin(s_79_25), .o(t_1259), .co(t_1260), .cout(t_1261));
compressor_4_2 u2_438(.a(s_79_34), .b(s_79_33), .c(s_79_32), .d(s_79_31), .cin(s_79_30), .o(t_1262), .co(t_1263), .cout(t_1264));
compressor_4_2 u2_439(.a(s_79_39), .b(s_79_38), .c(s_79_37), .d(s_79_36), .cin(s_79_35), .o(t_1265), .co(t_1266), .cout(t_1267));
compressor_4_2 u2_440(.a(s_80_2), .b(s_80_1), .c(s_80_0), .d(t_1240), .cin(t_1243), .o(t_1268), .co(t_1269), .cout(t_1270));
compressor_4_2 u2_441(.a(s_80_5), .b(s_80_4), .c(s_80_3), .d(t_1246), .cin(t_1249), .o(t_1271), .co(t_1272), .cout(t_1273));
compressor_4_2 u2_442(.a(s_80_8), .b(s_80_7), .c(s_80_6), .d(t_1252), .cin(t_1255), .o(t_1274), .co(t_1275), .cout(t_1276));
compressor_4_2 u2_443(.a(s_80_11), .b(s_80_10), .c(s_80_9), .d(t_1258), .cin(t_1261), .o(t_1277), .co(t_1278), .cout(t_1279));
compressor_4_2 u2_444(.a(s_80_14), .b(s_80_13), .c(s_80_12), .d(t_1264), .cin(t_1267), .o(t_1280), .co(t_1281), .cout(t_1282));
compressor_4_2 u2_445(.a(s_80_19), .b(s_80_18), .c(s_80_17), .d(s_80_16), .cin(s_80_15), .o(t_1283), .co(t_1284), .cout(t_1285));
compressor_4_2 u2_446(.a(s_80_24), .b(s_80_23), .c(s_80_22), .d(s_80_21), .cin(s_80_20), .o(t_1286), .co(t_1287), .cout(t_1288));
compressor_4_2 u2_447(.a(s_80_29), .b(s_80_28), .c(s_80_27), .d(s_80_26), .cin(s_80_25), .o(t_1289), .co(t_1290), .cout(t_1291));
compressor_4_2 u2_448(.a(s_80_34), .b(s_80_33), .c(s_80_32), .d(s_80_31), .cin(s_80_30), .o(t_1292), .co(t_1293), .cout(t_1294));
compressor_4_2 u2_449(.a(s_80_39), .b(s_80_38), .c(s_80_37), .d(s_80_36), .cin(s_80_35), .o(t_1295), .co(t_1296), .cout(t_1297));
half_adder u0_450(.a(s_80_41), .b(s_80_40), .o(t_1298), .cout(t_1299));
compressor_4_2 u2_451(.a(s_81_2), .b(s_81_1), .c(s_81_0), .d(t_1270), .cin(t_1273), .o(t_1300), .co(t_1301), .cout(t_1302));
compressor_4_2 u2_452(.a(s_81_5), .b(s_81_4), .c(s_81_3), .d(t_1276), .cin(t_1279), .o(t_1303), .co(t_1304), .cout(t_1305));
compressor_4_2 u2_453(.a(s_81_8), .b(s_81_7), .c(s_81_6), .d(t_1282), .cin(t_1285), .o(t_1306), .co(t_1307), .cout(t_1308));
compressor_4_2 u2_454(.a(s_81_11), .b(s_81_10), .c(s_81_9), .d(t_1288), .cin(t_1291), .o(t_1309), .co(t_1310), .cout(t_1311));
compressor_4_2 u2_455(.a(s_81_14), .b(s_81_13), .c(s_81_12), .d(t_1294), .cin(t_1297), .o(t_1312), .co(t_1313), .cout(t_1314));
compressor_4_2 u2_456(.a(s_81_18), .b(s_81_17), .c(s_81_16), .d(s_81_15), .cin(t_1299), .o(t_1315), .co(t_1316), .cout(t_1317));
compressor_4_2 u2_457(.a(s_81_23), .b(s_81_22), .c(s_81_21), .d(s_81_20), .cin(s_81_19), .o(t_1318), .co(t_1319), .cout(t_1320));
compressor_4_2 u2_458(.a(s_81_28), .b(s_81_27), .c(s_81_26), .d(s_81_25), .cin(s_81_24), .o(t_1321), .co(t_1322), .cout(t_1323));
compressor_4_2 u2_459(.a(s_81_33), .b(s_81_32), .c(s_81_31), .d(s_81_30), .cin(s_81_29), .o(t_1324), .co(t_1325), .cout(t_1326));
compressor_4_2 u2_460(.a(s_81_38), .b(s_81_37), .c(s_81_36), .d(s_81_35), .cin(s_81_34), .o(t_1327), .co(t_1328), .cout(t_1329));
half_adder u0_461(.a(s_81_40), .b(s_81_39), .o(t_1330), .cout(t_1331));
compressor_4_2 u2_462(.a(s_82_2), .b(s_82_1), .c(s_82_0), .d(t_1302), .cin(t_1305), .o(t_1332), .co(t_1333), .cout(t_1334));
compressor_4_2 u2_463(.a(s_82_5), .b(s_82_4), .c(s_82_3), .d(t_1308), .cin(t_1311), .o(t_1335), .co(t_1336), .cout(t_1337));
compressor_4_2 u2_464(.a(s_82_8), .b(s_82_7), .c(s_82_6), .d(t_1314), .cin(t_1317), .o(t_1338), .co(t_1339), .cout(t_1340));
compressor_4_2 u2_465(.a(s_82_11), .b(s_82_10), .c(s_82_9), .d(t_1320), .cin(t_1323), .o(t_1341), .co(t_1342), .cout(t_1343));
compressor_4_2 u2_466(.a(s_82_14), .b(s_82_13), .c(s_82_12), .d(t_1326), .cin(t_1329), .o(t_1344), .co(t_1345), .cout(t_1346));
compressor_4_2 u2_467(.a(s_82_18), .b(s_82_17), .c(s_82_16), .d(s_82_15), .cin(t_1331), .o(t_1347), .co(t_1348), .cout(t_1349));
compressor_4_2 u2_468(.a(s_82_23), .b(s_82_22), .c(s_82_21), .d(s_82_20), .cin(s_82_19), .o(t_1350), .co(t_1351), .cout(t_1352));
compressor_4_2 u2_469(.a(s_82_28), .b(s_82_27), .c(s_82_26), .d(s_82_25), .cin(s_82_24), .o(t_1353), .co(t_1354), .cout(t_1355));
compressor_4_2 u2_470(.a(s_82_33), .b(s_82_32), .c(s_82_31), .d(s_82_30), .cin(s_82_29), .o(t_1356), .co(t_1357), .cout(t_1358));
compressor_4_2 u2_471(.a(s_82_38), .b(s_82_37), .c(s_82_36), .d(s_82_35), .cin(s_82_34), .o(t_1359), .co(t_1360), .cout(t_1361));
compressor_3_2 u1_472(.a(s_82_41), .b(s_82_40), .cin(s_82_39), .o(t_1362), .cout(t_1363));
compressor_4_2 u2_473(.a(s_83_2), .b(s_83_1), .c(s_83_0), .d(t_1334), .cin(t_1337), .o(t_1364), .co(t_1365), .cout(t_1366));
compressor_4_2 u2_474(.a(s_83_5), .b(s_83_4), .c(s_83_3), .d(t_1340), .cin(t_1343), .o(t_1367), .co(t_1368), .cout(t_1369));
compressor_4_2 u2_475(.a(s_83_8), .b(s_83_7), .c(s_83_6), .d(t_1346), .cin(t_1349), .o(t_1370), .co(t_1371), .cout(t_1372));
compressor_4_2 u2_476(.a(s_83_11), .b(s_83_10), .c(s_83_9), .d(t_1352), .cin(t_1355), .o(t_1373), .co(t_1374), .cout(t_1375));
compressor_4_2 u2_477(.a(s_83_14), .b(s_83_13), .c(s_83_12), .d(t_1358), .cin(t_1361), .o(t_1376), .co(t_1377), .cout(t_1378));
compressor_4_2 u2_478(.a(s_83_18), .b(s_83_17), .c(s_83_16), .d(s_83_15), .cin(t_1363), .o(t_1379), .co(t_1380), .cout(t_1381));
compressor_4_2 u2_479(.a(s_83_23), .b(s_83_22), .c(s_83_21), .d(s_83_20), .cin(s_83_19), .o(t_1382), .co(t_1383), .cout(t_1384));
compressor_4_2 u2_480(.a(s_83_28), .b(s_83_27), .c(s_83_26), .d(s_83_25), .cin(s_83_24), .o(t_1385), .co(t_1386), .cout(t_1387));
compressor_4_2 u2_481(.a(s_83_33), .b(s_83_32), .c(s_83_31), .d(s_83_30), .cin(s_83_29), .o(t_1388), .co(t_1389), .cout(t_1390));
compressor_4_2 u2_482(.a(s_83_38), .b(s_83_37), .c(s_83_36), .d(s_83_35), .cin(s_83_34), .o(t_1391), .co(t_1392), .cout(t_1393));
compressor_3_2 u1_483(.a(s_83_41), .b(s_83_40), .cin(s_83_39), .o(t_1394), .cout(t_1395));
compressor_4_2 u2_484(.a(s_84_2), .b(s_84_1), .c(s_84_0), .d(t_1366), .cin(t_1369), .o(t_1396), .co(t_1397), .cout(t_1398));
compressor_4_2 u2_485(.a(s_84_5), .b(s_84_4), .c(s_84_3), .d(t_1372), .cin(t_1375), .o(t_1399), .co(t_1400), .cout(t_1401));
compressor_4_2 u2_486(.a(s_84_8), .b(s_84_7), .c(s_84_6), .d(t_1378), .cin(t_1381), .o(t_1402), .co(t_1403), .cout(t_1404));
compressor_4_2 u2_487(.a(s_84_11), .b(s_84_10), .c(s_84_9), .d(t_1384), .cin(t_1387), .o(t_1405), .co(t_1406), .cout(t_1407));
compressor_4_2 u2_488(.a(s_84_14), .b(s_84_13), .c(s_84_12), .d(t_1390), .cin(t_1393), .o(t_1408), .co(t_1409), .cout(t_1410));
compressor_4_2 u2_489(.a(s_84_18), .b(s_84_17), .c(s_84_16), .d(s_84_15), .cin(t_1395), .o(t_1411), .co(t_1412), .cout(t_1413));
compressor_4_2 u2_490(.a(s_84_23), .b(s_84_22), .c(s_84_21), .d(s_84_20), .cin(s_84_19), .o(t_1414), .co(t_1415), .cout(t_1416));
compressor_4_2 u2_491(.a(s_84_28), .b(s_84_27), .c(s_84_26), .d(s_84_25), .cin(s_84_24), .o(t_1417), .co(t_1418), .cout(t_1419));
compressor_4_2 u2_492(.a(s_84_33), .b(s_84_32), .c(s_84_31), .d(s_84_30), .cin(s_84_29), .o(t_1420), .co(t_1421), .cout(t_1422));
compressor_4_2 u2_493(.a(s_84_38), .b(s_84_37), .c(s_84_36), .d(s_84_35), .cin(s_84_34), .o(t_1423), .co(t_1424), .cout(t_1425));
compressor_4_2 u2_494(.a(s_84_43), .b(s_84_42), .c(s_84_41), .d(s_84_40), .cin(s_84_39), .o(t_1426), .co(t_1427), .cout(t_1428));
compressor_4_2 u2_495(.a(s_85_2), .b(s_85_1), .c(s_85_0), .d(t_1398), .cin(t_1401), .o(t_1429), .co(t_1430), .cout(t_1431));
compressor_4_2 u2_496(.a(s_85_5), .b(s_85_4), .c(s_85_3), .d(t_1404), .cin(t_1407), .o(t_1432), .co(t_1433), .cout(t_1434));
compressor_4_2 u2_497(.a(s_85_8), .b(s_85_7), .c(s_85_6), .d(t_1410), .cin(t_1413), .o(t_1435), .co(t_1436), .cout(t_1437));
compressor_4_2 u2_498(.a(s_85_11), .b(s_85_10), .c(s_85_9), .d(t_1416), .cin(t_1419), .o(t_1438), .co(t_1439), .cout(t_1440));
compressor_4_2 u2_499(.a(s_85_14), .b(s_85_13), .c(s_85_12), .d(t_1422), .cin(t_1425), .o(t_1441), .co(t_1442), .cout(t_1443));
compressor_4_2 u2_500(.a(s_85_18), .b(s_85_17), .c(s_85_16), .d(s_85_15), .cin(t_1428), .o(t_1444), .co(t_1445), .cout(t_1446));
compressor_4_2 u2_501(.a(s_85_23), .b(s_85_22), .c(s_85_21), .d(s_85_20), .cin(s_85_19), .o(t_1447), .co(t_1448), .cout(t_1449));
compressor_4_2 u2_502(.a(s_85_28), .b(s_85_27), .c(s_85_26), .d(s_85_25), .cin(s_85_24), .o(t_1450), .co(t_1451), .cout(t_1452));
compressor_4_2 u2_503(.a(s_85_33), .b(s_85_32), .c(s_85_31), .d(s_85_30), .cin(s_85_29), .o(t_1453), .co(t_1454), .cout(t_1455));
compressor_4_2 u2_504(.a(s_85_38), .b(s_85_37), .c(s_85_36), .d(s_85_35), .cin(s_85_34), .o(t_1456), .co(t_1457), .cout(t_1458));
compressor_3_2 u1_505(.a(s_85_41), .b(s_85_40), .cin(s_85_39), .o(t_1459), .cout(t_1460));
compressor_4_2 u2_506(.a(s_86_2), .b(s_86_1), .c(s_86_0), .d(t_1431), .cin(t_1434), .o(t_1461), .co(t_1462), .cout(t_1463));
compressor_4_2 u2_507(.a(s_86_5), .b(s_86_4), .c(s_86_3), .d(t_1437), .cin(t_1440), .o(t_1464), .co(t_1465), .cout(t_1466));
compressor_4_2 u2_508(.a(s_86_8), .b(s_86_7), .c(s_86_6), .d(t_1443), .cin(t_1446), .o(t_1467), .co(t_1468), .cout(t_1469));
compressor_4_2 u2_509(.a(s_86_11), .b(s_86_10), .c(s_86_9), .d(t_1449), .cin(t_1452), .o(t_1470), .co(t_1471), .cout(t_1472));
compressor_4_2 u2_510(.a(s_86_14), .b(s_86_13), .c(s_86_12), .d(t_1455), .cin(t_1458), .o(t_1473), .co(t_1474), .cout(t_1475));
compressor_4_2 u2_511(.a(s_86_18), .b(s_86_17), .c(s_86_16), .d(s_86_15), .cin(t_1460), .o(t_1476), .co(t_1477), .cout(t_1478));
compressor_4_2 u2_512(.a(s_86_23), .b(s_86_22), .c(s_86_21), .d(s_86_20), .cin(s_86_19), .o(t_1479), .co(t_1480), .cout(t_1481));
compressor_4_2 u2_513(.a(s_86_28), .b(s_86_27), .c(s_86_26), .d(s_86_25), .cin(s_86_24), .o(t_1482), .co(t_1483), .cout(t_1484));
compressor_4_2 u2_514(.a(s_86_33), .b(s_86_32), .c(s_86_31), .d(s_86_30), .cin(s_86_29), .o(t_1485), .co(t_1486), .cout(t_1487));
compressor_4_2 u2_515(.a(s_86_38), .b(s_86_37), .c(s_86_36), .d(s_86_35), .cin(s_86_34), .o(t_1488), .co(t_1489), .cout(t_1490));
compressor_4_2 u2_516(.a(s_86_43), .b(s_86_42), .c(s_86_41), .d(s_86_40), .cin(s_86_39), .o(t_1491), .co(t_1492), .cout(t_1493));
compressor_4_2 u2_517(.a(s_87_2), .b(s_87_1), .c(s_87_0), .d(t_1463), .cin(t_1466), .o(t_1494), .co(t_1495), .cout(t_1496));
compressor_4_2 u2_518(.a(s_87_5), .b(s_87_4), .c(s_87_3), .d(t_1469), .cin(t_1472), .o(t_1497), .co(t_1498), .cout(t_1499));
compressor_4_2 u2_519(.a(s_87_8), .b(s_87_7), .c(s_87_6), .d(t_1475), .cin(t_1478), .o(t_1500), .co(t_1501), .cout(t_1502));
compressor_4_2 u2_520(.a(s_87_11), .b(s_87_10), .c(s_87_9), .d(t_1481), .cin(t_1484), .o(t_1503), .co(t_1504), .cout(t_1505));
compressor_4_2 u2_521(.a(s_87_14), .b(s_87_13), .c(s_87_12), .d(t_1487), .cin(t_1490), .o(t_1506), .co(t_1507), .cout(t_1508));
compressor_4_2 u2_522(.a(s_87_18), .b(s_87_17), .c(s_87_16), .d(s_87_15), .cin(t_1493), .o(t_1509), .co(t_1510), .cout(t_1511));
compressor_4_2 u2_523(.a(s_87_23), .b(s_87_22), .c(s_87_21), .d(s_87_20), .cin(s_87_19), .o(t_1512), .co(t_1513), .cout(t_1514));
compressor_4_2 u2_524(.a(s_87_28), .b(s_87_27), .c(s_87_26), .d(s_87_25), .cin(s_87_24), .o(t_1515), .co(t_1516), .cout(t_1517));
compressor_4_2 u2_525(.a(s_87_33), .b(s_87_32), .c(s_87_31), .d(s_87_30), .cin(s_87_29), .o(t_1518), .co(t_1519), .cout(t_1520));
compressor_4_2 u2_526(.a(s_87_38), .b(s_87_37), .c(s_87_36), .d(s_87_35), .cin(s_87_34), .o(t_1521), .co(t_1522), .cout(t_1523));
compressor_4_2 u2_527(.a(s_87_43), .b(s_87_42), .c(s_87_41), .d(s_87_40), .cin(s_87_39), .o(t_1524), .co(t_1525), .cout(t_1526));
compressor_4_2 u2_528(.a(s_88_2), .b(s_88_1), .c(s_88_0), .d(t_1496), .cin(t_1499), .o(t_1527), .co(t_1528), .cout(t_1529));
compressor_4_2 u2_529(.a(s_88_5), .b(s_88_4), .c(s_88_3), .d(t_1502), .cin(t_1505), .o(t_1530), .co(t_1531), .cout(t_1532));
compressor_4_2 u2_530(.a(s_88_8), .b(s_88_7), .c(s_88_6), .d(t_1508), .cin(t_1511), .o(t_1533), .co(t_1534), .cout(t_1535));
compressor_4_2 u2_531(.a(s_88_11), .b(s_88_10), .c(s_88_9), .d(t_1514), .cin(t_1517), .o(t_1536), .co(t_1537), .cout(t_1538));
compressor_4_2 u2_532(.a(s_88_14), .b(s_88_13), .c(s_88_12), .d(t_1520), .cin(t_1523), .o(t_1539), .co(t_1540), .cout(t_1541));
compressor_4_2 u2_533(.a(s_88_18), .b(s_88_17), .c(s_88_16), .d(s_88_15), .cin(t_1526), .o(t_1542), .co(t_1543), .cout(t_1544));
compressor_4_2 u2_534(.a(s_88_23), .b(s_88_22), .c(s_88_21), .d(s_88_20), .cin(s_88_19), .o(t_1545), .co(t_1546), .cout(t_1547));
compressor_4_2 u2_535(.a(s_88_28), .b(s_88_27), .c(s_88_26), .d(s_88_25), .cin(s_88_24), .o(t_1548), .co(t_1549), .cout(t_1550));
compressor_4_2 u2_536(.a(s_88_33), .b(s_88_32), .c(s_88_31), .d(s_88_30), .cin(s_88_29), .o(t_1551), .co(t_1552), .cout(t_1553));
compressor_4_2 u2_537(.a(s_88_38), .b(s_88_37), .c(s_88_36), .d(s_88_35), .cin(s_88_34), .o(t_1554), .co(t_1555), .cout(t_1556));
compressor_4_2 u2_538(.a(s_88_43), .b(s_88_42), .c(s_88_41), .d(s_88_40), .cin(s_88_39), .o(t_1557), .co(t_1558), .cout(t_1559));
half_adder u0_539(.a(s_88_45), .b(s_88_44), .o(t_1560), .cout(t_1561));
compressor_4_2 u2_540(.a(s_89_2), .b(s_89_1), .c(s_89_0), .d(t_1529), .cin(t_1532), .o(t_1562), .co(t_1563), .cout(t_1564));
compressor_4_2 u2_541(.a(s_89_5), .b(s_89_4), .c(s_89_3), .d(t_1535), .cin(t_1538), .o(t_1565), .co(t_1566), .cout(t_1567));
compressor_4_2 u2_542(.a(s_89_8), .b(s_89_7), .c(s_89_6), .d(t_1541), .cin(t_1544), .o(t_1568), .co(t_1569), .cout(t_1570));
compressor_4_2 u2_543(.a(s_89_11), .b(s_89_10), .c(s_89_9), .d(t_1547), .cin(t_1550), .o(t_1571), .co(t_1572), .cout(t_1573));
compressor_4_2 u2_544(.a(s_89_14), .b(s_89_13), .c(s_89_12), .d(t_1553), .cin(t_1556), .o(t_1574), .co(t_1575), .cout(t_1576));
compressor_4_2 u2_545(.a(s_89_17), .b(s_89_16), .c(s_89_15), .d(t_1559), .cin(t_1561), .o(t_1577), .co(t_1578), .cout(t_1579));
compressor_4_2 u2_546(.a(s_89_22), .b(s_89_21), .c(s_89_20), .d(s_89_19), .cin(s_89_18), .o(t_1580), .co(t_1581), .cout(t_1582));
compressor_4_2 u2_547(.a(s_89_27), .b(s_89_26), .c(s_89_25), .d(s_89_24), .cin(s_89_23), .o(t_1583), .co(t_1584), .cout(t_1585));
compressor_4_2 u2_548(.a(s_89_32), .b(s_89_31), .c(s_89_30), .d(s_89_29), .cin(s_89_28), .o(t_1586), .co(t_1587), .cout(t_1588));
compressor_4_2 u2_549(.a(s_89_37), .b(s_89_36), .c(s_89_35), .d(s_89_34), .cin(s_89_33), .o(t_1589), .co(t_1590), .cout(t_1591));
compressor_4_2 u2_550(.a(s_89_42), .b(s_89_41), .c(s_89_40), .d(s_89_39), .cin(s_89_38), .o(t_1592), .co(t_1593), .cout(t_1594));
half_adder u0_551(.a(s_89_44), .b(s_89_43), .o(t_1595), .cout(t_1596));
compressor_4_2 u2_552(.a(s_90_2), .b(s_90_1), .c(s_90_0), .d(t_1564), .cin(t_1567), .o(t_1597), .co(t_1598), .cout(t_1599));
compressor_4_2 u2_553(.a(s_90_5), .b(s_90_4), .c(s_90_3), .d(t_1570), .cin(t_1573), .o(t_1600), .co(t_1601), .cout(t_1602));
compressor_4_2 u2_554(.a(s_90_8), .b(s_90_7), .c(s_90_6), .d(t_1576), .cin(t_1579), .o(t_1603), .co(t_1604), .cout(t_1605));
compressor_4_2 u2_555(.a(s_90_11), .b(s_90_10), .c(s_90_9), .d(t_1582), .cin(t_1585), .o(t_1606), .co(t_1607), .cout(t_1608));
compressor_4_2 u2_556(.a(s_90_14), .b(s_90_13), .c(s_90_12), .d(t_1588), .cin(t_1591), .o(t_1609), .co(t_1610), .cout(t_1611));
compressor_4_2 u2_557(.a(s_90_17), .b(s_90_16), .c(s_90_15), .d(t_1594), .cin(t_1596), .o(t_1612), .co(t_1613), .cout(t_1614));
compressor_4_2 u2_558(.a(s_90_22), .b(s_90_21), .c(s_90_20), .d(s_90_19), .cin(s_90_18), .o(t_1615), .co(t_1616), .cout(t_1617));
compressor_4_2 u2_559(.a(s_90_27), .b(s_90_26), .c(s_90_25), .d(s_90_24), .cin(s_90_23), .o(t_1618), .co(t_1619), .cout(t_1620));
compressor_4_2 u2_560(.a(s_90_32), .b(s_90_31), .c(s_90_30), .d(s_90_29), .cin(s_90_28), .o(t_1621), .co(t_1622), .cout(t_1623));
compressor_4_2 u2_561(.a(s_90_37), .b(s_90_36), .c(s_90_35), .d(s_90_34), .cin(s_90_33), .o(t_1624), .co(t_1625), .cout(t_1626));
compressor_4_2 u2_562(.a(s_90_42), .b(s_90_41), .c(s_90_40), .d(s_90_39), .cin(s_90_38), .o(t_1627), .co(t_1628), .cout(t_1629));
compressor_3_2 u1_563(.a(s_90_45), .b(s_90_44), .cin(s_90_43), .o(t_1630), .cout(t_1631));
compressor_4_2 u2_564(.a(s_91_2), .b(s_91_1), .c(s_91_0), .d(t_1599), .cin(t_1602), .o(t_1632), .co(t_1633), .cout(t_1634));
compressor_4_2 u2_565(.a(s_91_5), .b(s_91_4), .c(s_91_3), .d(t_1605), .cin(t_1608), .o(t_1635), .co(t_1636), .cout(t_1637));
compressor_4_2 u2_566(.a(s_91_8), .b(s_91_7), .c(s_91_6), .d(t_1611), .cin(t_1614), .o(t_1638), .co(t_1639), .cout(t_1640));
compressor_4_2 u2_567(.a(s_91_11), .b(s_91_10), .c(s_91_9), .d(t_1617), .cin(t_1620), .o(t_1641), .co(t_1642), .cout(t_1643));
compressor_4_2 u2_568(.a(s_91_14), .b(s_91_13), .c(s_91_12), .d(t_1623), .cin(t_1626), .o(t_1644), .co(t_1645), .cout(t_1646));
compressor_4_2 u2_569(.a(s_91_17), .b(s_91_16), .c(s_91_15), .d(t_1629), .cin(t_1631), .o(t_1647), .co(t_1648), .cout(t_1649));
compressor_4_2 u2_570(.a(s_91_22), .b(s_91_21), .c(s_91_20), .d(s_91_19), .cin(s_91_18), .o(t_1650), .co(t_1651), .cout(t_1652));
compressor_4_2 u2_571(.a(s_91_27), .b(s_91_26), .c(s_91_25), .d(s_91_24), .cin(s_91_23), .o(t_1653), .co(t_1654), .cout(t_1655));
compressor_4_2 u2_572(.a(s_91_32), .b(s_91_31), .c(s_91_30), .d(s_91_29), .cin(s_91_28), .o(t_1656), .co(t_1657), .cout(t_1658));
compressor_4_2 u2_573(.a(s_91_37), .b(s_91_36), .c(s_91_35), .d(s_91_34), .cin(s_91_33), .o(t_1659), .co(t_1660), .cout(t_1661));
compressor_4_2 u2_574(.a(s_91_42), .b(s_91_41), .c(s_91_40), .d(s_91_39), .cin(s_91_38), .o(t_1662), .co(t_1663), .cout(t_1664));
compressor_3_2 u1_575(.a(s_91_45), .b(s_91_44), .cin(s_91_43), .o(t_1665), .cout(t_1666));
compressor_4_2 u2_576(.a(s_92_2), .b(s_92_1), .c(s_92_0), .d(t_1634), .cin(t_1637), .o(t_1667), .co(t_1668), .cout(t_1669));
compressor_4_2 u2_577(.a(s_92_5), .b(s_92_4), .c(s_92_3), .d(t_1640), .cin(t_1643), .o(t_1670), .co(t_1671), .cout(t_1672));
compressor_4_2 u2_578(.a(s_92_8), .b(s_92_7), .c(s_92_6), .d(t_1646), .cin(t_1649), .o(t_1673), .co(t_1674), .cout(t_1675));
compressor_4_2 u2_579(.a(s_92_11), .b(s_92_10), .c(s_92_9), .d(t_1652), .cin(t_1655), .o(t_1676), .co(t_1677), .cout(t_1678));
compressor_4_2 u2_580(.a(s_92_14), .b(s_92_13), .c(s_92_12), .d(t_1658), .cin(t_1661), .o(t_1679), .co(t_1680), .cout(t_1681));
compressor_4_2 u2_581(.a(s_92_17), .b(s_92_16), .c(s_92_15), .d(t_1664), .cin(t_1666), .o(t_1682), .co(t_1683), .cout(t_1684));
compressor_4_2 u2_582(.a(s_92_22), .b(s_92_21), .c(s_92_20), .d(s_92_19), .cin(s_92_18), .o(t_1685), .co(t_1686), .cout(t_1687));
compressor_4_2 u2_583(.a(s_92_27), .b(s_92_26), .c(s_92_25), .d(s_92_24), .cin(s_92_23), .o(t_1688), .co(t_1689), .cout(t_1690));
compressor_4_2 u2_584(.a(s_92_32), .b(s_92_31), .c(s_92_30), .d(s_92_29), .cin(s_92_28), .o(t_1691), .co(t_1692), .cout(t_1693));
compressor_4_2 u2_585(.a(s_92_37), .b(s_92_36), .c(s_92_35), .d(s_92_34), .cin(s_92_33), .o(t_1694), .co(t_1695), .cout(t_1696));
compressor_4_2 u2_586(.a(s_92_42), .b(s_92_41), .c(s_92_40), .d(s_92_39), .cin(s_92_38), .o(t_1697), .co(t_1698), .cout(t_1699));
compressor_4_2 u2_587(.a(s_92_47), .b(s_92_46), .c(s_92_45), .d(s_92_44), .cin(s_92_43), .o(t_1700), .co(t_1701), .cout(t_1702));
compressor_4_2 u2_588(.a(s_93_2), .b(s_93_1), .c(s_93_0), .d(t_1669), .cin(t_1672), .o(t_1703), .co(t_1704), .cout(t_1705));
compressor_4_2 u2_589(.a(s_93_5), .b(s_93_4), .c(s_93_3), .d(t_1675), .cin(t_1678), .o(t_1706), .co(t_1707), .cout(t_1708));
compressor_4_2 u2_590(.a(s_93_8), .b(s_93_7), .c(s_93_6), .d(t_1681), .cin(t_1684), .o(t_1709), .co(t_1710), .cout(t_1711));
compressor_4_2 u2_591(.a(s_93_11), .b(s_93_10), .c(s_93_9), .d(t_1687), .cin(t_1690), .o(t_1712), .co(t_1713), .cout(t_1714));
compressor_4_2 u2_592(.a(s_93_14), .b(s_93_13), .c(s_93_12), .d(t_1693), .cin(t_1696), .o(t_1715), .co(t_1716), .cout(t_1717));
compressor_4_2 u2_593(.a(s_93_17), .b(s_93_16), .c(s_93_15), .d(t_1699), .cin(t_1702), .o(t_1718), .co(t_1719), .cout(t_1720));
compressor_4_2 u2_594(.a(s_93_22), .b(s_93_21), .c(s_93_20), .d(s_93_19), .cin(s_93_18), .o(t_1721), .co(t_1722), .cout(t_1723));
compressor_4_2 u2_595(.a(s_93_27), .b(s_93_26), .c(s_93_25), .d(s_93_24), .cin(s_93_23), .o(t_1724), .co(t_1725), .cout(t_1726));
compressor_4_2 u2_596(.a(s_93_32), .b(s_93_31), .c(s_93_30), .d(s_93_29), .cin(s_93_28), .o(t_1727), .co(t_1728), .cout(t_1729));
compressor_4_2 u2_597(.a(s_93_37), .b(s_93_36), .c(s_93_35), .d(s_93_34), .cin(s_93_33), .o(t_1730), .co(t_1731), .cout(t_1732));
compressor_4_2 u2_598(.a(s_93_42), .b(s_93_41), .c(s_93_40), .d(s_93_39), .cin(s_93_38), .o(t_1733), .co(t_1734), .cout(t_1735));
compressor_3_2 u1_599(.a(s_93_45), .b(s_93_44), .cin(s_93_43), .o(t_1736), .cout(t_1737));
compressor_4_2 u2_600(.a(s_94_2), .b(s_94_1), .c(s_94_0), .d(t_1705), .cin(t_1708), .o(t_1738), .co(t_1739), .cout(t_1740));
compressor_4_2 u2_601(.a(s_94_5), .b(s_94_4), .c(s_94_3), .d(t_1711), .cin(t_1714), .o(t_1741), .co(t_1742), .cout(t_1743));
compressor_4_2 u2_602(.a(s_94_8), .b(s_94_7), .c(s_94_6), .d(t_1717), .cin(t_1720), .o(t_1744), .co(t_1745), .cout(t_1746));
compressor_4_2 u2_603(.a(s_94_11), .b(s_94_10), .c(s_94_9), .d(t_1723), .cin(t_1726), .o(t_1747), .co(t_1748), .cout(t_1749));
compressor_4_2 u2_604(.a(s_94_14), .b(s_94_13), .c(s_94_12), .d(t_1729), .cin(t_1732), .o(t_1750), .co(t_1751), .cout(t_1752));
compressor_4_2 u2_605(.a(s_94_17), .b(s_94_16), .c(s_94_15), .d(t_1735), .cin(t_1737), .o(t_1753), .co(t_1754), .cout(t_1755));
compressor_4_2 u2_606(.a(s_94_22), .b(s_94_21), .c(s_94_20), .d(s_94_19), .cin(s_94_18), .o(t_1756), .co(t_1757), .cout(t_1758));
compressor_4_2 u2_607(.a(s_94_27), .b(s_94_26), .c(s_94_25), .d(s_94_24), .cin(s_94_23), .o(t_1759), .co(t_1760), .cout(t_1761));
compressor_4_2 u2_608(.a(s_94_32), .b(s_94_31), .c(s_94_30), .d(s_94_29), .cin(s_94_28), .o(t_1762), .co(t_1763), .cout(t_1764));
compressor_4_2 u2_609(.a(s_94_37), .b(s_94_36), .c(s_94_35), .d(s_94_34), .cin(s_94_33), .o(t_1765), .co(t_1766), .cout(t_1767));
compressor_4_2 u2_610(.a(s_94_42), .b(s_94_41), .c(s_94_40), .d(s_94_39), .cin(s_94_38), .o(t_1768), .co(t_1769), .cout(t_1770));
compressor_4_2 u2_611(.a(s_94_47), .b(s_94_46), .c(s_94_45), .d(s_94_44), .cin(s_94_43), .o(t_1771), .co(t_1772), .cout(t_1773));
compressor_4_2 u2_612(.a(s_95_2), .b(s_95_1), .c(s_95_0), .d(t_1740), .cin(t_1743), .o(t_1774), .co(t_1775), .cout(t_1776));
compressor_4_2 u2_613(.a(s_95_5), .b(s_95_4), .c(s_95_3), .d(t_1746), .cin(t_1749), .o(t_1777), .co(t_1778), .cout(t_1779));
compressor_4_2 u2_614(.a(s_95_8), .b(s_95_7), .c(s_95_6), .d(t_1752), .cin(t_1755), .o(t_1780), .co(t_1781), .cout(t_1782));
compressor_4_2 u2_615(.a(s_95_11), .b(s_95_10), .c(s_95_9), .d(t_1758), .cin(t_1761), .o(t_1783), .co(t_1784), .cout(t_1785));
compressor_4_2 u2_616(.a(s_95_14), .b(s_95_13), .c(s_95_12), .d(t_1764), .cin(t_1767), .o(t_1786), .co(t_1787), .cout(t_1788));
compressor_4_2 u2_617(.a(s_95_17), .b(s_95_16), .c(s_95_15), .d(t_1770), .cin(t_1773), .o(t_1789), .co(t_1790), .cout(t_1791));
compressor_4_2 u2_618(.a(s_95_22), .b(s_95_21), .c(s_95_20), .d(s_95_19), .cin(s_95_18), .o(t_1792), .co(t_1793), .cout(t_1794));
compressor_4_2 u2_619(.a(s_95_27), .b(s_95_26), .c(s_95_25), .d(s_95_24), .cin(s_95_23), .o(t_1795), .co(t_1796), .cout(t_1797));
compressor_4_2 u2_620(.a(s_95_32), .b(s_95_31), .c(s_95_30), .d(s_95_29), .cin(s_95_28), .o(t_1798), .co(t_1799), .cout(t_1800));
compressor_4_2 u2_621(.a(s_95_37), .b(s_95_36), .c(s_95_35), .d(s_95_34), .cin(s_95_33), .o(t_1801), .co(t_1802), .cout(t_1803));
compressor_4_2 u2_622(.a(s_95_42), .b(s_95_41), .c(s_95_40), .d(s_95_39), .cin(s_95_38), .o(t_1804), .co(t_1805), .cout(t_1806));
compressor_4_2 u2_623(.a(s_95_47), .b(s_95_46), .c(s_95_45), .d(s_95_44), .cin(s_95_43), .o(t_1807), .co(t_1808), .cout(t_1809));
compressor_4_2 u2_624(.a(s_96_2), .b(s_96_1), .c(s_96_0), .d(t_1776), .cin(t_1779), .o(t_1810), .co(t_1811), .cout(t_1812));
compressor_4_2 u2_625(.a(s_96_5), .b(s_96_4), .c(s_96_3), .d(t_1782), .cin(t_1785), .o(t_1813), .co(t_1814), .cout(t_1815));
compressor_4_2 u2_626(.a(s_96_8), .b(s_96_7), .c(s_96_6), .d(t_1788), .cin(t_1791), .o(t_1816), .co(t_1817), .cout(t_1818));
compressor_4_2 u2_627(.a(s_96_11), .b(s_96_10), .c(s_96_9), .d(t_1794), .cin(t_1797), .o(t_1819), .co(t_1820), .cout(t_1821));
compressor_4_2 u2_628(.a(s_96_14), .b(s_96_13), .c(s_96_12), .d(t_1800), .cin(t_1803), .o(t_1822), .co(t_1823), .cout(t_1824));
compressor_4_2 u2_629(.a(s_96_17), .b(s_96_16), .c(s_96_15), .d(t_1806), .cin(t_1809), .o(t_1825), .co(t_1826), .cout(t_1827));
compressor_4_2 u2_630(.a(s_96_22), .b(s_96_21), .c(s_96_20), .d(s_96_19), .cin(s_96_18), .o(t_1828), .co(t_1829), .cout(t_1830));
compressor_4_2 u2_631(.a(s_96_27), .b(s_96_26), .c(s_96_25), .d(s_96_24), .cin(s_96_23), .o(t_1831), .co(t_1832), .cout(t_1833));
compressor_4_2 u2_632(.a(s_96_32), .b(s_96_31), .c(s_96_30), .d(s_96_29), .cin(s_96_28), .o(t_1834), .co(t_1835), .cout(t_1836));
compressor_4_2 u2_633(.a(s_96_37), .b(s_96_36), .c(s_96_35), .d(s_96_34), .cin(s_96_33), .o(t_1837), .co(t_1838), .cout(t_1839));
compressor_4_2 u2_634(.a(s_96_42), .b(s_96_41), .c(s_96_40), .d(s_96_39), .cin(s_96_38), .o(t_1840), .co(t_1841), .cout(t_1842));
compressor_4_2 u2_635(.a(s_96_47), .b(s_96_46), .c(s_96_45), .d(s_96_44), .cin(s_96_43), .o(t_1843), .co(t_1844), .cout(t_1845));
half_adder u0_636(.a(s_96_49), .b(s_96_48), .o(t_1846), .cout(t_1847));
compressor_4_2 u2_637(.a(s_97_2), .b(s_97_1), .c(s_97_0), .d(t_1812), .cin(t_1815), .o(t_1848), .co(t_1849), .cout(t_1850));
compressor_4_2 u2_638(.a(s_97_5), .b(s_97_4), .c(s_97_3), .d(t_1818), .cin(t_1821), .o(t_1851), .co(t_1852), .cout(t_1853));
compressor_4_2 u2_639(.a(s_97_8), .b(s_97_7), .c(s_97_6), .d(t_1824), .cin(t_1827), .o(t_1854), .co(t_1855), .cout(t_1856));
compressor_4_2 u2_640(.a(s_97_11), .b(s_97_10), .c(s_97_9), .d(t_1830), .cin(t_1833), .o(t_1857), .co(t_1858), .cout(t_1859));
compressor_4_2 u2_641(.a(s_97_14), .b(s_97_13), .c(s_97_12), .d(t_1836), .cin(t_1839), .o(t_1860), .co(t_1861), .cout(t_1862));
compressor_4_2 u2_642(.a(s_97_17), .b(s_97_16), .c(s_97_15), .d(t_1842), .cin(t_1845), .o(t_1863), .co(t_1864), .cout(t_1865));
compressor_4_2 u2_643(.a(s_97_21), .b(s_97_20), .c(s_97_19), .d(s_97_18), .cin(t_1847), .o(t_1866), .co(t_1867), .cout(t_1868));
compressor_4_2 u2_644(.a(s_97_26), .b(s_97_25), .c(s_97_24), .d(s_97_23), .cin(s_97_22), .o(t_1869), .co(t_1870), .cout(t_1871));
compressor_4_2 u2_645(.a(s_97_31), .b(s_97_30), .c(s_97_29), .d(s_97_28), .cin(s_97_27), .o(t_1872), .co(t_1873), .cout(t_1874));
compressor_4_2 u2_646(.a(s_97_36), .b(s_97_35), .c(s_97_34), .d(s_97_33), .cin(s_97_32), .o(t_1875), .co(t_1876), .cout(t_1877));
compressor_4_2 u2_647(.a(s_97_41), .b(s_97_40), .c(s_97_39), .d(s_97_38), .cin(s_97_37), .o(t_1878), .co(t_1879), .cout(t_1880));
compressor_4_2 u2_648(.a(s_97_46), .b(s_97_45), .c(s_97_44), .d(s_97_43), .cin(s_97_42), .o(t_1881), .co(t_1882), .cout(t_1883));
half_adder u0_649(.a(s_97_48), .b(s_97_47), .o(t_1884), .cout(t_1885));
compressor_4_2 u2_650(.a(s_98_2), .b(s_98_1), .c(s_98_0), .d(t_1850), .cin(t_1853), .o(t_1886), .co(t_1887), .cout(t_1888));
compressor_4_2 u2_651(.a(s_98_5), .b(s_98_4), .c(s_98_3), .d(t_1856), .cin(t_1859), .o(t_1889), .co(t_1890), .cout(t_1891));
compressor_4_2 u2_652(.a(s_98_8), .b(s_98_7), .c(s_98_6), .d(t_1862), .cin(t_1865), .o(t_1892), .co(t_1893), .cout(t_1894));
compressor_4_2 u2_653(.a(s_98_11), .b(s_98_10), .c(s_98_9), .d(t_1868), .cin(t_1871), .o(t_1895), .co(t_1896), .cout(t_1897));
compressor_4_2 u2_654(.a(s_98_14), .b(s_98_13), .c(s_98_12), .d(t_1874), .cin(t_1877), .o(t_1898), .co(t_1899), .cout(t_1900));
compressor_4_2 u2_655(.a(s_98_17), .b(s_98_16), .c(s_98_15), .d(t_1880), .cin(t_1883), .o(t_1901), .co(t_1902), .cout(t_1903));
compressor_4_2 u2_656(.a(s_98_21), .b(s_98_20), .c(s_98_19), .d(s_98_18), .cin(t_1885), .o(t_1904), .co(t_1905), .cout(t_1906));
compressor_4_2 u2_657(.a(s_98_26), .b(s_98_25), .c(s_98_24), .d(s_98_23), .cin(s_98_22), .o(t_1907), .co(t_1908), .cout(t_1909));
compressor_4_2 u2_658(.a(s_98_31), .b(s_98_30), .c(s_98_29), .d(s_98_28), .cin(s_98_27), .o(t_1910), .co(t_1911), .cout(t_1912));
compressor_4_2 u2_659(.a(s_98_36), .b(s_98_35), .c(s_98_34), .d(s_98_33), .cin(s_98_32), .o(t_1913), .co(t_1914), .cout(t_1915));
compressor_4_2 u2_660(.a(s_98_41), .b(s_98_40), .c(s_98_39), .d(s_98_38), .cin(s_98_37), .o(t_1916), .co(t_1917), .cout(t_1918));
compressor_4_2 u2_661(.a(s_98_46), .b(s_98_45), .c(s_98_44), .d(s_98_43), .cin(s_98_42), .o(t_1919), .co(t_1920), .cout(t_1921));
compressor_3_2 u1_662(.a(s_98_49), .b(s_98_48), .cin(s_98_47), .o(t_1922), .cout(t_1923));
compressor_4_2 u2_663(.a(s_99_2), .b(s_99_1), .c(s_99_0), .d(t_1888), .cin(t_1891), .o(t_1924), .co(t_1925), .cout(t_1926));
compressor_4_2 u2_664(.a(s_99_5), .b(s_99_4), .c(s_99_3), .d(t_1894), .cin(t_1897), .o(t_1927), .co(t_1928), .cout(t_1929));
compressor_4_2 u2_665(.a(s_99_8), .b(s_99_7), .c(s_99_6), .d(t_1900), .cin(t_1903), .o(t_1930), .co(t_1931), .cout(t_1932));
compressor_4_2 u2_666(.a(s_99_11), .b(s_99_10), .c(s_99_9), .d(t_1906), .cin(t_1909), .o(t_1933), .co(t_1934), .cout(t_1935));
compressor_4_2 u2_667(.a(s_99_14), .b(s_99_13), .c(s_99_12), .d(t_1912), .cin(t_1915), .o(t_1936), .co(t_1937), .cout(t_1938));
compressor_4_2 u2_668(.a(s_99_17), .b(s_99_16), .c(s_99_15), .d(t_1918), .cin(t_1921), .o(t_1939), .co(t_1940), .cout(t_1941));
compressor_4_2 u2_669(.a(s_99_21), .b(s_99_20), .c(s_99_19), .d(s_99_18), .cin(t_1923), .o(t_1942), .co(t_1943), .cout(t_1944));
compressor_4_2 u2_670(.a(s_99_26), .b(s_99_25), .c(s_99_24), .d(s_99_23), .cin(s_99_22), .o(t_1945), .co(t_1946), .cout(t_1947));
compressor_4_2 u2_671(.a(s_99_31), .b(s_99_30), .c(s_99_29), .d(s_99_28), .cin(s_99_27), .o(t_1948), .co(t_1949), .cout(t_1950));
compressor_4_2 u2_672(.a(s_99_36), .b(s_99_35), .c(s_99_34), .d(s_99_33), .cin(s_99_32), .o(t_1951), .co(t_1952), .cout(t_1953));
compressor_4_2 u2_673(.a(s_99_41), .b(s_99_40), .c(s_99_39), .d(s_99_38), .cin(s_99_37), .o(t_1954), .co(t_1955), .cout(t_1956));
compressor_4_2 u2_674(.a(s_99_46), .b(s_99_45), .c(s_99_44), .d(s_99_43), .cin(s_99_42), .o(t_1957), .co(t_1958), .cout(t_1959));
compressor_3_2 u1_675(.a(s_99_49), .b(s_99_48), .cin(s_99_47), .o(t_1960), .cout(t_1961));
compressor_4_2 u2_676(.a(s_100_2), .b(s_100_1), .c(s_100_0), .d(t_1926), .cin(t_1929), .o(t_1962), .co(t_1963), .cout(t_1964));
compressor_4_2 u2_677(.a(s_100_5), .b(s_100_4), .c(s_100_3), .d(t_1932), .cin(t_1935), .o(t_1965), .co(t_1966), .cout(t_1967));
compressor_4_2 u2_678(.a(s_100_8), .b(s_100_7), .c(s_100_6), .d(t_1938), .cin(t_1941), .o(t_1968), .co(t_1969), .cout(t_1970));
compressor_4_2 u2_679(.a(s_100_11), .b(s_100_10), .c(s_100_9), .d(t_1944), .cin(t_1947), .o(t_1971), .co(t_1972), .cout(t_1973));
compressor_4_2 u2_680(.a(s_100_14), .b(s_100_13), .c(s_100_12), .d(t_1950), .cin(t_1953), .o(t_1974), .co(t_1975), .cout(t_1976));
compressor_4_2 u2_681(.a(s_100_17), .b(s_100_16), .c(s_100_15), .d(t_1956), .cin(t_1959), .o(t_1977), .co(t_1978), .cout(t_1979));
compressor_4_2 u2_682(.a(s_100_21), .b(s_100_20), .c(s_100_19), .d(s_100_18), .cin(t_1961), .o(t_1980), .co(t_1981), .cout(t_1982));
compressor_4_2 u2_683(.a(s_100_26), .b(s_100_25), .c(s_100_24), .d(s_100_23), .cin(s_100_22), .o(t_1983), .co(t_1984), .cout(t_1985));
compressor_4_2 u2_684(.a(s_100_31), .b(s_100_30), .c(s_100_29), .d(s_100_28), .cin(s_100_27), .o(t_1986), .co(t_1987), .cout(t_1988));
compressor_4_2 u2_685(.a(s_100_36), .b(s_100_35), .c(s_100_34), .d(s_100_33), .cin(s_100_32), .o(t_1989), .co(t_1990), .cout(t_1991));
compressor_4_2 u2_686(.a(s_100_41), .b(s_100_40), .c(s_100_39), .d(s_100_38), .cin(s_100_37), .o(t_1992), .co(t_1993), .cout(t_1994));
compressor_4_2 u2_687(.a(s_100_46), .b(s_100_45), .c(s_100_44), .d(s_100_43), .cin(s_100_42), .o(t_1995), .co(t_1996), .cout(t_1997));
compressor_4_2 u2_688(.a(s_100_51), .b(s_100_50), .c(s_100_49), .d(s_100_48), .cin(s_100_47), .o(t_1998), .co(t_1999), .cout(t_2000));
compressor_4_2 u2_689(.a(s_101_2), .b(s_101_1), .c(s_101_0), .d(t_1964), .cin(t_1967), .o(t_2001), .co(t_2002), .cout(t_2003));
compressor_4_2 u2_690(.a(s_101_5), .b(s_101_4), .c(s_101_3), .d(t_1970), .cin(t_1973), .o(t_2004), .co(t_2005), .cout(t_2006));
compressor_4_2 u2_691(.a(s_101_8), .b(s_101_7), .c(s_101_6), .d(t_1976), .cin(t_1979), .o(t_2007), .co(t_2008), .cout(t_2009));
compressor_4_2 u2_692(.a(s_101_11), .b(s_101_10), .c(s_101_9), .d(t_1982), .cin(t_1985), .o(t_2010), .co(t_2011), .cout(t_2012));
compressor_4_2 u2_693(.a(s_101_14), .b(s_101_13), .c(s_101_12), .d(t_1988), .cin(t_1991), .o(t_2013), .co(t_2014), .cout(t_2015));
compressor_4_2 u2_694(.a(s_101_17), .b(s_101_16), .c(s_101_15), .d(t_1994), .cin(t_1997), .o(t_2016), .co(t_2017), .cout(t_2018));
compressor_4_2 u2_695(.a(s_101_21), .b(s_101_20), .c(s_101_19), .d(s_101_18), .cin(t_2000), .o(t_2019), .co(t_2020), .cout(t_2021));
compressor_4_2 u2_696(.a(s_101_26), .b(s_101_25), .c(s_101_24), .d(s_101_23), .cin(s_101_22), .o(t_2022), .co(t_2023), .cout(t_2024));
compressor_4_2 u2_697(.a(s_101_31), .b(s_101_30), .c(s_101_29), .d(s_101_28), .cin(s_101_27), .o(t_2025), .co(t_2026), .cout(t_2027));
compressor_4_2 u2_698(.a(s_101_36), .b(s_101_35), .c(s_101_34), .d(s_101_33), .cin(s_101_32), .o(t_2028), .co(t_2029), .cout(t_2030));
compressor_4_2 u2_699(.a(s_101_41), .b(s_101_40), .c(s_101_39), .d(s_101_38), .cin(s_101_37), .o(t_2031), .co(t_2032), .cout(t_2033));
compressor_4_2 u2_700(.a(s_101_46), .b(s_101_45), .c(s_101_44), .d(s_101_43), .cin(s_101_42), .o(t_2034), .co(t_2035), .cout(t_2036));
compressor_3_2 u1_701(.a(s_101_49), .b(s_101_48), .cin(s_101_47), .o(t_2037), .cout(t_2038));
compressor_4_2 u2_702(.a(s_102_2), .b(s_102_1), .c(s_102_0), .d(t_2003), .cin(t_2006), .o(t_2039), .co(t_2040), .cout(t_2041));
compressor_4_2 u2_703(.a(s_102_5), .b(s_102_4), .c(s_102_3), .d(t_2009), .cin(t_2012), .o(t_2042), .co(t_2043), .cout(t_2044));
compressor_4_2 u2_704(.a(s_102_8), .b(s_102_7), .c(s_102_6), .d(t_2015), .cin(t_2018), .o(t_2045), .co(t_2046), .cout(t_2047));
compressor_4_2 u2_705(.a(s_102_11), .b(s_102_10), .c(s_102_9), .d(t_2021), .cin(t_2024), .o(t_2048), .co(t_2049), .cout(t_2050));
compressor_4_2 u2_706(.a(s_102_14), .b(s_102_13), .c(s_102_12), .d(t_2027), .cin(t_2030), .o(t_2051), .co(t_2052), .cout(t_2053));
compressor_4_2 u2_707(.a(s_102_17), .b(s_102_16), .c(s_102_15), .d(t_2033), .cin(t_2036), .o(t_2054), .co(t_2055), .cout(t_2056));
compressor_4_2 u2_708(.a(s_102_21), .b(s_102_20), .c(s_102_19), .d(s_102_18), .cin(t_2038), .o(t_2057), .co(t_2058), .cout(t_2059));
compressor_4_2 u2_709(.a(s_102_26), .b(s_102_25), .c(s_102_24), .d(s_102_23), .cin(s_102_22), .o(t_2060), .co(t_2061), .cout(t_2062));
compressor_4_2 u2_710(.a(s_102_31), .b(s_102_30), .c(s_102_29), .d(s_102_28), .cin(s_102_27), .o(t_2063), .co(t_2064), .cout(t_2065));
compressor_4_2 u2_711(.a(s_102_36), .b(s_102_35), .c(s_102_34), .d(s_102_33), .cin(s_102_32), .o(t_2066), .co(t_2067), .cout(t_2068));
compressor_4_2 u2_712(.a(s_102_41), .b(s_102_40), .c(s_102_39), .d(s_102_38), .cin(s_102_37), .o(t_2069), .co(t_2070), .cout(t_2071));
compressor_4_2 u2_713(.a(s_102_46), .b(s_102_45), .c(s_102_44), .d(s_102_43), .cin(s_102_42), .o(t_2072), .co(t_2073), .cout(t_2074));
compressor_4_2 u2_714(.a(s_102_51), .b(s_102_50), .c(s_102_49), .d(s_102_48), .cin(s_102_47), .o(t_2075), .co(t_2076), .cout(t_2077));
compressor_4_2 u2_715(.a(s_103_2), .b(s_103_1), .c(s_103_0), .d(t_2041), .cin(t_2044), .o(t_2078), .co(t_2079), .cout(t_2080));
compressor_4_2 u2_716(.a(s_103_5), .b(s_103_4), .c(s_103_3), .d(t_2047), .cin(t_2050), .o(t_2081), .co(t_2082), .cout(t_2083));
compressor_4_2 u2_717(.a(s_103_8), .b(s_103_7), .c(s_103_6), .d(t_2053), .cin(t_2056), .o(t_2084), .co(t_2085), .cout(t_2086));
compressor_4_2 u2_718(.a(s_103_11), .b(s_103_10), .c(s_103_9), .d(t_2059), .cin(t_2062), .o(t_2087), .co(t_2088), .cout(t_2089));
compressor_4_2 u2_719(.a(s_103_14), .b(s_103_13), .c(s_103_12), .d(t_2065), .cin(t_2068), .o(t_2090), .co(t_2091), .cout(t_2092));
compressor_4_2 u2_720(.a(s_103_17), .b(s_103_16), .c(s_103_15), .d(t_2071), .cin(t_2074), .o(t_2093), .co(t_2094), .cout(t_2095));
compressor_4_2 u2_721(.a(s_103_21), .b(s_103_20), .c(s_103_19), .d(s_103_18), .cin(t_2077), .o(t_2096), .co(t_2097), .cout(t_2098));
compressor_4_2 u2_722(.a(s_103_26), .b(s_103_25), .c(s_103_24), .d(s_103_23), .cin(s_103_22), .o(t_2099), .co(t_2100), .cout(t_2101));
compressor_4_2 u2_723(.a(s_103_31), .b(s_103_30), .c(s_103_29), .d(s_103_28), .cin(s_103_27), .o(t_2102), .co(t_2103), .cout(t_2104));
compressor_4_2 u2_724(.a(s_103_36), .b(s_103_35), .c(s_103_34), .d(s_103_33), .cin(s_103_32), .o(t_2105), .co(t_2106), .cout(t_2107));
compressor_4_2 u2_725(.a(s_103_41), .b(s_103_40), .c(s_103_39), .d(s_103_38), .cin(s_103_37), .o(t_2108), .co(t_2109), .cout(t_2110));
compressor_4_2 u2_726(.a(s_103_46), .b(s_103_45), .c(s_103_44), .d(s_103_43), .cin(s_103_42), .o(t_2111), .co(t_2112), .cout(t_2113));
compressor_4_2 u2_727(.a(s_103_51), .b(s_103_50), .c(s_103_49), .d(s_103_48), .cin(s_103_47), .o(t_2114), .co(t_2115), .cout(t_2116));
compressor_4_2 u2_728(.a(s_104_2), .b(s_104_1), .c(s_104_0), .d(t_2080), .cin(t_2083), .o(t_2117), .co(t_2118), .cout(t_2119));
compressor_4_2 u2_729(.a(s_104_5), .b(s_104_4), .c(s_104_3), .d(t_2086), .cin(t_2089), .o(t_2120), .co(t_2121), .cout(t_2122));
compressor_4_2 u2_730(.a(s_104_8), .b(s_104_7), .c(s_104_6), .d(t_2092), .cin(t_2095), .o(t_2123), .co(t_2124), .cout(t_2125));
compressor_4_2 u2_731(.a(s_104_11), .b(s_104_10), .c(s_104_9), .d(t_2098), .cin(t_2101), .o(t_2126), .co(t_2127), .cout(t_2128));
compressor_4_2 u2_732(.a(s_104_14), .b(s_104_13), .c(s_104_12), .d(t_2104), .cin(t_2107), .o(t_2129), .co(t_2130), .cout(t_2131));
compressor_4_2 u2_733(.a(s_104_17), .b(s_104_16), .c(s_104_15), .d(t_2110), .cin(t_2113), .o(t_2132), .co(t_2133), .cout(t_2134));
compressor_4_2 u2_734(.a(s_104_21), .b(s_104_20), .c(s_104_19), .d(s_104_18), .cin(t_2116), .o(t_2135), .co(t_2136), .cout(t_2137));
compressor_4_2 u2_735(.a(s_104_26), .b(s_104_25), .c(s_104_24), .d(s_104_23), .cin(s_104_22), .o(t_2138), .co(t_2139), .cout(t_2140));
compressor_4_2 u2_736(.a(s_104_31), .b(s_104_30), .c(s_104_29), .d(s_104_28), .cin(s_104_27), .o(t_2141), .co(t_2142), .cout(t_2143));
compressor_4_2 u2_737(.a(s_104_36), .b(s_104_35), .c(s_104_34), .d(s_104_33), .cin(s_104_32), .o(t_2144), .co(t_2145), .cout(t_2146));
compressor_4_2 u2_738(.a(s_104_41), .b(s_104_40), .c(s_104_39), .d(s_104_38), .cin(s_104_37), .o(t_2147), .co(t_2148), .cout(t_2149));
compressor_4_2 u2_739(.a(s_104_46), .b(s_104_45), .c(s_104_44), .d(s_104_43), .cin(s_104_42), .o(t_2150), .co(t_2151), .cout(t_2152));
compressor_4_2 u2_740(.a(s_104_51), .b(s_104_50), .c(s_104_49), .d(s_104_48), .cin(s_104_47), .o(t_2153), .co(t_2154), .cout(t_2155));
half_adder u0_741(.a(s_104_53), .b(s_104_52), .o(t_2156), .cout(t_2157));
compressor_4_2 u2_742(.a(s_105_2), .b(s_105_1), .c(s_105_0), .d(t_2119), .cin(t_2122), .o(t_2158), .co(t_2159), .cout(t_2160));
compressor_4_2 u2_743(.a(s_105_5), .b(s_105_4), .c(s_105_3), .d(t_2125), .cin(t_2128), .o(t_2161), .co(t_2162), .cout(t_2163));
compressor_4_2 u2_744(.a(s_105_8), .b(s_105_7), .c(s_105_6), .d(t_2131), .cin(t_2134), .o(t_2164), .co(t_2165), .cout(t_2166));
compressor_4_2 u2_745(.a(s_105_11), .b(s_105_10), .c(s_105_9), .d(t_2137), .cin(t_2140), .o(t_2167), .co(t_2168), .cout(t_2169));
compressor_4_2 u2_746(.a(s_105_14), .b(s_105_13), .c(s_105_12), .d(t_2143), .cin(t_2146), .o(t_2170), .co(t_2171), .cout(t_2172));
compressor_4_2 u2_747(.a(s_105_17), .b(s_105_16), .c(s_105_15), .d(t_2149), .cin(t_2152), .o(t_2173), .co(t_2174), .cout(t_2175));
compressor_4_2 u2_748(.a(s_105_20), .b(s_105_19), .c(s_105_18), .d(t_2155), .cin(t_2157), .o(t_2176), .co(t_2177), .cout(t_2178));
compressor_4_2 u2_749(.a(s_105_25), .b(s_105_24), .c(s_105_23), .d(s_105_22), .cin(s_105_21), .o(t_2179), .co(t_2180), .cout(t_2181));
compressor_4_2 u2_750(.a(s_105_30), .b(s_105_29), .c(s_105_28), .d(s_105_27), .cin(s_105_26), .o(t_2182), .co(t_2183), .cout(t_2184));
compressor_4_2 u2_751(.a(s_105_35), .b(s_105_34), .c(s_105_33), .d(s_105_32), .cin(s_105_31), .o(t_2185), .co(t_2186), .cout(t_2187));
compressor_4_2 u2_752(.a(s_105_40), .b(s_105_39), .c(s_105_38), .d(s_105_37), .cin(s_105_36), .o(t_2188), .co(t_2189), .cout(t_2190));
compressor_4_2 u2_753(.a(s_105_45), .b(s_105_44), .c(s_105_43), .d(s_105_42), .cin(s_105_41), .o(t_2191), .co(t_2192), .cout(t_2193));
compressor_4_2 u2_754(.a(s_105_50), .b(s_105_49), .c(s_105_48), .d(s_105_47), .cin(s_105_46), .o(t_2194), .co(t_2195), .cout(t_2196));
half_adder u0_755(.a(s_105_52), .b(s_105_51), .o(t_2197), .cout(t_2198));
compressor_4_2 u2_756(.a(s_106_2), .b(s_106_1), .c(s_106_0), .d(t_2160), .cin(t_2163), .o(t_2199), .co(t_2200), .cout(t_2201));
compressor_4_2 u2_757(.a(s_106_5), .b(s_106_4), .c(s_106_3), .d(t_2166), .cin(t_2169), .o(t_2202), .co(t_2203), .cout(t_2204));
compressor_4_2 u2_758(.a(s_106_8), .b(s_106_7), .c(s_106_6), .d(t_2172), .cin(t_2175), .o(t_2205), .co(t_2206), .cout(t_2207));
compressor_4_2 u2_759(.a(s_106_11), .b(s_106_10), .c(s_106_9), .d(t_2178), .cin(t_2181), .o(t_2208), .co(t_2209), .cout(t_2210));
compressor_4_2 u2_760(.a(s_106_14), .b(s_106_13), .c(s_106_12), .d(t_2184), .cin(t_2187), .o(t_2211), .co(t_2212), .cout(t_2213));
compressor_4_2 u2_761(.a(s_106_17), .b(s_106_16), .c(s_106_15), .d(t_2190), .cin(t_2193), .o(t_2214), .co(t_2215), .cout(t_2216));
compressor_4_2 u2_762(.a(s_106_20), .b(s_106_19), .c(s_106_18), .d(t_2196), .cin(t_2198), .o(t_2217), .co(t_2218), .cout(t_2219));
compressor_4_2 u2_763(.a(s_106_25), .b(s_106_24), .c(s_106_23), .d(s_106_22), .cin(s_106_21), .o(t_2220), .co(t_2221), .cout(t_2222));
compressor_4_2 u2_764(.a(s_106_30), .b(s_106_29), .c(s_106_28), .d(s_106_27), .cin(s_106_26), .o(t_2223), .co(t_2224), .cout(t_2225));
compressor_4_2 u2_765(.a(s_106_35), .b(s_106_34), .c(s_106_33), .d(s_106_32), .cin(s_106_31), .o(t_2226), .co(t_2227), .cout(t_2228));
compressor_4_2 u2_766(.a(s_106_40), .b(s_106_39), .c(s_106_38), .d(s_106_37), .cin(s_106_36), .o(t_2229), .co(t_2230), .cout(t_2231));
compressor_4_2 u2_767(.a(s_106_45), .b(s_106_44), .c(s_106_43), .d(s_106_42), .cin(s_106_41), .o(t_2232), .co(t_2233), .cout(t_2234));
compressor_4_2 u2_768(.a(s_106_50), .b(s_106_49), .c(s_106_48), .d(s_106_47), .cin(s_106_46), .o(t_2235), .co(t_2236), .cout(t_2237));
compressor_3_2 u1_769(.a(s_106_53), .b(s_106_52), .cin(s_106_51), .o(t_2238), .cout(t_2239));
compressor_4_2 u2_770(.a(s_107_2), .b(s_107_1), .c(s_107_0), .d(t_2201), .cin(t_2204), .o(t_2240), .co(t_2241), .cout(t_2242));
compressor_4_2 u2_771(.a(s_107_5), .b(s_107_4), .c(s_107_3), .d(t_2207), .cin(t_2210), .o(t_2243), .co(t_2244), .cout(t_2245));
compressor_4_2 u2_772(.a(s_107_8), .b(s_107_7), .c(s_107_6), .d(t_2213), .cin(t_2216), .o(t_2246), .co(t_2247), .cout(t_2248));
compressor_4_2 u2_773(.a(s_107_11), .b(s_107_10), .c(s_107_9), .d(t_2219), .cin(t_2222), .o(t_2249), .co(t_2250), .cout(t_2251));
compressor_4_2 u2_774(.a(s_107_14), .b(s_107_13), .c(s_107_12), .d(t_2225), .cin(t_2228), .o(t_2252), .co(t_2253), .cout(t_2254));
compressor_4_2 u2_775(.a(s_107_17), .b(s_107_16), .c(s_107_15), .d(t_2231), .cin(t_2234), .o(t_2255), .co(t_2256), .cout(t_2257));
compressor_4_2 u2_776(.a(s_107_20), .b(s_107_19), .c(s_107_18), .d(t_2237), .cin(t_2239), .o(t_2258), .co(t_2259), .cout(t_2260));
compressor_4_2 u2_777(.a(s_107_25), .b(s_107_24), .c(s_107_23), .d(s_107_22), .cin(s_107_21), .o(t_2261), .co(t_2262), .cout(t_2263));
compressor_4_2 u2_778(.a(s_107_30), .b(s_107_29), .c(s_107_28), .d(s_107_27), .cin(s_107_26), .o(t_2264), .co(t_2265), .cout(t_2266));
compressor_4_2 u2_779(.a(s_107_35), .b(s_107_34), .c(s_107_33), .d(s_107_32), .cin(s_107_31), .o(t_2267), .co(t_2268), .cout(t_2269));
compressor_4_2 u2_780(.a(s_107_40), .b(s_107_39), .c(s_107_38), .d(s_107_37), .cin(s_107_36), .o(t_2270), .co(t_2271), .cout(t_2272));
compressor_4_2 u2_781(.a(s_107_45), .b(s_107_44), .c(s_107_43), .d(s_107_42), .cin(s_107_41), .o(t_2273), .co(t_2274), .cout(t_2275));
compressor_4_2 u2_782(.a(s_107_50), .b(s_107_49), .c(s_107_48), .d(s_107_47), .cin(s_107_46), .o(t_2276), .co(t_2277), .cout(t_2278));
compressor_3_2 u1_783(.a(s_107_53), .b(s_107_52), .cin(s_107_51), .o(t_2279), .cout(t_2280));
compressor_4_2 u2_784(.a(s_108_2), .b(s_108_1), .c(s_108_0), .d(t_2242), .cin(t_2245), .o(t_2281), .co(t_2282), .cout(t_2283));
compressor_4_2 u2_785(.a(s_108_5), .b(s_108_4), .c(s_108_3), .d(t_2248), .cin(t_2251), .o(t_2284), .co(t_2285), .cout(t_2286));
compressor_4_2 u2_786(.a(s_108_8), .b(s_108_7), .c(s_108_6), .d(t_2254), .cin(t_2257), .o(t_2287), .co(t_2288), .cout(t_2289));
compressor_4_2 u2_787(.a(s_108_11), .b(s_108_10), .c(s_108_9), .d(t_2260), .cin(t_2263), .o(t_2290), .co(t_2291), .cout(t_2292));
compressor_4_2 u2_788(.a(s_108_14), .b(s_108_13), .c(s_108_12), .d(t_2266), .cin(t_2269), .o(t_2293), .co(t_2294), .cout(t_2295));
compressor_4_2 u2_789(.a(s_108_17), .b(s_108_16), .c(s_108_15), .d(t_2272), .cin(t_2275), .o(t_2296), .co(t_2297), .cout(t_2298));
compressor_4_2 u2_790(.a(s_108_20), .b(s_108_19), .c(s_108_18), .d(t_2278), .cin(t_2280), .o(t_2299), .co(t_2300), .cout(t_2301));
compressor_4_2 u2_791(.a(s_108_25), .b(s_108_24), .c(s_108_23), .d(s_108_22), .cin(s_108_21), .o(t_2302), .co(t_2303), .cout(t_2304));
compressor_4_2 u2_792(.a(s_108_30), .b(s_108_29), .c(s_108_28), .d(s_108_27), .cin(s_108_26), .o(t_2305), .co(t_2306), .cout(t_2307));
compressor_4_2 u2_793(.a(s_108_35), .b(s_108_34), .c(s_108_33), .d(s_108_32), .cin(s_108_31), .o(t_2308), .co(t_2309), .cout(t_2310));
compressor_4_2 u2_794(.a(s_108_40), .b(s_108_39), .c(s_108_38), .d(s_108_37), .cin(s_108_36), .o(t_2311), .co(t_2312), .cout(t_2313));
compressor_4_2 u2_795(.a(s_108_45), .b(s_108_44), .c(s_108_43), .d(s_108_42), .cin(s_108_41), .o(t_2314), .co(t_2315), .cout(t_2316));
compressor_4_2 u2_796(.a(s_108_50), .b(s_108_49), .c(s_108_48), .d(s_108_47), .cin(s_108_46), .o(t_2317), .co(t_2318), .cout(t_2319));
compressor_4_2 u2_797(.a(s_108_55), .b(s_108_54), .c(s_108_53), .d(s_108_52), .cin(s_108_51), .o(t_2320), .co(t_2321), .cout(t_2322));
compressor_4_2 u2_798(.a(s_109_2), .b(s_109_1), .c(s_109_0), .d(t_2283), .cin(t_2286), .o(t_2323), .co(t_2324), .cout(t_2325));
compressor_4_2 u2_799(.a(s_109_5), .b(s_109_4), .c(s_109_3), .d(t_2289), .cin(t_2292), .o(t_2326), .co(t_2327), .cout(t_2328));
compressor_4_2 u2_800(.a(s_109_8), .b(s_109_7), .c(s_109_6), .d(t_2295), .cin(t_2298), .o(t_2329), .co(t_2330), .cout(t_2331));
compressor_4_2 u2_801(.a(s_109_11), .b(s_109_10), .c(s_109_9), .d(t_2301), .cin(t_2304), .o(t_2332), .co(t_2333), .cout(t_2334));
compressor_4_2 u2_802(.a(s_109_14), .b(s_109_13), .c(s_109_12), .d(t_2307), .cin(t_2310), .o(t_2335), .co(t_2336), .cout(t_2337));
compressor_4_2 u2_803(.a(s_109_17), .b(s_109_16), .c(s_109_15), .d(t_2313), .cin(t_2316), .o(t_2338), .co(t_2339), .cout(t_2340));
compressor_4_2 u2_804(.a(s_109_20), .b(s_109_19), .c(s_109_18), .d(t_2319), .cin(t_2322), .o(t_2341), .co(t_2342), .cout(t_2343));
compressor_4_2 u2_805(.a(s_109_25), .b(s_109_24), .c(s_109_23), .d(s_109_22), .cin(s_109_21), .o(t_2344), .co(t_2345), .cout(t_2346));
compressor_4_2 u2_806(.a(s_109_30), .b(s_109_29), .c(s_109_28), .d(s_109_27), .cin(s_109_26), .o(t_2347), .co(t_2348), .cout(t_2349));
compressor_4_2 u2_807(.a(s_109_35), .b(s_109_34), .c(s_109_33), .d(s_109_32), .cin(s_109_31), .o(t_2350), .co(t_2351), .cout(t_2352));
compressor_4_2 u2_808(.a(s_109_40), .b(s_109_39), .c(s_109_38), .d(s_109_37), .cin(s_109_36), .o(t_2353), .co(t_2354), .cout(t_2355));
compressor_4_2 u2_809(.a(s_109_45), .b(s_109_44), .c(s_109_43), .d(s_109_42), .cin(s_109_41), .o(t_2356), .co(t_2357), .cout(t_2358));
compressor_4_2 u2_810(.a(s_109_50), .b(s_109_49), .c(s_109_48), .d(s_109_47), .cin(s_109_46), .o(t_2359), .co(t_2360), .cout(t_2361));
compressor_3_2 u1_811(.a(s_109_53), .b(s_109_52), .cin(s_109_51), .o(t_2362), .cout(t_2363));
compressor_4_2 u2_812(.a(s_110_2), .b(s_110_1), .c(s_110_0), .d(t_2325), .cin(t_2328), .o(t_2364), .co(t_2365), .cout(t_2366));
compressor_4_2 u2_813(.a(s_110_5), .b(s_110_4), .c(s_110_3), .d(t_2331), .cin(t_2334), .o(t_2367), .co(t_2368), .cout(t_2369));
compressor_4_2 u2_814(.a(s_110_8), .b(s_110_7), .c(s_110_6), .d(t_2337), .cin(t_2340), .o(t_2370), .co(t_2371), .cout(t_2372));
compressor_4_2 u2_815(.a(s_110_11), .b(s_110_10), .c(s_110_9), .d(t_2343), .cin(t_2346), .o(t_2373), .co(t_2374), .cout(t_2375));
compressor_4_2 u2_816(.a(s_110_14), .b(s_110_13), .c(s_110_12), .d(t_2349), .cin(t_2352), .o(t_2376), .co(t_2377), .cout(t_2378));
compressor_4_2 u2_817(.a(s_110_17), .b(s_110_16), .c(s_110_15), .d(t_2355), .cin(t_2358), .o(t_2379), .co(t_2380), .cout(t_2381));
compressor_4_2 u2_818(.a(s_110_20), .b(s_110_19), .c(s_110_18), .d(t_2361), .cin(t_2363), .o(t_2382), .co(t_2383), .cout(t_2384));
compressor_4_2 u2_819(.a(s_110_25), .b(s_110_24), .c(s_110_23), .d(s_110_22), .cin(s_110_21), .o(t_2385), .co(t_2386), .cout(t_2387));
compressor_4_2 u2_820(.a(s_110_30), .b(s_110_29), .c(s_110_28), .d(s_110_27), .cin(s_110_26), .o(t_2388), .co(t_2389), .cout(t_2390));
compressor_4_2 u2_821(.a(s_110_35), .b(s_110_34), .c(s_110_33), .d(s_110_32), .cin(s_110_31), .o(t_2391), .co(t_2392), .cout(t_2393));
compressor_4_2 u2_822(.a(s_110_40), .b(s_110_39), .c(s_110_38), .d(s_110_37), .cin(s_110_36), .o(t_2394), .co(t_2395), .cout(t_2396));
compressor_4_2 u2_823(.a(s_110_45), .b(s_110_44), .c(s_110_43), .d(s_110_42), .cin(s_110_41), .o(t_2397), .co(t_2398), .cout(t_2399));
compressor_4_2 u2_824(.a(s_110_50), .b(s_110_49), .c(s_110_48), .d(s_110_47), .cin(s_110_46), .o(t_2400), .co(t_2401), .cout(t_2402));
compressor_4_2 u2_825(.a(s_110_55), .b(s_110_54), .c(s_110_53), .d(s_110_52), .cin(s_110_51), .o(t_2403), .co(t_2404), .cout(t_2405));
compressor_4_2 u2_826(.a(s_111_2), .b(s_111_1), .c(s_111_0), .d(t_2366), .cin(t_2369), .o(t_2406), .co(t_2407), .cout(t_2408));
compressor_4_2 u2_827(.a(s_111_5), .b(s_111_4), .c(s_111_3), .d(t_2372), .cin(t_2375), .o(t_2409), .co(t_2410), .cout(t_2411));
compressor_4_2 u2_828(.a(s_111_8), .b(s_111_7), .c(s_111_6), .d(t_2378), .cin(t_2381), .o(t_2412), .co(t_2413), .cout(t_2414));
compressor_4_2 u2_829(.a(s_111_11), .b(s_111_10), .c(s_111_9), .d(t_2384), .cin(t_2387), .o(t_2415), .co(t_2416), .cout(t_2417));
compressor_4_2 u2_830(.a(s_111_14), .b(s_111_13), .c(s_111_12), .d(t_2390), .cin(t_2393), .o(t_2418), .co(t_2419), .cout(t_2420));
compressor_4_2 u2_831(.a(s_111_17), .b(s_111_16), .c(s_111_15), .d(t_2396), .cin(t_2399), .o(t_2421), .co(t_2422), .cout(t_2423));
compressor_4_2 u2_832(.a(s_111_20), .b(s_111_19), .c(s_111_18), .d(t_2402), .cin(t_2405), .o(t_2424), .co(t_2425), .cout(t_2426));
compressor_4_2 u2_833(.a(s_111_25), .b(s_111_24), .c(s_111_23), .d(s_111_22), .cin(s_111_21), .o(t_2427), .co(t_2428), .cout(t_2429));
compressor_4_2 u2_834(.a(s_111_30), .b(s_111_29), .c(s_111_28), .d(s_111_27), .cin(s_111_26), .o(t_2430), .co(t_2431), .cout(t_2432));
compressor_4_2 u2_835(.a(s_111_35), .b(s_111_34), .c(s_111_33), .d(s_111_32), .cin(s_111_31), .o(t_2433), .co(t_2434), .cout(t_2435));
compressor_4_2 u2_836(.a(s_111_40), .b(s_111_39), .c(s_111_38), .d(s_111_37), .cin(s_111_36), .o(t_2436), .co(t_2437), .cout(t_2438));
compressor_4_2 u2_837(.a(s_111_45), .b(s_111_44), .c(s_111_43), .d(s_111_42), .cin(s_111_41), .o(t_2439), .co(t_2440), .cout(t_2441));
compressor_4_2 u2_838(.a(s_111_50), .b(s_111_49), .c(s_111_48), .d(s_111_47), .cin(s_111_46), .o(t_2442), .co(t_2443), .cout(t_2444));
compressor_4_2 u2_839(.a(s_111_55), .b(s_111_54), .c(s_111_53), .d(s_111_52), .cin(s_111_51), .o(t_2445), .co(t_2446), .cout(t_2447));
compressor_4_2 u2_840(.a(s_112_2), .b(s_112_1), .c(s_112_0), .d(t_2408), .cin(t_2411), .o(t_2448), .co(t_2449), .cout(t_2450));
compressor_4_2 u2_841(.a(s_112_5), .b(s_112_4), .c(s_112_3), .d(t_2414), .cin(t_2417), .o(t_2451), .co(t_2452), .cout(t_2453));
compressor_4_2 u2_842(.a(s_112_8), .b(s_112_7), .c(s_112_6), .d(t_2420), .cin(t_2423), .o(t_2454), .co(t_2455), .cout(t_2456));
compressor_4_2 u2_843(.a(s_112_11), .b(s_112_10), .c(s_112_9), .d(t_2426), .cin(t_2429), .o(t_2457), .co(t_2458), .cout(t_2459));
compressor_4_2 u2_844(.a(s_112_14), .b(s_112_13), .c(s_112_12), .d(t_2432), .cin(t_2435), .o(t_2460), .co(t_2461), .cout(t_2462));
compressor_4_2 u2_845(.a(s_112_17), .b(s_112_16), .c(s_112_15), .d(t_2438), .cin(t_2441), .o(t_2463), .co(t_2464), .cout(t_2465));
compressor_4_2 u2_846(.a(s_112_20), .b(s_112_19), .c(s_112_18), .d(t_2444), .cin(t_2447), .o(t_2466), .co(t_2467), .cout(t_2468));
compressor_4_2 u2_847(.a(s_112_25), .b(s_112_24), .c(s_112_23), .d(s_112_22), .cin(s_112_21), .o(t_2469), .co(t_2470), .cout(t_2471));
compressor_4_2 u2_848(.a(s_112_30), .b(s_112_29), .c(s_112_28), .d(s_112_27), .cin(s_112_26), .o(t_2472), .co(t_2473), .cout(t_2474));
compressor_4_2 u2_849(.a(s_112_35), .b(s_112_34), .c(s_112_33), .d(s_112_32), .cin(s_112_31), .o(t_2475), .co(t_2476), .cout(t_2477));
compressor_4_2 u2_850(.a(s_112_40), .b(s_112_39), .c(s_112_38), .d(s_112_37), .cin(s_112_36), .o(t_2478), .co(t_2479), .cout(t_2480));
compressor_4_2 u2_851(.a(s_112_45), .b(s_112_44), .c(s_112_43), .d(s_112_42), .cin(s_112_41), .o(t_2481), .co(t_2482), .cout(t_2483));
compressor_4_2 u2_852(.a(s_112_50), .b(s_112_49), .c(s_112_48), .d(s_112_47), .cin(s_112_46), .o(t_2484), .co(t_2485), .cout(t_2486));
compressor_4_2 u2_853(.a(s_112_55), .b(s_112_54), .c(s_112_53), .d(s_112_52), .cin(s_112_51), .o(t_2487), .co(t_2488), .cout(t_2489));
half_adder u0_854(.a(s_112_57), .b(s_112_56), .o(t_2490), .cout(t_2491));
compressor_4_2 u2_855(.a(s_113_2), .b(s_113_1), .c(s_113_0), .d(t_2450), .cin(t_2453), .o(t_2492), .co(t_2493), .cout(t_2494));
compressor_4_2 u2_856(.a(s_113_5), .b(s_113_4), .c(s_113_3), .d(t_2456), .cin(t_2459), .o(t_2495), .co(t_2496), .cout(t_2497));
compressor_4_2 u2_857(.a(s_113_8), .b(s_113_7), .c(s_113_6), .d(t_2462), .cin(t_2465), .o(t_2498), .co(t_2499), .cout(t_2500));
compressor_4_2 u2_858(.a(s_113_11), .b(s_113_10), .c(s_113_9), .d(t_2468), .cin(t_2471), .o(t_2501), .co(t_2502), .cout(t_2503));
compressor_4_2 u2_859(.a(s_113_14), .b(s_113_13), .c(s_113_12), .d(t_2474), .cin(t_2477), .o(t_2504), .co(t_2505), .cout(t_2506));
compressor_4_2 u2_860(.a(s_113_17), .b(s_113_16), .c(s_113_15), .d(t_2480), .cin(t_2483), .o(t_2507), .co(t_2508), .cout(t_2509));
compressor_4_2 u2_861(.a(s_113_20), .b(s_113_19), .c(s_113_18), .d(t_2486), .cin(t_2489), .o(t_2510), .co(t_2511), .cout(t_2512));
compressor_4_2 u2_862(.a(s_113_24), .b(s_113_23), .c(s_113_22), .d(s_113_21), .cin(t_2491), .o(t_2513), .co(t_2514), .cout(t_2515));
compressor_4_2 u2_863(.a(s_113_29), .b(s_113_28), .c(s_113_27), .d(s_113_26), .cin(s_113_25), .o(t_2516), .co(t_2517), .cout(t_2518));
compressor_4_2 u2_864(.a(s_113_34), .b(s_113_33), .c(s_113_32), .d(s_113_31), .cin(s_113_30), .o(t_2519), .co(t_2520), .cout(t_2521));
compressor_4_2 u2_865(.a(s_113_39), .b(s_113_38), .c(s_113_37), .d(s_113_36), .cin(s_113_35), .o(t_2522), .co(t_2523), .cout(t_2524));
compressor_4_2 u2_866(.a(s_113_44), .b(s_113_43), .c(s_113_42), .d(s_113_41), .cin(s_113_40), .o(t_2525), .co(t_2526), .cout(t_2527));
compressor_4_2 u2_867(.a(s_113_49), .b(s_113_48), .c(s_113_47), .d(s_113_46), .cin(s_113_45), .o(t_2528), .co(t_2529), .cout(t_2530));
compressor_4_2 u2_868(.a(s_113_54), .b(s_113_53), .c(s_113_52), .d(s_113_51), .cin(s_113_50), .o(t_2531), .co(t_2532), .cout(t_2533));
half_adder u0_869(.a(s_113_56), .b(s_113_55), .o(t_2534), .cout(t_2535));
compressor_4_2 u2_870(.a(s_114_2), .b(s_114_1), .c(s_114_0), .d(t_2494), .cin(t_2497), .o(t_2536), .co(t_2537), .cout(t_2538));
compressor_4_2 u2_871(.a(s_114_5), .b(s_114_4), .c(s_114_3), .d(t_2500), .cin(t_2503), .o(t_2539), .co(t_2540), .cout(t_2541));
compressor_4_2 u2_872(.a(s_114_8), .b(s_114_7), .c(s_114_6), .d(t_2506), .cin(t_2509), .o(t_2542), .co(t_2543), .cout(t_2544));
compressor_4_2 u2_873(.a(s_114_11), .b(s_114_10), .c(s_114_9), .d(t_2512), .cin(t_2515), .o(t_2545), .co(t_2546), .cout(t_2547));
compressor_4_2 u2_874(.a(s_114_14), .b(s_114_13), .c(s_114_12), .d(t_2518), .cin(t_2521), .o(t_2548), .co(t_2549), .cout(t_2550));
compressor_4_2 u2_875(.a(s_114_17), .b(s_114_16), .c(s_114_15), .d(t_2524), .cin(t_2527), .o(t_2551), .co(t_2552), .cout(t_2553));
compressor_4_2 u2_876(.a(s_114_20), .b(s_114_19), .c(s_114_18), .d(t_2530), .cin(t_2533), .o(t_2554), .co(t_2555), .cout(t_2556));
compressor_4_2 u2_877(.a(s_114_24), .b(s_114_23), .c(s_114_22), .d(s_114_21), .cin(t_2535), .o(t_2557), .co(t_2558), .cout(t_2559));
compressor_4_2 u2_878(.a(s_114_29), .b(s_114_28), .c(s_114_27), .d(s_114_26), .cin(s_114_25), .o(t_2560), .co(t_2561), .cout(t_2562));
compressor_4_2 u2_879(.a(s_114_34), .b(s_114_33), .c(s_114_32), .d(s_114_31), .cin(s_114_30), .o(t_2563), .co(t_2564), .cout(t_2565));
compressor_4_2 u2_880(.a(s_114_39), .b(s_114_38), .c(s_114_37), .d(s_114_36), .cin(s_114_35), .o(t_2566), .co(t_2567), .cout(t_2568));
compressor_4_2 u2_881(.a(s_114_44), .b(s_114_43), .c(s_114_42), .d(s_114_41), .cin(s_114_40), .o(t_2569), .co(t_2570), .cout(t_2571));
compressor_4_2 u2_882(.a(s_114_49), .b(s_114_48), .c(s_114_47), .d(s_114_46), .cin(s_114_45), .o(t_2572), .co(t_2573), .cout(t_2574));
compressor_4_2 u2_883(.a(s_114_54), .b(s_114_53), .c(s_114_52), .d(s_114_51), .cin(s_114_50), .o(t_2575), .co(t_2576), .cout(t_2577));
compressor_3_2 u1_884(.a(s_114_57), .b(s_114_56), .cin(s_114_55), .o(t_2578), .cout(t_2579));
compressor_4_2 u2_885(.a(s_115_2), .b(s_115_1), .c(s_115_0), .d(t_2538), .cin(t_2541), .o(t_2580), .co(t_2581), .cout(t_2582));
compressor_4_2 u2_886(.a(s_115_5), .b(s_115_4), .c(s_115_3), .d(t_2544), .cin(t_2547), .o(t_2583), .co(t_2584), .cout(t_2585));
compressor_4_2 u2_887(.a(s_115_8), .b(s_115_7), .c(s_115_6), .d(t_2550), .cin(t_2553), .o(t_2586), .co(t_2587), .cout(t_2588));
compressor_4_2 u2_888(.a(s_115_11), .b(s_115_10), .c(s_115_9), .d(t_2556), .cin(t_2559), .o(t_2589), .co(t_2590), .cout(t_2591));
compressor_4_2 u2_889(.a(s_115_14), .b(s_115_13), .c(s_115_12), .d(t_2562), .cin(t_2565), .o(t_2592), .co(t_2593), .cout(t_2594));
compressor_4_2 u2_890(.a(s_115_17), .b(s_115_16), .c(s_115_15), .d(t_2568), .cin(t_2571), .o(t_2595), .co(t_2596), .cout(t_2597));
compressor_4_2 u2_891(.a(s_115_20), .b(s_115_19), .c(s_115_18), .d(t_2574), .cin(t_2577), .o(t_2598), .co(t_2599), .cout(t_2600));
compressor_4_2 u2_892(.a(s_115_24), .b(s_115_23), .c(s_115_22), .d(s_115_21), .cin(t_2579), .o(t_2601), .co(t_2602), .cout(t_2603));
compressor_4_2 u2_893(.a(s_115_29), .b(s_115_28), .c(s_115_27), .d(s_115_26), .cin(s_115_25), .o(t_2604), .co(t_2605), .cout(t_2606));
compressor_4_2 u2_894(.a(s_115_34), .b(s_115_33), .c(s_115_32), .d(s_115_31), .cin(s_115_30), .o(t_2607), .co(t_2608), .cout(t_2609));
compressor_4_2 u2_895(.a(s_115_39), .b(s_115_38), .c(s_115_37), .d(s_115_36), .cin(s_115_35), .o(t_2610), .co(t_2611), .cout(t_2612));
compressor_4_2 u2_896(.a(s_115_44), .b(s_115_43), .c(s_115_42), .d(s_115_41), .cin(s_115_40), .o(t_2613), .co(t_2614), .cout(t_2615));
compressor_4_2 u2_897(.a(s_115_49), .b(s_115_48), .c(s_115_47), .d(s_115_46), .cin(s_115_45), .o(t_2616), .co(t_2617), .cout(t_2618));
compressor_4_2 u2_898(.a(s_115_54), .b(s_115_53), .c(s_115_52), .d(s_115_51), .cin(s_115_50), .o(t_2619), .co(t_2620), .cout(t_2621));
compressor_3_2 u1_899(.a(s_115_57), .b(s_115_56), .cin(s_115_55), .o(t_2622), .cout(t_2623));
compressor_4_2 u2_900(.a(s_116_2), .b(s_116_1), .c(s_116_0), .d(t_2582), .cin(t_2585), .o(t_2624), .co(t_2625), .cout(t_2626));
compressor_4_2 u2_901(.a(s_116_5), .b(s_116_4), .c(s_116_3), .d(t_2588), .cin(t_2591), .o(t_2627), .co(t_2628), .cout(t_2629));
compressor_4_2 u2_902(.a(s_116_8), .b(s_116_7), .c(s_116_6), .d(t_2594), .cin(t_2597), .o(t_2630), .co(t_2631), .cout(t_2632));
compressor_4_2 u2_903(.a(s_116_11), .b(s_116_10), .c(s_116_9), .d(t_2600), .cin(t_2603), .o(t_2633), .co(t_2634), .cout(t_2635));
compressor_4_2 u2_904(.a(s_116_14), .b(s_116_13), .c(s_116_12), .d(t_2606), .cin(t_2609), .o(t_2636), .co(t_2637), .cout(t_2638));
compressor_4_2 u2_905(.a(s_116_17), .b(s_116_16), .c(s_116_15), .d(t_2612), .cin(t_2615), .o(t_2639), .co(t_2640), .cout(t_2641));
compressor_4_2 u2_906(.a(s_116_20), .b(s_116_19), .c(s_116_18), .d(t_2618), .cin(t_2621), .o(t_2642), .co(t_2643), .cout(t_2644));
compressor_4_2 u2_907(.a(s_116_24), .b(s_116_23), .c(s_116_22), .d(s_116_21), .cin(t_2623), .o(t_2645), .co(t_2646), .cout(t_2647));
compressor_4_2 u2_908(.a(s_116_29), .b(s_116_28), .c(s_116_27), .d(s_116_26), .cin(s_116_25), .o(t_2648), .co(t_2649), .cout(t_2650));
compressor_4_2 u2_909(.a(s_116_34), .b(s_116_33), .c(s_116_32), .d(s_116_31), .cin(s_116_30), .o(t_2651), .co(t_2652), .cout(t_2653));
compressor_4_2 u2_910(.a(s_116_39), .b(s_116_38), .c(s_116_37), .d(s_116_36), .cin(s_116_35), .o(t_2654), .co(t_2655), .cout(t_2656));
compressor_4_2 u2_911(.a(s_116_44), .b(s_116_43), .c(s_116_42), .d(s_116_41), .cin(s_116_40), .o(t_2657), .co(t_2658), .cout(t_2659));
compressor_4_2 u2_912(.a(s_116_49), .b(s_116_48), .c(s_116_47), .d(s_116_46), .cin(s_116_45), .o(t_2660), .co(t_2661), .cout(t_2662));
compressor_4_2 u2_913(.a(s_116_54), .b(s_116_53), .c(s_116_52), .d(s_116_51), .cin(s_116_50), .o(t_2663), .co(t_2664), .cout(t_2665));
compressor_4_2 u2_914(.a(s_116_59), .b(s_116_58), .c(s_116_57), .d(s_116_56), .cin(s_116_55), .o(t_2666), .co(t_2667), .cout(t_2668));
compressor_4_2 u2_915(.a(s_117_2), .b(s_117_1), .c(s_117_0), .d(t_2626), .cin(t_2629), .o(t_2669), .co(t_2670), .cout(t_2671));
compressor_4_2 u2_916(.a(s_117_5), .b(s_117_4), .c(s_117_3), .d(t_2632), .cin(t_2635), .o(t_2672), .co(t_2673), .cout(t_2674));
compressor_4_2 u2_917(.a(s_117_8), .b(s_117_7), .c(s_117_6), .d(t_2638), .cin(t_2641), .o(t_2675), .co(t_2676), .cout(t_2677));
compressor_4_2 u2_918(.a(s_117_11), .b(s_117_10), .c(s_117_9), .d(t_2644), .cin(t_2647), .o(t_2678), .co(t_2679), .cout(t_2680));
compressor_4_2 u2_919(.a(s_117_14), .b(s_117_13), .c(s_117_12), .d(t_2650), .cin(t_2653), .o(t_2681), .co(t_2682), .cout(t_2683));
compressor_4_2 u2_920(.a(s_117_17), .b(s_117_16), .c(s_117_15), .d(t_2656), .cin(t_2659), .o(t_2684), .co(t_2685), .cout(t_2686));
compressor_4_2 u2_921(.a(s_117_20), .b(s_117_19), .c(s_117_18), .d(t_2662), .cin(t_2665), .o(t_2687), .co(t_2688), .cout(t_2689));
compressor_4_2 u2_922(.a(s_117_24), .b(s_117_23), .c(s_117_22), .d(s_117_21), .cin(t_2668), .o(t_2690), .co(t_2691), .cout(t_2692));
compressor_4_2 u2_923(.a(s_117_29), .b(s_117_28), .c(s_117_27), .d(s_117_26), .cin(s_117_25), .o(t_2693), .co(t_2694), .cout(t_2695));
compressor_4_2 u2_924(.a(s_117_34), .b(s_117_33), .c(s_117_32), .d(s_117_31), .cin(s_117_30), .o(t_2696), .co(t_2697), .cout(t_2698));
compressor_4_2 u2_925(.a(s_117_39), .b(s_117_38), .c(s_117_37), .d(s_117_36), .cin(s_117_35), .o(t_2699), .co(t_2700), .cout(t_2701));
compressor_4_2 u2_926(.a(s_117_44), .b(s_117_43), .c(s_117_42), .d(s_117_41), .cin(s_117_40), .o(t_2702), .co(t_2703), .cout(t_2704));
compressor_4_2 u2_927(.a(s_117_49), .b(s_117_48), .c(s_117_47), .d(s_117_46), .cin(s_117_45), .o(t_2705), .co(t_2706), .cout(t_2707));
compressor_4_2 u2_928(.a(s_117_54), .b(s_117_53), .c(s_117_52), .d(s_117_51), .cin(s_117_50), .o(t_2708), .co(t_2709), .cout(t_2710));
compressor_3_2 u1_929(.a(s_117_57), .b(s_117_56), .cin(s_117_55), .o(t_2711), .cout(t_2712));
compressor_4_2 u2_930(.a(s_118_2), .b(s_118_1), .c(s_118_0), .d(t_2671), .cin(t_2674), .o(t_2713), .co(t_2714), .cout(t_2715));
compressor_4_2 u2_931(.a(s_118_5), .b(s_118_4), .c(s_118_3), .d(t_2677), .cin(t_2680), .o(t_2716), .co(t_2717), .cout(t_2718));
compressor_4_2 u2_932(.a(s_118_8), .b(s_118_7), .c(s_118_6), .d(t_2683), .cin(t_2686), .o(t_2719), .co(t_2720), .cout(t_2721));
compressor_4_2 u2_933(.a(s_118_11), .b(s_118_10), .c(s_118_9), .d(t_2689), .cin(t_2692), .o(t_2722), .co(t_2723), .cout(t_2724));
compressor_4_2 u2_934(.a(s_118_14), .b(s_118_13), .c(s_118_12), .d(t_2695), .cin(t_2698), .o(t_2725), .co(t_2726), .cout(t_2727));
compressor_4_2 u2_935(.a(s_118_17), .b(s_118_16), .c(s_118_15), .d(t_2701), .cin(t_2704), .o(t_2728), .co(t_2729), .cout(t_2730));
compressor_4_2 u2_936(.a(s_118_20), .b(s_118_19), .c(s_118_18), .d(t_2707), .cin(t_2710), .o(t_2731), .co(t_2732), .cout(t_2733));
compressor_4_2 u2_937(.a(s_118_24), .b(s_118_23), .c(s_118_22), .d(s_118_21), .cin(t_2712), .o(t_2734), .co(t_2735), .cout(t_2736));
compressor_4_2 u2_938(.a(s_118_29), .b(s_118_28), .c(s_118_27), .d(s_118_26), .cin(s_118_25), .o(t_2737), .co(t_2738), .cout(t_2739));
compressor_4_2 u2_939(.a(s_118_34), .b(s_118_33), .c(s_118_32), .d(s_118_31), .cin(s_118_30), .o(t_2740), .co(t_2741), .cout(t_2742));
compressor_4_2 u2_940(.a(s_118_39), .b(s_118_38), .c(s_118_37), .d(s_118_36), .cin(s_118_35), .o(t_2743), .co(t_2744), .cout(t_2745));
compressor_4_2 u2_941(.a(s_118_44), .b(s_118_43), .c(s_118_42), .d(s_118_41), .cin(s_118_40), .o(t_2746), .co(t_2747), .cout(t_2748));
compressor_4_2 u2_942(.a(s_118_49), .b(s_118_48), .c(s_118_47), .d(s_118_46), .cin(s_118_45), .o(t_2749), .co(t_2750), .cout(t_2751));
compressor_4_2 u2_943(.a(s_118_54), .b(s_118_53), .c(s_118_52), .d(s_118_51), .cin(s_118_50), .o(t_2752), .co(t_2753), .cout(t_2754));
compressor_4_2 u2_944(.a(s_118_59), .b(s_118_58), .c(s_118_57), .d(s_118_56), .cin(s_118_55), .o(t_2755), .co(t_2756), .cout(t_2757));
compressor_4_2 u2_945(.a(s_119_2), .b(s_119_1), .c(s_119_0), .d(t_2715), .cin(t_2718), .o(t_2758), .co(t_2759), .cout(t_2760));
compressor_4_2 u2_946(.a(s_119_5), .b(s_119_4), .c(s_119_3), .d(t_2721), .cin(t_2724), .o(t_2761), .co(t_2762), .cout(t_2763));
compressor_4_2 u2_947(.a(s_119_8), .b(s_119_7), .c(s_119_6), .d(t_2727), .cin(t_2730), .o(t_2764), .co(t_2765), .cout(t_2766));
compressor_4_2 u2_948(.a(s_119_11), .b(s_119_10), .c(s_119_9), .d(t_2733), .cin(t_2736), .o(t_2767), .co(t_2768), .cout(t_2769));
compressor_4_2 u2_949(.a(s_119_14), .b(s_119_13), .c(s_119_12), .d(t_2739), .cin(t_2742), .o(t_2770), .co(t_2771), .cout(t_2772));
compressor_4_2 u2_950(.a(s_119_17), .b(s_119_16), .c(s_119_15), .d(t_2745), .cin(t_2748), .o(t_2773), .co(t_2774), .cout(t_2775));
compressor_4_2 u2_951(.a(s_119_20), .b(s_119_19), .c(s_119_18), .d(t_2751), .cin(t_2754), .o(t_2776), .co(t_2777), .cout(t_2778));
compressor_4_2 u2_952(.a(s_119_24), .b(s_119_23), .c(s_119_22), .d(s_119_21), .cin(t_2757), .o(t_2779), .co(t_2780), .cout(t_2781));
compressor_4_2 u2_953(.a(s_119_29), .b(s_119_28), .c(s_119_27), .d(s_119_26), .cin(s_119_25), .o(t_2782), .co(t_2783), .cout(t_2784));
compressor_4_2 u2_954(.a(s_119_34), .b(s_119_33), .c(s_119_32), .d(s_119_31), .cin(s_119_30), .o(t_2785), .co(t_2786), .cout(t_2787));
compressor_4_2 u2_955(.a(s_119_39), .b(s_119_38), .c(s_119_37), .d(s_119_36), .cin(s_119_35), .o(t_2788), .co(t_2789), .cout(t_2790));
compressor_4_2 u2_956(.a(s_119_44), .b(s_119_43), .c(s_119_42), .d(s_119_41), .cin(s_119_40), .o(t_2791), .co(t_2792), .cout(t_2793));
compressor_4_2 u2_957(.a(s_119_49), .b(s_119_48), .c(s_119_47), .d(s_119_46), .cin(s_119_45), .o(t_2794), .co(t_2795), .cout(t_2796));
compressor_4_2 u2_958(.a(s_119_54), .b(s_119_53), .c(s_119_52), .d(s_119_51), .cin(s_119_50), .o(t_2797), .co(t_2798), .cout(t_2799));
compressor_4_2 u2_959(.a(s_119_59), .b(s_119_58), .c(s_119_57), .d(s_119_56), .cin(s_119_55), .o(t_2800), .co(t_2801), .cout(t_2802));
compressor_4_2 u2_960(.a(s_120_2), .b(s_120_1), .c(s_120_0), .d(t_2760), .cin(t_2763), .o(t_2803), .co(t_2804), .cout(t_2805));
compressor_4_2 u2_961(.a(s_120_5), .b(s_120_4), .c(s_120_3), .d(t_2766), .cin(t_2769), .o(t_2806), .co(t_2807), .cout(t_2808));
compressor_4_2 u2_962(.a(s_120_8), .b(s_120_7), .c(s_120_6), .d(t_2772), .cin(t_2775), .o(t_2809), .co(t_2810), .cout(t_2811));
compressor_4_2 u2_963(.a(s_120_11), .b(s_120_10), .c(s_120_9), .d(t_2778), .cin(t_2781), .o(t_2812), .co(t_2813), .cout(t_2814));
compressor_4_2 u2_964(.a(s_120_14), .b(s_120_13), .c(s_120_12), .d(t_2784), .cin(t_2787), .o(t_2815), .co(t_2816), .cout(t_2817));
compressor_4_2 u2_965(.a(s_120_17), .b(s_120_16), .c(s_120_15), .d(t_2790), .cin(t_2793), .o(t_2818), .co(t_2819), .cout(t_2820));
compressor_4_2 u2_966(.a(s_120_20), .b(s_120_19), .c(s_120_18), .d(t_2796), .cin(t_2799), .o(t_2821), .co(t_2822), .cout(t_2823));
compressor_4_2 u2_967(.a(s_120_24), .b(s_120_23), .c(s_120_22), .d(s_120_21), .cin(t_2802), .o(t_2824), .co(t_2825), .cout(t_2826));
compressor_4_2 u2_968(.a(s_120_29), .b(s_120_28), .c(s_120_27), .d(s_120_26), .cin(s_120_25), .o(t_2827), .co(t_2828), .cout(t_2829));
compressor_4_2 u2_969(.a(s_120_34), .b(s_120_33), .c(s_120_32), .d(s_120_31), .cin(s_120_30), .o(t_2830), .co(t_2831), .cout(t_2832));
compressor_4_2 u2_970(.a(s_120_39), .b(s_120_38), .c(s_120_37), .d(s_120_36), .cin(s_120_35), .o(t_2833), .co(t_2834), .cout(t_2835));
compressor_4_2 u2_971(.a(s_120_44), .b(s_120_43), .c(s_120_42), .d(s_120_41), .cin(s_120_40), .o(t_2836), .co(t_2837), .cout(t_2838));
compressor_4_2 u2_972(.a(s_120_49), .b(s_120_48), .c(s_120_47), .d(s_120_46), .cin(s_120_45), .o(t_2839), .co(t_2840), .cout(t_2841));
compressor_4_2 u2_973(.a(s_120_54), .b(s_120_53), .c(s_120_52), .d(s_120_51), .cin(s_120_50), .o(t_2842), .co(t_2843), .cout(t_2844));
compressor_4_2 u2_974(.a(s_120_59), .b(s_120_58), .c(s_120_57), .d(s_120_56), .cin(s_120_55), .o(t_2845), .co(t_2846), .cout(t_2847));
half_adder u0_975(.a(s_120_61), .b(s_120_60), .o(t_2848), .cout(t_2849));
compressor_4_2 u2_976(.a(s_121_2), .b(s_121_1), .c(s_121_0), .d(t_2805), .cin(t_2808), .o(t_2850), .co(t_2851), .cout(t_2852));
compressor_4_2 u2_977(.a(s_121_5), .b(s_121_4), .c(s_121_3), .d(t_2811), .cin(t_2814), .o(t_2853), .co(t_2854), .cout(t_2855));
compressor_4_2 u2_978(.a(s_121_8), .b(s_121_7), .c(s_121_6), .d(t_2817), .cin(t_2820), .o(t_2856), .co(t_2857), .cout(t_2858));
compressor_4_2 u2_979(.a(s_121_11), .b(s_121_10), .c(s_121_9), .d(t_2823), .cin(t_2826), .o(t_2859), .co(t_2860), .cout(t_2861));
compressor_4_2 u2_980(.a(s_121_14), .b(s_121_13), .c(s_121_12), .d(t_2829), .cin(t_2832), .o(t_2862), .co(t_2863), .cout(t_2864));
compressor_4_2 u2_981(.a(s_121_17), .b(s_121_16), .c(s_121_15), .d(t_2835), .cin(t_2838), .o(t_2865), .co(t_2866), .cout(t_2867));
compressor_4_2 u2_982(.a(s_121_20), .b(s_121_19), .c(s_121_18), .d(t_2841), .cin(t_2844), .o(t_2868), .co(t_2869), .cout(t_2870));
compressor_4_2 u2_983(.a(s_121_23), .b(s_121_22), .c(s_121_21), .d(t_2847), .cin(t_2849), .o(t_2871), .co(t_2872), .cout(t_2873));
compressor_4_2 u2_984(.a(s_121_28), .b(s_121_27), .c(s_121_26), .d(s_121_25), .cin(s_121_24), .o(t_2874), .co(t_2875), .cout(t_2876));
compressor_4_2 u2_985(.a(s_121_33), .b(s_121_32), .c(s_121_31), .d(s_121_30), .cin(s_121_29), .o(t_2877), .co(t_2878), .cout(t_2879));
compressor_4_2 u2_986(.a(s_121_38), .b(s_121_37), .c(s_121_36), .d(s_121_35), .cin(s_121_34), .o(t_2880), .co(t_2881), .cout(t_2882));
compressor_4_2 u2_987(.a(s_121_43), .b(s_121_42), .c(s_121_41), .d(s_121_40), .cin(s_121_39), .o(t_2883), .co(t_2884), .cout(t_2885));
compressor_4_2 u2_988(.a(s_121_48), .b(s_121_47), .c(s_121_46), .d(s_121_45), .cin(s_121_44), .o(t_2886), .co(t_2887), .cout(t_2888));
compressor_4_2 u2_989(.a(s_121_53), .b(s_121_52), .c(s_121_51), .d(s_121_50), .cin(s_121_49), .o(t_2889), .co(t_2890), .cout(t_2891));
compressor_4_2 u2_990(.a(s_121_58), .b(s_121_57), .c(s_121_56), .d(s_121_55), .cin(s_121_54), .o(t_2892), .co(t_2893), .cout(t_2894));
half_adder u0_991(.a(s_121_60), .b(s_121_59), .o(t_2895), .cout(t_2896));
compressor_4_2 u2_992(.a(s_122_2), .b(s_122_1), .c(s_122_0), .d(t_2852), .cin(t_2855), .o(t_2897), .co(t_2898), .cout(t_2899));
compressor_4_2 u2_993(.a(s_122_5), .b(s_122_4), .c(s_122_3), .d(t_2858), .cin(t_2861), .o(t_2900), .co(t_2901), .cout(t_2902));
compressor_4_2 u2_994(.a(s_122_8), .b(s_122_7), .c(s_122_6), .d(t_2864), .cin(t_2867), .o(t_2903), .co(t_2904), .cout(t_2905));
compressor_4_2 u2_995(.a(s_122_11), .b(s_122_10), .c(s_122_9), .d(t_2870), .cin(t_2873), .o(t_2906), .co(t_2907), .cout(t_2908));
compressor_4_2 u2_996(.a(s_122_14), .b(s_122_13), .c(s_122_12), .d(t_2876), .cin(t_2879), .o(t_2909), .co(t_2910), .cout(t_2911));
compressor_4_2 u2_997(.a(s_122_17), .b(s_122_16), .c(s_122_15), .d(t_2882), .cin(t_2885), .o(t_2912), .co(t_2913), .cout(t_2914));
compressor_4_2 u2_998(.a(s_122_20), .b(s_122_19), .c(s_122_18), .d(t_2888), .cin(t_2891), .o(t_2915), .co(t_2916), .cout(t_2917));
compressor_4_2 u2_999(.a(s_122_23), .b(s_122_22), .c(s_122_21), .d(t_2894), .cin(t_2896), .o(t_2918), .co(t_2919), .cout(t_2920));
compressor_4_2 u2_1000(.a(s_122_28), .b(s_122_27), .c(s_122_26), .d(s_122_25), .cin(s_122_24), .o(t_2921), .co(t_2922), .cout(t_2923));
compressor_4_2 u2_1001(.a(s_122_33), .b(s_122_32), .c(s_122_31), .d(s_122_30), .cin(s_122_29), .o(t_2924), .co(t_2925), .cout(t_2926));
compressor_4_2 u2_1002(.a(s_122_38), .b(s_122_37), .c(s_122_36), .d(s_122_35), .cin(s_122_34), .o(t_2927), .co(t_2928), .cout(t_2929));
compressor_4_2 u2_1003(.a(s_122_43), .b(s_122_42), .c(s_122_41), .d(s_122_40), .cin(s_122_39), .o(t_2930), .co(t_2931), .cout(t_2932));
compressor_4_2 u2_1004(.a(s_122_48), .b(s_122_47), .c(s_122_46), .d(s_122_45), .cin(s_122_44), .o(t_2933), .co(t_2934), .cout(t_2935));
compressor_4_2 u2_1005(.a(s_122_53), .b(s_122_52), .c(s_122_51), .d(s_122_50), .cin(s_122_49), .o(t_2936), .co(t_2937), .cout(t_2938));
compressor_4_2 u2_1006(.a(s_122_58), .b(s_122_57), .c(s_122_56), .d(s_122_55), .cin(s_122_54), .o(t_2939), .co(t_2940), .cout(t_2941));
compressor_3_2 u1_1007(.a(s_122_61), .b(s_122_60), .cin(s_122_59), .o(t_2942), .cout(t_2943));
compressor_4_2 u2_1008(.a(s_123_2), .b(s_123_1), .c(s_123_0), .d(t_2899), .cin(t_2902), .o(t_2944), .co(t_2945), .cout(t_2946));
compressor_4_2 u2_1009(.a(s_123_5), .b(s_123_4), .c(s_123_3), .d(t_2905), .cin(t_2908), .o(t_2947), .co(t_2948), .cout(t_2949));
compressor_4_2 u2_1010(.a(s_123_8), .b(s_123_7), .c(s_123_6), .d(t_2911), .cin(t_2914), .o(t_2950), .co(t_2951), .cout(t_2952));
compressor_4_2 u2_1011(.a(s_123_11), .b(s_123_10), .c(s_123_9), .d(t_2917), .cin(t_2920), .o(t_2953), .co(t_2954), .cout(t_2955));
compressor_4_2 u2_1012(.a(s_123_14), .b(s_123_13), .c(s_123_12), .d(t_2923), .cin(t_2926), .o(t_2956), .co(t_2957), .cout(t_2958));
compressor_4_2 u2_1013(.a(s_123_17), .b(s_123_16), .c(s_123_15), .d(t_2929), .cin(t_2932), .o(t_2959), .co(t_2960), .cout(t_2961));
compressor_4_2 u2_1014(.a(s_123_20), .b(s_123_19), .c(s_123_18), .d(t_2935), .cin(t_2938), .o(t_2962), .co(t_2963), .cout(t_2964));
compressor_4_2 u2_1015(.a(s_123_23), .b(s_123_22), .c(s_123_21), .d(t_2941), .cin(t_2943), .o(t_2965), .co(t_2966), .cout(t_2967));
compressor_4_2 u2_1016(.a(s_123_28), .b(s_123_27), .c(s_123_26), .d(s_123_25), .cin(s_123_24), .o(t_2968), .co(t_2969), .cout(t_2970));
compressor_4_2 u2_1017(.a(s_123_33), .b(s_123_32), .c(s_123_31), .d(s_123_30), .cin(s_123_29), .o(t_2971), .co(t_2972), .cout(t_2973));
compressor_4_2 u2_1018(.a(s_123_38), .b(s_123_37), .c(s_123_36), .d(s_123_35), .cin(s_123_34), .o(t_2974), .co(t_2975), .cout(t_2976));
compressor_4_2 u2_1019(.a(s_123_43), .b(s_123_42), .c(s_123_41), .d(s_123_40), .cin(s_123_39), .o(t_2977), .co(t_2978), .cout(t_2979));
compressor_4_2 u2_1020(.a(s_123_48), .b(s_123_47), .c(s_123_46), .d(s_123_45), .cin(s_123_44), .o(t_2980), .co(t_2981), .cout(t_2982));
compressor_4_2 u2_1021(.a(s_123_53), .b(s_123_52), .c(s_123_51), .d(s_123_50), .cin(s_123_49), .o(t_2983), .co(t_2984), .cout(t_2985));
compressor_4_2 u2_1022(.a(s_123_58), .b(s_123_57), .c(s_123_56), .d(s_123_55), .cin(s_123_54), .o(t_2986), .co(t_2987), .cout(t_2988));
compressor_3_2 u1_1023(.a(s_123_61), .b(s_123_60), .cin(s_123_59), .o(t_2989), .cout(t_2990));
compressor_4_2 u2_1024(.a(s_124_2), .b(s_124_1), .c(s_124_0), .d(t_2946), .cin(t_2949), .o(t_2991), .co(t_2992), .cout(t_2993));
compressor_4_2 u2_1025(.a(s_124_5), .b(s_124_4), .c(s_124_3), .d(t_2952), .cin(t_2955), .o(t_2994), .co(t_2995), .cout(t_2996));
compressor_4_2 u2_1026(.a(s_124_8), .b(s_124_7), .c(s_124_6), .d(t_2958), .cin(t_2961), .o(t_2997), .co(t_2998), .cout(t_2999));
compressor_4_2 u2_1027(.a(s_124_11), .b(s_124_10), .c(s_124_9), .d(t_2964), .cin(t_2967), .o(t_3000), .co(t_3001), .cout(t_3002));
compressor_4_2 u2_1028(.a(s_124_14), .b(s_124_13), .c(s_124_12), .d(t_2970), .cin(t_2973), .o(t_3003), .co(t_3004), .cout(t_3005));
compressor_4_2 u2_1029(.a(s_124_17), .b(s_124_16), .c(s_124_15), .d(t_2976), .cin(t_2979), .o(t_3006), .co(t_3007), .cout(t_3008));
compressor_4_2 u2_1030(.a(s_124_20), .b(s_124_19), .c(s_124_18), .d(t_2982), .cin(t_2985), .o(t_3009), .co(t_3010), .cout(t_3011));
compressor_4_2 u2_1031(.a(s_124_23), .b(s_124_22), .c(s_124_21), .d(t_2988), .cin(t_2990), .o(t_3012), .co(t_3013), .cout(t_3014));
compressor_4_2 u2_1032(.a(s_124_28), .b(s_124_27), .c(s_124_26), .d(s_124_25), .cin(s_124_24), .o(t_3015), .co(t_3016), .cout(t_3017));
compressor_4_2 u2_1033(.a(s_124_33), .b(s_124_32), .c(s_124_31), .d(s_124_30), .cin(s_124_29), .o(t_3018), .co(t_3019), .cout(t_3020));
compressor_4_2 u2_1034(.a(s_124_38), .b(s_124_37), .c(s_124_36), .d(s_124_35), .cin(s_124_34), .o(t_3021), .co(t_3022), .cout(t_3023));
compressor_4_2 u2_1035(.a(s_124_43), .b(s_124_42), .c(s_124_41), .d(s_124_40), .cin(s_124_39), .o(t_3024), .co(t_3025), .cout(t_3026));
compressor_4_2 u2_1036(.a(s_124_48), .b(s_124_47), .c(s_124_46), .d(s_124_45), .cin(s_124_44), .o(t_3027), .co(t_3028), .cout(t_3029));
compressor_4_2 u2_1037(.a(s_124_53), .b(s_124_52), .c(s_124_51), .d(s_124_50), .cin(s_124_49), .o(t_3030), .co(t_3031), .cout(t_3032));
compressor_4_2 u2_1038(.a(s_124_58), .b(s_124_57), .c(s_124_56), .d(s_124_55), .cin(s_124_54), .o(t_3033), .co(t_3034), .cout(t_3035));
compressor_4_2 u2_1039(.a(s_124_63), .b(s_124_62), .c(s_124_61), .d(s_124_60), .cin(s_124_59), .o(t_3036), .co(t_3037), .cout(t_3038));
compressor_4_2 u2_1040(.a(s_125_2), .b(s_125_1), .c(s_125_0), .d(t_2993), .cin(t_2996), .o(t_3039), .co(t_3040), .cout(t_3041));
compressor_4_2 u2_1041(.a(s_125_5), .b(s_125_4), .c(s_125_3), .d(t_2999), .cin(t_3002), .o(t_3042), .co(t_3043), .cout(t_3044));
compressor_4_2 u2_1042(.a(s_125_8), .b(s_125_7), .c(s_125_6), .d(t_3005), .cin(t_3008), .o(t_3045), .co(t_3046), .cout(t_3047));
compressor_4_2 u2_1043(.a(s_125_11), .b(s_125_10), .c(s_125_9), .d(t_3011), .cin(t_3014), .o(t_3048), .co(t_3049), .cout(t_3050));
compressor_4_2 u2_1044(.a(s_125_14), .b(s_125_13), .c(s_125_12), .d(t_3017), .cin(t_3020), .o(t_3051), .co(t_3052), .cout(t_3053));
compressor_4_2 u2_1045(.a(s_125_17), .b(s_125_16), .c(s_125_15), .d(t_3023), .cin(t_3026), .o(t_3054), .co(t_3055), .cout(t_3056));
compressor_4_2 u2_1046(.a(s_125_20), .b(s_125_19), .c(s_125_18), .d(t_3029), .cin(t_3032), .o(t_3057), .co(t_3058), .cout(t_3059));
compressor_4_2 u2_1047(.a(s_125_23), .b(s_125_22), .c(s_125_21), .d(t_3035), .cin(t_3038), .o(t_3060), .co(t_3061), .cout(t_3062));
compressor_4_2 u2_1048(.a(s_125_28), .b(s_125_27), .c(s_125_26), .d(s_125_25), .cin(s_125_24), .o(t_3063), .co(t_3064), .cout(t_3065));
compressor_4_2 u2_1049(.a(s_125_33), .b(s_125_32), .c(s_125_31), .d(s_125_30), .cin(s_125_29), .o(t_3066), .co(t_3067), .cout(t_3068));
compressor_4_2 u2_1050(.a(s_125_38), .b(s_125_37), .c(s_125_36), .d(s_125_35), .cin(s_125_34), .o(t_3069), .co(t_3070), .cout(t_3071));
compressor_4_2 u2_1051(.a(s_125_43), .b(s_125_42), .c(s_125_41), .d(s_125_40), .cin(s_125_39), .o(t_3072), .co(t_3073), .cout(t_3074));
compressor_4_2 u2_1052(.a(s_125_48), .b(s_125_47), .c(s_125_46), .d(s_125_45), .cin(s_125_44), .o(t_3075), .co(t_3076), .cout(t_3077));
compressor_4_2 u2_1053(.a(s_125_53), .b(s_125_52), .c(s_125_51), .d(s_125_50), .cin(s_125_49), .o(t_3078), .co(t_3079), .cout(t_3080));
compressor_4_2 u2_1054(.a(s_125_58), .b(s_125_57), .c(s_125_56), .d(s_125_55), .cin(s_125_54), .o(t_3081), .co(t_3082), .cout(t_3083));
compressor_3_2 u1_1055(.a(s_125_61), .b(s_125_60), .cin(s_125_59), .o(t_3084), .cout(t_3085));
compressor_4_2 u2_1056(.a(s_126_2), .b(s_126_1), .c(s_126_0), .d(t_3041), .cin(t_3044), .o(t_3086), .co(t_3087), .cout(t_3088));
compressor_4_2 u2_1057(.a(s_126_5), .b(s_126_4), .c(s_126_3), .d(t_3047), .cin(t_3050), .o(t_3089), .co(t_3090), .cout(t_3091));
compressor_4_2 u2_1058(.a(s_126_8), .b(s_126_7), .c(s_126_6), .d(t_3053), .cin(t_3056), .o(t_3092), .co(t_3093), .cout(t_3094));
compressor_4_2 u2_1059(.a(s_126_11), .b(s_126_10), .c(s_126_9), .d(t_3059), .cin(t_3062), .o(t_3095), .co(t_3096), .cout(t_3097));
compressor_4_2 u2_1060(.a(s_126_14), .b(s_126_13), .c(s_126_12), .d(t_3065), .cin(t_3068), .o(t_3098), .co(t_3099), .cout(t_3100));
compressor_4_2 u2_1061(.a(s_126_17), .b(s_126_16), .c(s_126_15), .d(t_3071), .cin(t_3074), .o(t_3101), .co(t_3102), .cout(t_3103));
compressor_4_2 u2_1062(.a(s_126_20), .b(s_126_19), .c(s_126_18), .d(t_3077), .cin(t_3080), .o(t_3104), .co(t_3105), .cout(t_3106));
compressor_4_2 u2_1063(.a(s_126_23), .b(s_126_22), .c(s_126_21), .d(t_3083), .cin(t_3085), .o(t_3107), .co(t_3108), .cout(t_3109));
compressor_4_2 u2_1064(.a(s_126_28), .b(s_126_27), .c(s_126_26), .d(s_126_25), .cin(s_126_24), .o(t_3110), .co(t_3111), .cout(t_3112));
compressor_4_2 u2_1065(.a(s_126_33), .b(s_126_32), .c(s_126_31), .d(s_126_30), .cin(s_126_29), .o(t_3113), .co(t_3114), .cout(t_3115));
compressor_4_2 u2_1066(.a(s_126_38), .b(s_126_37), .c(s_126_36), .d(s_126_35), .cin(s_126_34), .o(t_3116), .co(t_3117), .cout(t_3118));
compressor_4_2 u2_1067(.a(s_126_43), .b(s_126_42), .c(s_126_41), .d(s_126_40), .cin(s_126_39), .o(t_3119), .co(t_3120), .cout(t_3121));
compressor_4_2 u2_1068(.a(s_126_48), .b(s_126_47), .c(s_126_46), .d(s_126_45), .cin(s_126_44), .o(t_3122), .co(t_3123), .cout(t_3124));
compressor_4_2 u2_1069(.a(s_126_53), .b(s_126_52), .c(s_126_51), .d(s_126_50), .cin(s_126_49), .o(t_3125), .co(t_3126), .cout(t_3127));
compressor_4_2 u2_1070(.a(s_126_58), .b(s_126_57), .c(s_126_56), .d(s_126_55), .cin(s_126_54), .o(t_3128), .co(t_3129), .cout(t_3130));
compressor_4_2 u2_1071(.a(s_126_63), .b(s_126_62), .c(s_126_61), .d(s_126_60), .cin(s_126_59), .o(t_3131), .co(t_3132), .cout(t_3133));
compressor_4_2 u2_1072(.a(s_127_2), .b(s_127_1), .c(s_127_0), .d(t_3088), .cin(t_3091), .o(t_3134), .co(t_3135), .cout(t_3136));
compressor_4_2 u2_1073(.a(s_127_5), .b(s_127_4), .c(s_127_3), .d(t_3094), .cin(t_3097), .o(t_3137), .co(t_3138), .cout(t_3139));
compressor_4_2 u2_1074(.a(s_127_8), .b(s_127_7), .c(s_127_6), .d(t_3100), .cin(t_3103), .o(t_3140), .co(t_3141), .cout(t_3142));
compressor_4_2 u2_1075(.a(s_127_11), .b(s_127_10), .c(s_127_9), .d(t_3106), .cin(t_3109), .o(t_3143), .co(t_3144), .cout(t_3145));
compressor_4_2 u2_1076(.a(s_127_14), .b(s_127_13), .c(s_127_12), .d(t_3112), .cin(t_3115), .o(t_3146), .co(t_3147), .cout(t_3148));
compressor_4_2 u2_1077(.a(s_127_17), .b(s_127_16), .c(s_127_15), .d(t_3118), .cin(t_3121), .o(t_3149), .co(t_3150), .cout(t_3151));
compressor_4_2 u2_1078(.a(s_127_20), .b(s_127_19), .c(s_127_18), .d(t_3124), .cin(t_3127), .o(t_3152), .co(t_3153), .cout(t_3154));
compressor_4_2 u2_1079(.a(s_127_23), .b(s_127_22), .c(s_127_21), .d(t_3130), .cin(t_3133), .o(t_3155), .co(t_3156), .cout(t_3157));
compressor_4_2 u2_1080(.a(s_127_28), .b(s_127_27), .c(s_127_26), .d(s_127_25), .cin(s_127_24), .o(t_3158), .co(t_3159), .cout(t_3160));
compressor_4_2 u2_1081(.a(s_127_33), .b(s_127_32), .c(s_127_31), .d(s_127_30), .cin(s_127_29), .o(t_3161), .co(t_3162), .cout(t_3163));
compressor_4_2 u2_1082(.a(s_127_38), .b(s_127_37), .c(s_127_36), .d(s_127_35), .cin(s_127_34), .o(t_3164), .co(t_3165), .cout(t_3166));
compressor_4_2 u2_1083(.a(s_127_43), .b(s_127_42), .c(s_127_41), .d(s_127_40), .cin(s_127_39), .o(t_3167), .co(t_3168), .cout(t_3169));
compressor_4_2 u2_1084(.a(s_127_48), .b(s_127_47), .c(s_127_46), .d(s_127_45), .cin(s_127_44), .o(t_3170), .co(t_3171), .cout(t_3172));
compressor_4_2 u2_1085(.a(s_127_53), .b(s_127_52), .c(s_127_51), .d(s_127_50), .cin(s_127_49), .o(t_3173), .co(t_3174), .cout(t_3175));
compressor_4_2 u2_1086(.a(s_127_58), .b(s_127_57), .c(s_127_56), .d(s_127_55), .cin(s_127_54), .o(t_3176), .co(t_3177), .cout(t_3178));
compressor_4_2 u2_1087(.a(s_127_63), .b(s_127_62), .c(s_127_61), .d(s_127_60), .cin(s_127_59), .o(t_3179), .co(t_3180), .cout(t_3181));
compressor_4_2 u2_1088(.a(s_128_2), .b(s_128_1), .c(s_128_0), .d(t_3136), .cin(t_3139), .o(t_3182), .co(t_3183), .cout(t_3184));
compressor_4_2 u2_1089(.a(s_128_5), .b(s_128_4), .c(s_128_3), .d(t_3142), .cin(t_3145), .o(t_3185), .co(t_3186), .cout(t_3187));
compressor_4_2 u2_1090(.a(s_128_8), .b(s_128_7), .c(s_128_6), .d(t_3148), .cin(t_3151), .o(t_3188), .co(t_3189), .cout(t_3190));
compressor_4_2 u2_1091(.a(s_128_11), .b(s_128_10), .c(s_128_9), .d(t_3154), .cin(t_3157), .o(t_3191), .co(t_3192), .cout(t_3193));
compressor_4_2 u2_1092(.a(s_128_14), .b(s_128_13), .c(s_128_12), .d(t_3160), .cin(t_3163), .o(t_3194), .co(t_3195), .cout(t_3196));
compressor_4_2 u2_1093(.a(s_128_17), .b(s_128_16), .c(s_128_15), .d(t_3166), .cin(t_3169), .o(t_3197), .co(t_3198), .cout(t_3199));
compressor_4_2 u2_1094(.a(s_128_20), .b(s_128_19), .c(s_128_18), .d(t_3172), .cin(t_3175), .o(t_3200), .co(t_3201), .cout(t_3202));
compressor_4_2 u2_1095(.a(s_128_23), .b(s_128_22), .c(s_128_21), .d(t_3178), .cin(t_3181), .o(t_3203), .co(t_3204), .cout(t_3205));
compressor_4_2 u2_1096(.a(s_128_28), .b(s_128_27), .c(s_128_26), .d(s_128_25), .cin(s_128_24), .o(t_3206), .co(t_3207), .cout(t_3208));
compressor_4_2 u2_1097(.a(s_128_33), .b(s_128_32), .c(s_128_31), .d(s_128_30), .cin(s_128_29), .o(t_3209), .co(t_3210), .cout(t_3211));
compressor_4_2 u2_1098(.a(s_128_38), .b(s_128_37), .c(s_128_36), .d(s_128_35), .cin(s_128_34), .o(t_3212), .co(t_3213), .cout(t_3214));
compressor_4_2 u2_1099(.a(s_128_43), .b(s_128_42), .c(s_128_41), .d(s_128_40), .cin(s_128_39), .o(t_3215), .co(t_3216), .cout(t_3217));
compressor_4_2 u2_1100(.a(s_128_48), .b(s_128_47), .c(s_128_46), .d(s_128_45), .cin(s_128_44), .o(t_3218), .co(t_3219), .cout(t_3220));
compressor_4_2 u2_1101(.a(s_128_53), .b(s_128_52), .c(s_128_51), .d(s_128_50), .cin(s_128_49), .o(t_3221), .co(t_3222), .cout(t_3223));
compressor_4_2 u2_1102(.a(s_128_58), .b(s_128_57), .c(s_128_56), .d(s_128_55), .cin(s_128_54), .o(t_3224), .co(t_3225), .cout(t_3226));
compressor_4_2 u2_1103(.a(s_128_63), .b(s_128_62), .c(s_128_61), .d(s_128_60), .cin(s_128_59), .o(t_3227), .co(t_3228), .cout(t_3229));
compressor_4_2 u2_1104(.a(s_129_2), .b(s_129_1), .c(s_129_0), .d(t_3184), .cin(t_3187), .o(t_3230), .co(t_3231), .cout(t_3232));
compressor_4_2 u2_1105(.a(s_129_5), .b(s_129_4), .c(s_129_3), .d(t_3190), .cin(t_3193), .o(t_3233), .co(t_3234), .cout(t_3235));
compressor_4_2 u2_1106(.a(s_129_8), .b(s_129_7), .c(s_129_6), .d(t_3196), .cin(t_3199), .o(t_3236), .co(t_3237), .cout(t_3238));
compressor_4_2 u2_1107(.a(s_129_11), .b(s_129_10), .c(s_129_9), .d(t_3202), .cin(t_3205), .o(t_3239), .co(t_3240), .cout(t_3241));
compressor_4_2 u2_1108(.a(s_129_14), .b(s_129_13), .c(s_129_12), .d(t_3208), .cin(t_3211), .o(t_3242), .co(t_3243), .cout(t_3244));
compressor_4_2 u2_1109(.a(s_129_17), .b(s_129_16), .c(s_129_15), .d(t_3214), .cin(t_3217), .o(t_3245), .co(t_3246), .cout(t_3247));
compressor_4_2 u2_1110(.a(s_129_20), .b(s_129_19), .c(s_129_18), .d(t_3220), .cin(t_3223), .o(t_3248), .co(t_3249), .cout(t_3250));
compressor_4_2 u2_1111(.a(s_129_23), .b(s_129_22), .c(s_129_21), .d(t_3226), .cin(t_3229), .o(t_3251), .co(t_3252), .cout(t_3253));
compressor_4_2 u2_1112(.a(s_129_28), .b(s_129_27), .c(s_129_26), .d(s_129_25), .cin(s_129_24), .o(t_3254), .co(t_3255), .cout(t_3256));
compressor_4_2 u2_1113(.a(s_129_33), .b(s_129_32), .c(s_129_31), .d(s_129_30), .cin(s_129_29), .o(t_3257), .co(t_3258), .cout(t_3259));
compressor_4_2 u2_1114(.a(s_129_38), .b(s_129_37), .c(s_129_36), .d(s_129_35), .cin(s_129_34), .o(t_3260), .co(t_3261), .cout(t_3262));
compressor_4_2 u2_1115(.a(s_129_43), .b(s_129_42), .c(s_129_41), .d(s_129_40), .cin(s_129_39), .o(t_3263), .co(t_3264), .cout(t_3265));
compressor_4_2 u2_1116(.a(s_129_48), .b(s_129_47), .c(s_129_46), .d(s_129_45), .cin(s_129_44), .o(t_3266), .co(t_3267), .cout(t_3268));
compressor_4_2 u2_1117(.a(s_129_53), .b(s_129_52), .c(s_129_51), .d(s_129_50), .cin(s_129_49), .o(t_3269), .co(t_3270), .cout(t_3271));
compressor_4_2 u2_1118(.a(s_129_58), .b(s_129_57), .c(s_129_56), .d(s_129_55), .cin(s_129_54), .o(t_3272), .co(t_3273), .cout(t_3274));
compressor_4_2 u2_1119(.a(s_129_63), .b(s_129_62), .c(s_129_61), .d(s_129_60), .cin(s_129_59), .o(t_3275), .co(t_3276), .cout(t_3277));
compressor_4_2 u2_1120(.a(s_130_2), .b(s_130_1), .c(s_130_0), .d(t_3232), .cin(t_3235), .o(t_3278), .co(t_3279), .cout(t_3280));
compressor_4_2 u2_1121(.a(s_130_5), .b(s_130_4), .c(s_130_3), .d(t_3238), .cin(t_3241), .o(t_3281), .co(t_3282), .cout(t_3283));
compressor_4_2 u2_1122(.a(s_130_8), .b(s_130_7), .c(s_130_6), .d(t_3244), .cin(t_3247), .o(t_3284), .co(t_3285), .cout(t_3286));
compressor_4_2 u2_1123(.a(s_130_11), .b(s_130_10), .c(s_130_9), .d(t_3250), .cin(t_3253), .o(t_3287), .co(t_3288), .cout(t_3289));
compressor_4_2 u2_1124(.a(s_130_14), .b(s_130_13), .c(s_130_12), .d(t_3256), .cin(t_3259), .o(t_3290), .co(t_3291), .cout(t_3292));
compressor_4_2 u2_1125(.a(s_130_17), .b(s_130_16), .c(s_130_15), .d(t_3262), .cin(t_3265), .o(t_3293), .co(t_3294), .cout(t_3295));
compressor_4_2 u2_1126(.a(s_130_20), .b(s_130_19), .c(s_130_18), .d(t_3268), .cin(t_3271), .o(t_3296), .co(t_3297), .cout(t_3298));
compressor_4_2 u2_1127(.a(s_130_23), .b(s_130_22), .c(s_130_21), .d(t_3274), .cin(t_3277), .o(t_3299), .co(t_3300), .cout(t_3301));
compressor_4_2 u2_1128(.a(s_130_28), .b(s_130_27), .c(s_130_26), .d(s_130_25), .cin(s_130_24), .o(t_3302), .co(t_3303), .cout(t_3304));
compressor_4_2 u2_1129(.a(s_130_33), .b(s_130_32), .c(s_130_31), .d(s_130_30), .cin(s_130_29), .o(t_3305), .co(t_3306), .cout(t_3307));
compressor_4_2 u2_1130(.a(s_130_38), .b(s_130_37), .c(s_130_36), .d(s_130_35), .cin(s_130_34), .o(t_3308), .co(t_3309), .cout(t_3310));
compressor_4_2 u2_1131(.a(s_130_43), .b(s_130_42), .c(s_130_41), .d(s_130_40), .cin(s_130_39), .o(t_3311), .co(t_3312), .cout(t_3313));
compressor_4_2 u2_1132(.a(s_130_48), .b(s_130_47), .c(s_130_46), .d(s_130_45), .cin(s_130_44), .o(t_3314), .co(t_3315), .cout(t_3316));
compressor_4_2 u2_1133(.a(s_130_53), .b(s_130_52), .c(s_130_51), .d(s_130_50), .cin(s_130_49), .o(t_3317), .co(t_3318), .cout(t_3319));
compressor_4_2 u2_1134(.a(s_130_58), .b(s_130_57), .c(s_130_56), .d(s_130_55), .cin(s_130_54), .o(t_3320), .co(t_3321), .cout(t_3322));
compressor_4_2 u2_1135(.a(s_130_63), .b(s_130_62), .c(s_130_61), .d(s_130_60), .cin(s_130_59), .o(t_3323), .co(t_3324), .cout(t_3325));
compressor_4_2 u2_1136(.a(s_131_2), .b(s_131_1), .c(s_131_0), .d(t_3280), .cin(t_3283), .o(t_3326), .co(t_3327), .cout(t_3328));
compressor_4_2 u2_1137(.a(s_131_5), .b(s_131_4), .c(s_131_3), .d(t_3286), .cin(t_3289), .o(t_3329), .co(t_3330), .cout(t_3331));
compressor_4_2 u2_1138(.a(s_131_8), .b(s_131_7), .c(s_131_6), .d(t_3292), .cin(t_3295), .o(t_3332), .co(t_3333), .cout(t_3334));
compressor_4_2 u2_1139(.a(s_131_11), .b(s_131_10), .c(s_131_9), .d(t_3298), .cin(t_3301), .o(t_3335), .co(t_3336), .cout(t_3337));
compressor_4_2 u2_1140(.a(s_131_14), .b(s_131_13), .c(s_131_12), .d(t_3304), .cin(t_3307), .o(t_3338), .co(t_3339), .cout(t_3340));
compressor_4_2 u2_1141(.a(s_131_17), .b(s_131_16), .c(s_131_15), .d(t_3310), .cin(t_3313), .o(t_3341), .co(t_3342), .cout(t_3343));
compressor_4_2 u2_1142(.a(s_131_20), .b(s_131_19), .c(s_131_18), .d(t_3316), .cin(t_3319), .o(t_3344), .co(t_3345), .cout(t_3346));
compressor_4_2 u2_1143(.a(s_131_23), .b(s_131_22), .c(s_131_21), .d(t_3322), .cin(t_3325), .o(t_3347), .co(t_3348), .cout(t_3349));
compressor_4_2 u2_1144(.a(s_131_28), .b(s_131_27), .c(s_131_26), .d(s_131_25), .cin(s_131_24), .o(t_3350), .co(t_3351), .cout(t_3352));
compressor_4_2 u2_1145(.a(s_131_33), .b(s_131_32), .c(s_131_31), .d(s_131_30), .cin(s_131_29), .o(t_3353), .co(t_3354), .cout(t_3355));
compressor_4_2 u2_1146(.a(s_131_38), .b(s_131_37), .c(s_131_36), .d(s_131_35), .cin(s_131_34), .o(t_3356), .co(t_3357), .cout(t_3358));
compressor_4_2 u2_1147(.a(s_131_43), .b(s_131_42), .c(s_131_41), .d(s_131_40), .cin(s_131_39), .o(t_3359), .co(t_3360), .cout(t_3361));
compressor_4_2 u2_1148(.a(s_131_48), .b(s_131_47), .c(s_131_46), .d(s_131_45), .cin(s_131_44), .o(t_3362), .co(t_3363), .cout(t_3364));
compressor_4_2 u2_1149(.a(s_131_53), .b(s_131_52), .c(s_131_51), .d(s_131_50), .cin(s_131_49), .o(t_3365), .co(t_3366), .cout(t_3367));
compressor_4_2 u2_1150(.a(s_131_58), .b(s_131_57), .c(s_131_56), .d(s_131_55), .cin(s_131_54), .o(t_3368), .co(t_3369), .cout(t_3370));
compressor_4_2 u2_1151(.a(s_131_63), .b(s_131_62), .c(s_131_61), .d(s_131_60), .cin(s_131_59), .o(t_3371), .co(t_3372), .cout(t_3373));
compressor_4_2 u2_1152(.a(s_132_2), .b(s_132_1), .c(s_132_0), .d(t_3328), .cin(t_3331), .o(t_3374), .co(t_3375), .cout(t_3376));
compressor_4_2 u2_1153(.a(s_132_5), .b(s_132_4), .c(s_132_3), .d(t_3334), .cin(t_3337), .o(t_3377), .co(t_3378), .cout(t_3379));
compressor_4_2 u2_1154(.a(s_132_8), .b(s_132_7), .c(s_132_6), .d(t_3340), .cin(t_3343), .o(t_3380), .co(t_3381), .cout(t_3382));
compressor_4_2 u2_1155(.a(s_132_11), .b(s_132_10), .c(s_132_9), .d(t_3346), .cin(t_3349), .o(t_3383), .co(t_3384), .cout(t_3385));
compressor_4_2 u2_1156(.a(s_132_14), .b(s_132_13), .c(s_132_12), .d(t_3352), .cin(t_3355), .o(t_3386), .co(t_3387), .cout(t_3388));
compressor_4_2 u2_1157(.a(s_132_17), .b(s_132_16), .c(s_132_15), .d(t_3358), .cin(t_3361), .o(t_3389), .co(t_3390), .cout(t_3391));
compressor_4_2 u2_1158(.a(s_132_20), .b(s_132_19), .c(s_132_18), .d(t_3364), .cin(t_3367), .o(t_3392), .co(t_3393), .cout(t_3394));
compressor_4_2 u2_1159(.a(s_132_23), .b(s_132_22), .c(s_132_21), .d(t_3370), .cin(t_3373), .o(t_3395), .co(t_3396), .cout(t_3397));
compressor_4_2 u2_1160(.a(s_132_28), .b(s_132_27), .c(s_132_26), .d(s_132_25), .cin(s_132_24), .o(t_3398), .co(t_3399), .cout(t_3400));
compressor_4_2 u2_1161(.a(s_132_33), .b(s_132_32), .c(s_132_31), .d(s_132_30), .cin(s_132_29), .o(t_3401), .co(t_3402), .cout(t_3403));
compressor_4_2 u2_1162(.a(s_132_38), .b(s_132_37), .c(s_132_36), .d(s_132_35), .cin(s_132_34), .o(t_3404), .co(t_3405), .cout(t_3406));
compressor_4_2 u2_1163(.a(s_132_43), .b(s_132_42), .c(s_132_41), .d(s_132_40), .cin(s_132_39), .o(t_3407), .co(t_3408), .cout(t_3409));
compressor_4_2 u2_1164(.a(s_132_48), .b(s_132_47), .c(s_132_46), .d(s_132_45), .cin(s_132_44), .o(t_3410), .co(t_3411), .cout(t_3412));
compressor_4_2 u2_1165(.a(s_132_53), .b(s_132_52), .c(s_132_51), .d(s_132_50), .cin(s_132_49), .o(t_3413), .co(t_3414), .cout(t_3415));
compressor_4_2 u2_1166(.a(s_132_58), .b(s_132_57), .c(s_132_56), .d(s_132_55), .cin(s_132_54), .o(t_3416), .co(t_3417), .cout(t_3418));
compressor_3_2 u1_1167(.a(s_132_61), .b(s_132_60), .cin(s_132_59), .o(t_3419), .cout(t_3420));
compressor_4_2 u2_1168(.a(s_133_2), .b(s_133_1), .c(s_133_0), .d(t_3376), .cin(t_3379), .o(t_3421), .co(t_3422), .cout(t_3423));
compressor_4_2 u2_1169(.a(s_133_5), .b(s_133_4), .c(s_133_3), .d(t_3382), .cin(t_3385), .o(t_3424), .co(t_3425), .cout(t_3426));
compressor_4_2 u2_1170(.a(s_133_8), .b(s_133_7), .c(s_133_6), .d(t_3388), .cin(t_3391), .o(t_3427), .co(t_3428), .cout(t_3429));
compressor_4_2 u2_1171(.a(s_133_11), .b(s_133_10), .c(s_133_9), .d(t_3394), .cin(t_3397), .o(t_3430), .co(t_3431), .cout(t_3432));
compressor_4_2 u2_1172(.a(s_133_14), .b(s_133_13), .c(s_133_12), .d(t_3400), .cin(t_3403), .o(t_3433), .co(t_3434), .cout(t_3435));
compressor_4_2 u2_1173(.a(s_133_17), .b(s_133_16), .c(s_133_15), .d(t_3406), .cin(t_3409), .o(t_3436), .co(t_3437), .cout(t_3438));
compressor_4_2 u2_1174(.a(s_133_20), .b(s_133_19), .c(s_133_18), .d(t_3412), .cin(t_3415), .o(t_3439), .co(t_3440), .cout(t_3441));
compressor_4_2 u2_1175(.a(s_133_23), .b(s_133_22), .c(s_133_21), .d(t_3418), .cin(t_3420), .o(t_3442), .co(t_3443), .cout(t_3444));
compressor_4_2 u2_1176(.a(s_133_28), .b(s_133_27), .c(s_133_26), .d(s_133_25), .cin(s_133_24), .o(t_3445), .co(t_3446), .cout(t_3447));
compressor_4_2 u2_1177(.a(s_133_33), .b(s_133_32), .c(s_133_31), .d(s_133_30), .cin(s_133_29), .o(t_3448), .co(t_3449), .cout(t_3450));
compressor_4_2 u2_1178(.a(s_133_38), .b(s_133_37), .c(s_133_36), .d(s_133_35), .cin(s_133_34), .o(t_3451), .co(t_3452), .cout(t_3453));
compressor_4_2 u2_1179(.a(s_133_43), .b(s_133_42), .c(s_133_41), .d(s_133_40), .cin(s_133_39), .o(t_3454), .co(t_3455), .cout(t_3456));
compressor_4_2 u2_1180(.a(s_133_48), .b(s_133_47), .c(s_133_46), .d(s_133_45), .cin(s_133_44), .o(t_3457), .co(t_3458), .cout(t_3459));
compressor_4_2 u2_1181(.a(s_133_53), .b(s_133_52), .c(s_133_51), .d(s_133_50), .cin(s_133_49), .o(t_3460), .co(t_3461), .cout(t_3462));
compressor_4_2 u2_1182(.a(s_133_58), .b(s_133_57), .c(s_133_56), .d(s_133_55), .cin(s_133_54), .o(t_3463), .co(t_3464), .cout(t_3465));
compressor_3_2 u1_1183(.a(s_133_61), .b(s_133_60), .cin(s_133_59), .o(t_3466), .cout(t_3467));
compressor_4_2 u2_1184(.a(s_134_2), .b(s_134_1), .c(s_134_0), .d(t_3423), .cin(t_3426), .o(t_3468), .co(t_3469), .cout(t_3470));
compressor_4_2 u2_1185(.a(s_134_5), .b(s_134_4), .c(s_134_3), .d(t_3429), .cin(t_3432), .o(t_3471), .co(t_3472), .cout(t_3473));
compressor_4_2 u2_1186(.a(s_134_8), .b(s_134_7), .c(s_134_6), .d(t_3435), .cin(t_3438), .o(t_3474), .co(t_3475), .cout(t_3476));
compressor_4_2 u2_1187(.a(s_134_11), .b(s_134_10), .c(s_134_9), .d(t_3441), .cin(t_3444), .o(t_3477), .co(t_3478), .cout(t_3479));
compressor_4_2 u2_1188(.a(s_134_14), .b(s_134_13), .c(s_134_12), .d(t_3447), .cin(t_3450), .o(t_3480), .co(t_3481), .cout(t_3482));
compressor_4_2 u2_1189(.a(s_134_17), .b(s_134_16), .c(s_134_15), .d(t_3453), .cin(t_3456), .o(t_3483), .co(t_3484), .cout(t_3485));
compressor_4_2 u2_1190(.a(s_134_20), .b(s_134_19), .c(s_134_18), .d(t_3459), .cin(t_3462), .o(t_3486), .co(t_3487), .cout(t_3488));
compressor_4_2 u2_1191(.a(s_134_23), .b(s_134_22), .c(s_134_21), .d(t_3465), .cin(t_3467), .o(t_3489), .co(t_3490), .cout(t_3491));
compressor_4_2 u2_1192(.a(s_134_28), .b(s_134_27), .c(s_134_26), .d(s_134_25), .cin(s_134_24), .o(t_3492), .co(t_3493), .cout(t_3494));
compressor_4_2 u2_1193(.a(s_134_33), .b(s_134_32), .c(s_134_31), .d(s_134_30), .cin(s_134_29), .o(t_3495), .co(t_3496), .cout(t_3497));
compressor_4_2 u2_1194(.a(s_134_38), .b(s_134_37), .c(s_134_36), .d(s_134_35), .cin(s_134_34), .o(t_3498), .co(t_3499), .cout(t_3500));
compressor_4_2 u2_1195(.a(s_134_43), .b(s_134_42), .c(s_134_41), .d(s_134_40), .cin(s_134_39), .o(t_3501), .co(t_3502), .cout(t_3503));
compressor_4_2 u2_1196(.a(s_134_48), .b(s_134_47), .c(s_134_46), .d(s_134_45), .cin(s_134_44), .o(t_3504), .co(t_3505), .cout(t_3506));
compressor_4_2 u2_1197(.a(s_134_53), .b(s_134_52), .c(s_134_51), .d(s_134_50), .cin(s_134_49), .o(t_3507), .co(t_3508), .cout(t_3509));
compressor_4_2 u2_1198(.a(s_134_58), .b(s_134_57), .c(s_134_56), .d(s_134_55), .cin(s_134_54), .o(t_3510), .co(t_3511), .cout(t_3512));
compressor_3_2 u1_1199(.a(s_134_61), .b(s_134_60), .cin(s_134_59), .o(t_3513), .cout(t_3514));
compressor_4_2 u2_1200(.a(s_135_2), .b(s_135_1), .c(s_135_0), .d(t_3470), .cin(t_3473), .o(t_3515), .co(t_3516), .cout(t_3517));
compressor_4_2 u2_1201(.a(s_135_5), .b(s_135_4), .c(s_135_3), .d(t_3476), .cin(t_3479), .o(t_3518), .co(t_3519), .cout(t_3520));
compressor_4_2 u2_1202(.a(s_135_8), .b(s_135_7), .c(s_135_6), .d(t_3482), .cin(t_3485), .o(t_3521), .co(t_3522), .cout(t_3523));
compressor_4_2 u2_1203(.a(s_135_11), .b(s_135_10), .c(s_135_9), .d(t_3488), .cin(t_3491), .o(t_3524), .co(t_3525), .cout(t_3526));
compressor_4_2 u2_1204(.a(s_135_14), .b(s_135_13), .c(s_135_12), .d(t_3494), .cin(t_3497), .o(t_3527), .co(t_3528), .cout(t_3529));
compressor_4_2 u2_1205(.a(s_135_17), .b(s_135_16), .c(s_135_15), .d(t_3500), .cin(t_3503), .o(t_3530), .co(t_3531), .cout(t_3532));
compressor_4_2 u2_1206(.a(s_135_20), .b(s_135_19), .c(s_135_18), .d(t_3506), .cin(t_3509), .o(t_3533), .co(t_3534), .cout(t_3535));
compressor_4_2 u2_1207(.a(s_135_23), .b(s_135_22), .c(s_135_21), .d(t_3512), .cin(t_3514), .o(t_3536), .co(t_3537), .cout(t_3538));
compressor_4_2 u2_1208(.a(s_135_28), .b(s_135_27), .c(s_135_26), .d(s_135_25), .cin(s_135_24), .o(t_3539), .co(t_3540), .cout(t_3541));
compressor_4_2 u2_1209(.a(s_135_33), .b(s_135_32), .c(s_135_31), .d(s_135_30), .cin(s_135_29), .o(t_3542), .co(t_3543), .cout(t_3544));
compressor_4_2 u2_1210(.a(s_135_38), .b(s_135_37), .c(s_135_36), .d(s_135_35), .cin(s_135_34), .o(t_3545), .co(t_3546), .cout(t_3547));
compressor_4_2 u2_1211(.a(s_135_43), .b(s_135_42), .c(s_135_41), .d(s_135_40), .cin(s_135_39), .o(t_3548), .co(t_3549), .cout(t_3550));
compressor_4_2 u2_1212(.a(s_135_48), .b(s_135_47), .c(s_135_46), .d(s_135_45), .cin(s_135_44), .o(t_3551), .co(t_3552), .cout(t_3553));
compressor_4_2 u2_1213(.a(s_135_53), .b(s_135_52), .c(s_135_51), .d(s_135_50), .cin(s_135_49), .o(t_3554), .co(t_3555), .cout(t_3556));
compressor_4_2 u2_1214(.a(s_135_58), .b(s_135_57), .c(s_135_56), .d(s_135_55), .cin(s_135_54), .o(t_3557), .co(t_3558), .cout(t_3559));
compressor_3_2 u1_1215(.a(s_135_61), .b(s_135_60), .cin(s_135_59), .o(t_3560), .cout(t_3561));
compressor_4_2 u2_1216(.a(s_136_2), .b(s_136_1), .c(s_136_0), .d(t_3517), .cin(t_3520), .o(t_3562), .co(t_3563), .cout(t_3564));
compressor_4_2 u2_1217(.a(s_136_5), .b(s_136_4), .c(s_136_3), .d(t_3523), .cin(t_3526), .o(t_3565), .co(t_3566), .cout(t_3567));
compressor_4_2 u2_1218(.a(s_136_8), .b(s_136_7), .c(s_136_6), .d(t_3529), .cin(t_3532), .o(t_3568), .co(t_3569), .cout(t_3570));
compressor_4_2 u2_1219(.a(s_136_11), .b(s_136_10), .c(s_136_9), .d(t_3535), .cin(t_3538), .o(t_3571), .co(t_3572), .cout(t_3573));
compressor_4_2 u2_1220(.a(s_136_14), .b(s_136_13), .c(s_136_12), .d(t_3541), .cin(t_3544), .o(t_3574), .co(t_3575), .cout(t_3576));
compressor_4_2 u2_1221(.a(s_136_17), .b(s_136_16), .c(s_136_15), .d(t_3547), .cin(t_3550), .o(t_3577), .co(t_3578), .cout(t_3579));
compressor_4_2 u2_1222(.a(s_136_20), .b(s_136_19), .c(s_136_18), .d(t_3553), .cin(t_3556), .o(t_3580), .co(t_3581), .cout(t_3582));
compressor_4_2 u2_1223(.a(s_136_23), .b(s_136_22), .c(s_136_21), .d(t_3559), .cin(t_3561), .o(t_3583), .co(t_3584), .cout(t_3585));
compressor_4_2 u2_1224(.a(s_136_28), .b(s_136_27), .c(s_136_26), .d(s_136_25), .cin(s_136_24), .o(t_3586), .co(t_3587), .cout(t_3588));
compressor_4_2 u2_1225(.a(s_136_33), .b(s_136_32), .c(s_136_31), .d(s_136_30), .cin(s_136_29), .o(t_3589), .co(t_3590), .cout(t_3591));
compressor_4_2 u2_1226(.a(s_136_38), .b(s_136_37), .c(s_136_36), .d(s_136_35), .cin(s_136_34), .o(t_3592), .co(t_3593), .cout(t_3594));
compressor_4_2 u2_1227(.a(s_136_43), .b(s_136_42), .c(s_136_41), .d(s_136_40), .cin(s_136_39), .o(t_3595), .co(t_3596), .cout(t_3597));
compressor_4_2 u2_1228(.a(s_136_48), .b(s_136_47), .c(s_136_46), .d(s_136_45), .cin(s_136_44), .o(t_3598), .co(t_3599), .cout(t_3600));
compressor_4_2 u2_1229(.a(s_136_53), .b(s_136_52), .c(s_136_51), .d(s_136_50), .cin(s_136_49), .o(t_3601), .co(t_3602), .cout(t_3603));
compressor_4_2 u2_1230(.a(s_136_58), .b(s_136_57), .c(s_136_56), .d(s_136_55), .cin(s_136_54), .o(t_3604), .co(t_3605), .cout(t_3606));
half_adder u0_1231(.a(s_136_60), .b(s_136_59), .o(t_3607), .cout(t_3608));
compressor_4_2 u2_1232(.a(s_137_2), .b(s_137_1), .c(s_137_0), .d(t_3564), .cin(t_3567), .o(t_3609), .co(t_3610), .cout(t_3611));
compressor_4_2 u2_1233(.a(s_137_5), .b(s_137_4), .c(s_137_3), .d(t_3570), .cin(t_3573), .o(t_3612), .co(t_3613), .cout(t_3614));
compressor_4_2 u2_1234(.a(s_137_8), .b(s_137_7), .c(s_137_6), .d(t_3576), .cin(t_3579), .o(t_3615), .co(t_3616), .cout(t_3617));
compressor_4_2 u2_1235(.a(s_137_11), .b(s_137_10), .c(s_137_9), .d(t_3582), .cin(t_3585), .o(t_3618), .co(t_3619), .cout(t_3620));
compressor_4_2 u2_1236(.a(s_137_14), .b(s_137_13), .c(s_137_12), .d(t_3588), .cin(t_3591), .o(t_3621), .co(t_3622), .cout(t_3623));
compressor_4_2 u2_1237(.a(s_137_17), .b(s_137_16), .c(s_137_15), .d(t_3594), .cin(t_3597), .o(t_3624), .co(t_3625), .cout(t_3626));
compressor_4_2 u2_1238(.a(s_137_20), .b(s_137_19), .c(s_137_18), .d(t_3600), .cin(t_3603), .o(t_3627), .co(t_3628), .cout(t_3629));
compressor_4_2 u2_1239(.a(s_137_23), .b(s_137_22), .c(s_137_21), .d(t_3606), .cin(t_3608), .o(t_3630), .co(t_3631), .cout(t_3632));
compressor_4_2 u2_1240(.a(s_137_28), .b(s_137_27), .c(s_137_26), .d(s_137_25), .cin(s_137_24), .o(t_3633), .co(t_3634), .cout(t_3635));
compressor_4_2 u2_1241(.a(s_137_33), .b(s_137_32), .c(s_137_31), .d(s_137_30), .cin(s_137_29), .o(t_3636), .co(t_3637), .cout(t_3638));
compressor_4_2 u2_1242(.a(s_137_38), .b(s_137_37), .c(s_137_36), .d(s_137_35), .cin(s_137_34), .o(t_3639), .co(t_3640), .cout(t_3641));
compressor_4_2 u2_1243(.a(s_137_43), .b(s_137_42), .c(s_137_41), .d(s_137_40), .cin(s_137_39), .o(t_3642), .co(t_3643), .cout(t_3644));
compressor_4_2 u2_1244(.a(s_137_48), .b(s_137_47), .c(s_137_46), .d(s_137_45), .cin(s_137_44), .o(t_3645), .co(t_3646), .cout(t_3647));
compressor_4_2 u2_1245(.a(s_137_53), .b(s_137_52), .c(s_137_51), .d(s_137_50), .cin(s_137_49), .o(t_3648), .co(t_3649), .cout(t_3650));
compressor_4_2 u2_1246(.a(s_137_58), .b(s_137_57), .c(s_137_56), .d(s_137_55), .cin(s_137_54), .o(t_3651), .co(t_3652), .cout(t_3653));
half_adder u0_1247(.a(s_137_60), .b(s_137_59), .o(t_3654), .cout(t_3655));
compressor_4_2 u2_1248(.a(s_138_2), .b(s_138_1), .c(s_138_0), .d(t_3611), .cin(t_3614), .o(t_3656), .co(t_3657), .cout(t_3658));
compressor_4_2 u2_1249(.a(s_138_5), .b(s_138_4), .c(s_138_3), .d(t_3617), .cin(t_3620), .o(t_3659), .co(t_3660), .cout(t_3661));
compressor_4_2 u2_1250(.a(s_138_8), .b(s_138_7), .c(s_138_6), .d(t_3623), .cin(t_3626), .o(t_3662), .co(t_3663), .cout(t_3664));
compressor_4_2 u2_1251(.a(s_138_11), .b(s_138_10), .c(s_138_9), .d(t_3629), .cin(t_3632), .o(t_3665), .co(t_3666), .cout(t_3667));
compressor_4_2 u2_1252(.a(s_138_14), .b(s_138_13), .c(s_138_12), .d(t_3635), .cin(t_3638), .o(t_3668), .co(t_3669), .cout(t_3670));
compressor_4_2 u2_1253(.a(s_138_17), .b(s_138_16), .c(s_138_15), .d(t_3641), .cin(t_3644), .o(t_3671), .co(t_3672), .cout(t_3673));
compressor_4_2 u2_1254(.a(s_138_20), .b(s_138_19), .c(s_138_18), .d(t_3647), .cin(t_3650), .o(t_3674), .co(t_3675), .cout(t_3676));
compressor_4_2 u2_1255(.a(s_138_23), .b(s_138_22), .c(s_138_21), .d(t_3653), .cin(t_3655), .o(t_3677), .co(t_3678), .cout(t_3679));
compressor_4_2 u2_1256(.a(s_138_28), .b(s_138_27), .c(s_138_26), .d(s_138_25), .cin(s_138_24), .o(t_3680), .co(t_3681), .cout(t_3682));
compressor_4_2 u2_1257(.a(s_138_33), .b(s_138_32), .c(s_138_31), .d(s_138_30), .cin(s_138_29), .o(t_3683), .co(t_3684), .cout(t_3685));
compressor_4_2 u2_1258(.a(s_138_38), .b(s_138_37), .c(s_138_36), .d(s_138_35), .cin(s_138_34), .o(t_3686), .co(t_3687), .cout(t_3688));
compressor_4_2 u2_1259(.a(s_138_43), .b(s_138_42), .c(s_138_41), .d(s_138_40), .cin(s_138_39), .o(t_3689), .co(t_3690), .cout(t_3691));
compressor_4_2 u2_1260(.a(s_138_48), .b(s_138_47), .c(s_138_46), .d(s_138_45), .cin(s_138_44), .o(t_3692), .co(t_3693), .cout(t_3694));
compressor_4_2 u2_1261(.a(s_138_53), .b(s_138_52), .c(s_138_51), .d(s_138_50), .cin(s_138_49), .o(t_3695), .co(t_3696), .cout(t_3697));
compressor_4_2 u2_1262(.a(s_138_58), .b(s_138_57), .c(s_138_56), .d(s_138_55), .cin(s_138_54), .o(t_3698), .co(t_3699), .cout(t_3700));
compressor_4_2 u2_1263(.a(s_139_2), .b(s_139_1), .c(s_139_0), .d(t_3658), .cin(t_3661), .o(t_3701), .co(t_3702), .cout(t_3703));
compressor_4_2 u2_1264(.a(s_139_5), .b(s_139_4), .c(s_139_3), .d(t_3664), .cin(t_3667), .o(t_3704), .co(t_3705), .cout(t_3706));
compressor_4_2 u2_1265(.a(s_139_8), .b(s_139_7), .c(s_139_6), .d(t_3670), .cin(t_3673), .o(t_3707), .co(t_3708), .cout(t_3709));
compressor_4_2 u2_1266(.a(s_139_11), .b(s_139_10), .c(s_139_9), .d(t_3676), .cin(t_3679), .o(t_3710), .co(t_3711), .cout(t_3712));
compressor_4_2 u2_1267(.a(s_139_14), .b(s_139_13), .c(s_139_12), .d(t_3682), .cin(t_3685), .o(t_3713), .co(t_3714), .cout(t_3715));
compressor_4_2 u2_1268(.a(s_139_17), .b(s_139_16), .c(s_139_15), .d(t_3688), .cin(t_3691), .o(t_3716), .co(t_3717), .cout(t_3718));
compressor_4_2 u2_1269(.a(s_139_20), .b(s_139_19), .c(s_139_18), .d(t_3694), .cin(t_3697), .o(t_3719), .co(t_3720), .cout(t_3721));
compressor_4_2 u2_1270(.a(s_139_24), .b(s_139_23), .c(s_139_22), .d(s_139_21), .cin(t_3700), .o(t_3722), .co(t_3723), .cout(t_3724));
compressor_4_2 u2_1271(.a(s_139_29), .b(s_139_28), .c(s_139_27), .d(s_139_26), .cin(s_139_25), .o(t_3725), .co(t_3726), .cout(t_3727));
compressor_4_2 u2_1272(.a(s_139_34), .b(s_139_33), .c(s_139_32), .d(s_139_31), .cin(s_139_30), .o(t_3728), .co(t_3729), .cout(t_3730));
compressor_4_2 u2_1273(.a(s_139_39), .b(s_139_38), .c(s_139_37), .d(s_139_36), .cin(s_139_35), .o(t_3731), .co(t_3732), .cout(t_3733));
compressor_4_2 u2_1274(.a(s_139_44), .b(s_139_43), .c(s_139_42), .d(s_139_41), .cin(s_139_40), .o(t_3734), .co(t_3735), .cout(t_3736));
compressor_4_2 u2_1275(.a(s_139_49), .b(s_139_48), .c(s_139_47), .d(s_139_46), .cin(s_139_45), .o(t_3737), .co(t_3738), .cout(t_3739));
compressor_4_2 u2_1276(.a(s_139_54), .b(s_139_53), .c(s_139_52), .d(s_139_51), .cin(s_139_50), .o(t_3740), .co(t_3741), .cout(t_3742));
compressor_4_2 u2_1277(.a(s_139_59), .b(s_139_58), .c(s_139_57), .d(s_139_56), .cin(s_139_55), .o(t_3743), .co(t_3744), .cout(t_3745));
compressor_4_2 u2_1278(.a(s_140_2), .b(s_140_1), .c(s_140_0), .d(t_3703), .cin(t_3706), .o(t_3746), .co(t_3747), .cout(t_3748));
compressor_4_2 u2_1279(.a(s_140_5), .b(s_140_4), .c(s_140_3), .d(t_3709), .cin(t_3712), .o(t_3749), .co(t_3750), .cout(t_3751));
compressor_4_2 u2_1280(.a(s_140_8), .b(s_140_7), .c(s_140_6), .d(t_3715), .cin(t_3718), .o(t_3752), .co(t_3753), .cout(t_3754));
compressor_4_2 u2_1281(.a(s_140_11), .b(s_140_10), .c(s_140_9), .d(t_3721), .cin(t_3724), .o(t_3755), .co(t_3756), .cout(t_3757));
compressor_4_2 u2_1282(.a(s_140_14), .b(s_140_13), .c(s_140_12), .d(t_3727), .cin(t_3730), .o(t_3758), .co(t_3759), .cout(t_3760));
compressor_4_2 u2_1283(.a(s_140_17), .b(s_140_16), .c(s_140_15), .d(t_3733), .cin(t_3736), .o(t_3761), .co(t_3762), .cout(t_3763));
compressor_4_2 u2_1284(.a(s_140_20), .b(s_140_19), .c(s_140_18), .d(t_3739), .cin(t_3742), .o(t_3764), .co(t_3765), .cout(t_3766));
compressor_4_2 u2_1285(.a(s_140_24), .b(s_140_23), .c(s_140_22), .d(s_140_21), .cin(t_3745), .o(t_3767), .co(t_3768), .cout(t_3769));
compressor_4_2 u2_1286(.a(s_140_29), .b(s_140_28), .c(s_140_27), .d(s_140_26), .cin(s_140_25), .o(t_3770), .co(t_3771), .cout(t_3772));
compressor_4_2 u2_1287(.a(s_140_34), .b(s_140_33), .c(s_140_32), .d(s_140_31), .cin(s_140_30), .o(t_3773), .co(t_3774), .cout(t_3775));
compressor_4_2 u2_1288(.a(s_140_39), .b(s_140_38), .c(s_140_37), .d(s_140_36), .cin(s_140_35), .o(t_3776), .co(t_3777), .cout(t_3778));
compressor_4_2 u2_1289(.a(s_140_44), .b(s_140_43), .c(s_140_42), .d(s_140_41), .cin(s_140_40), .o(t_3779), .co(t_3780), .cout(t_3781));
compressor_4_2 u2_1290(.a(s_140_49), .b(s_140_48), .c(s_140_47), .d(s_140_46), .cin(s_140_45), .o(t_3782), .co(t_3783), .cout(t_3784));
compressor_4_2 u2_1291(.a(s_140_54), .b(s_140_53), .c(s_140_52), .d(s_140_51), .cin(s_140_50), .o(t_3785), .co(t_3786), .cout(t_3787));
compressor_3_2 u1_1292(.a(s_140_57), .b(s_140_56), .cin(s_140_55), .o(t_3788), .cout(t_3789));
compressor_4_2 u2_1293(.a(s_141_2), .b(s_141_1), .c(s_141_0), .d(t_3748), .cin(t_3751), .o(t_3790), .co(t_3791), .cout(t_3792));
compressor_4_2 u2_1294(.a(s_141_5), .b(s_141_4), .c(s_141_3), .d(t_3754), .cin(t_3757), .o(t_3793), .co(t_3794), .cout(t_3795));
compressor_4_2 u2_1295(.a(s_141_8), .b(s_141_7), .c(s_141_6), .d(t_3760), .cin(t_3763), .o(t_3796), .co(t_3797), .cout(t_3798));
compressor_4_2 u2_1296(.a(s_141_11), .b(s_141_10), .c(s_141_9), .d(t_3766), .cin(t_3769), .o(t_3799), .co(t_3800), .cout(t_3801));
compressor_4_2 u2_1297(.a(s_141_14), .b(s_141_13), .c(s_141_12), .d(t_3772), .cin(t_3775), .o(t_3802), .co(t_3803), .cout(t_3804));
compressor_4_2 u2_1298(.a(s_141_17), .b(s_141_16), .c(s_141_15), .d(t_3778), .cin(t_3781), .o(t_3805), .co(t_3806), .cout(t_3807));
compressor_4_2 u2_1299(.a(s_141_20), .b(s_141_19), .c(s_141_18), .d(t_3784), .cin(t_3787), .o(t_3808), .co(t_3809), .cout(t_3810));
compressor_4_2 u2_1300(.a(s_141_24), .b(s_141_23), .c(s_141_22), .d(s_141_21), .cin(t_3789), .o(t_3811), .co(t_3812), .cout(t_3813));
compressor_4_2 u2_1301(.a(s_141_29), .b(s_141_28), .c(s_141_27), .d(s_141_26), .cin(s_141_25), .o(t_3814), .co(t_3815), .cout(t_3816));
compressor_4_2 u2_1302(.a(s_141_34), .b(s_141_33), .c(s_141_32), .d(s_141_31), .cin(s_141_30), .o(t_3817), .co(t_3818), .cout(t_3819));
compressor_4_2 u2_1303(.a(s_141_39), .b(s_141_38), .c(s_141_37), .d(s_141_36), .cin(s_141_35), .o(t_3820), .co(t_3821), .cout(t_3822));
compressor_4_2 u2_1304(.a(s_141_44), .b(s_141_43), .c(s_141_42), .d(s_141_41), .cin(s_141_40), .o(t_3823), .co(t_3824), .cout(t_3825));
compressor_4_2 u2_1305(.a(s_141_49), .b(s_141_48), .c(s_141_47), .d(s_141_46), .cin(s_141_45), .o(t_3826), .co(t_3827), .cout(t_3828));
compressor_4_2 u2_1306(.a(s_141_54), .b(s_141_53), .c(s_141_52), .d(s_141_51), .cin(s_141_50), .o(t_3829), .co(t_3830), .cout(t_3831));
compressor_3_2 u1_1307(.a(s_141_57), .b(s_141_56), .cin(s_141_55), .o(t_3832), .cout(t_3833));
compressor_4_2 u2_1308(.a(s_142_2), .b(s_142_1), .c(s_142_0), .d(t_3792), .cin(t_3795), .o(t_3834), .co(t_3835), .cout(t_3836));
compressor_4_2 u2_1309(.a(s_142_5), .b(s_142_4), .c(s_142_3), .d(t_3798), .cin(t_3801), .o(t_3837), .co(t_3838), .cout(t_3839));
compressor_4_2 u2_1310(.a(s_142_8), .b(s_142_7), .c(s_142_6), .d(t_3804), .cin(t_3807), .o(t_3840), .co(t_3841), .cout(t_3842));
compressor_4_2 u2_1311(.a(s_142_11), .b(s_142_10), .c(s_142_9), .d(t_3810), .cin(t_3813), .o(t_3843), .co(t_3844), .cout(t_3845));
compressor_4_2 u2_1312(.a(s_142_14), .b(s_142_13), .c(s_142_12), .d(t_3816), .cin(t_3819), .o(t_3846), .co(t_3847), .cout(t_3848));
compressor_4_2 u2_1313(.a(s_142_17), .b(s_142_16), .c(s_142_15), .d(t_3822), .cin(t_3825), .o(t_3849), .co(t_3850), .cout(t_3851));
compressor_4_2 u2_1314(.a(s_142_20), .b(s_142_19), .c(s_142_18), .d(t_3828), .cin(t_3831), .o(t_3852), .co(t_3853), .cout(t_3854));
compressor_4_2 u2_1315(.a(s_142_24), .b(s_142_23), .c(s_142_22), .d(s_142_21), .cin(t_3833), .o(t_3855), .co(t_3856), .cout(t_3857));
compressor_4_2 u2_1316(.a(s_142_29), .b(s_142_28), .c(s_142_27), .d(s_142_26), .cin(s_142_25), .o(t_3858), .co(t_3859), .cout(t_3860));
compressor_4_2 u2_1317(.a(s_142_34), .b(s_142_33), .c(s_142_32), .d(s_142_31), .cin(s_142_30), .o(t_3861), .co(t_3862), .cout(t_3863));
compressor_4_2 u2_1318(.a(s_142_39), .b(s_142_38), .c(s_142_37), .d(s_142_36), .cin(s_142_35), .o(t_3864), .co(t_3865), .cout(t_3866));
compressor_4_2 u2_1319(.a(s_142_44), .b(s_142_43), .c(s_142_42), .d(s_142_41), .cin(s_142_40), .o(t_3867), .co(t_3868), .cout(t_3869));
compressor_4_2 u2_1320(.a(s_142_49), .b(s_142_48), .c(s_142_47), .d(s_142_46), .cin(s_142_45), .o(t_3870), .co(t_3871), .cout(t_3872));
compressor_4_2 u2_1321(.a(s_142_54), .b(s_142_53), .c(s_142_52), .d(s_142_51), .cin(s_142_50), .o(t_3873), .co(t_3874), .cout(t_3875));
compressor_3_2 u1_1322(.a(s_142_57), .b(s_142_56), .cin(s_142_55), .o(t_3876), .cout(t_3877));
compressor_4_2 u2_1323(.a(s_143_2), .b(s_143_1), .c(s_143_0), .d(t_3836), .cin(t_3839), .o(t_3878), .co(t_3879), .cout(t_3880));
compressor_4_2 u2_1324(.a(s_143_5), .b(s_143_4), .c(s_143_3), .d(t_3842), .cin(t_3845), .o(t_3881), .co(t_3882), .cout(t_3883));
compressor_4_2 u2_1325(.a(s_143_8), .b(s_143_7), .c(s_143_6), .d(t_3848), .cin(t_3851), .o(t_3884), .co(t_3885), .cout(t_3886));
compressor_4_2 u2_1326(.a(s_143_11), .b(s_143_10), .c(s_143_9), .d(t_3854), .cin(t_3857), .o(t_3887), .co(t_3888), .cout(t_3889));
compressor_4_2 u2_1327(.a(s_143_14), .b(s_143_13), .c(s_143_12), .d(t_3860), .cin(t_3863), .o(t_3890), .co(t_3891), .cout(t_3892));
compressor_4_2 u2_1328(.a(s_143_17), .b(s_143_16), .c(s_143_15), .d(t_3866), .cin(t_3869), .o(t_3893), .co(t_3894), .cout(t_3895));
compressor_4_2 u2_1329(.a(s_143_20), .b(s_143_19), .c(s_143_18), .d(t_3872), .cin(t_3875), .o(t_3896), .co(t_3897), .cout(t_3898));
compressor_4_2 u2_1330(.a(s_143_24), .b(s_143_23), .c(s_143_22), .d(s_143_21), .cin(t_3877), .o(t_3899), .co(t_3900), .cout(t_3901));
compressor_4_2 u2_1331(.a(s_143_29), .b(s_143_28), .c(s_143_27), .d(s_143_26), .cin(s_143_25), .o(t_3902), .co(t_3903), .cout(t_3904));
compressor_4_2 u2_1332(.a(s_143_34), .b(s_143_33), .c(s_143_32), .d(s_143_31), .cin(s_143_30), .o(t_3905), .co(t_3906), .cout(t_3907));
compressor_4_2 u2_1333(.a(s_143_39), .b(s_143_38), .c(s_143_37), .d(s_143_36), .cin(s_143_35), .o(t_3908), .co(t_3909), .cout(t_3910));
compressor_4_2 u2_1334(.a(s_143_44), .b(s_143_43), .c(s_143_42), .d(s_143_41), .cin(s_143_40), .o(t_3911), .co(t_3912), .cout(t_3913));
compressor_4_2 u2_1335(.a(s_143_49), .b(s_143_48), .c(s_143_47), .d(s_143_46), .cin(s_143_45), .o(t_3914), .co(t_3915), .cout(t_3916));
compressor_4_2 u2_1336(.a(s_143_54), .b(s_143_53), .c(s_143_52), .d(s_143_51), .cin(s_143_50), .o(t_3917), .co(t_3918), .cout(t_3919));
compressor_3_2 u1_1337(.a(s_143_57), .b(s_143_56), .cin(s_143_55), .o(t_3920), .cout(t_3921));
compressor_4_2 u2_1338(.a(s_144_2), .b(s_144_1), .c(s_144_0), .d(t_3880), .cin(t_3883), .o(t_3922), .co(t_3923), .cout(t_3924));
compressor_4_2 u2_1339(.a(s_144_5), .b(s_144_4), .c(s_144_3), .d(t_3886), .cin(t_3889), .o(t_3925), .co(t_3926), .cout(t_3927));
compressor_4_2 u2_1340(.a(s_144_8), .b(s_144_7), .c(s_144_6), .d(t_3892), .cin(t_3895), .o(t_3928), .co(t_3929), .cout(t_3930));
compressor_4_2 u2_1341(.a(s_144_11), .b(s_144_10), .c(s_144_9), .d(t_3898), .cin(t_3901), .o(t_3931), .co(t_3932), .cout(t_3933));
compressor_4_2 u2_1342(.a(s_144_14), .b(s_144_13), .c(s_144_12), .d(t_3904), .cin(t_3907), .o(t_3934), .co(t_3935), .cout(t_3936));
compressor_4_2 u2_1343(.a(s_144_17), .b(s_144_16), .c(s_144_15), .d(t_3910), .cin(t_3913), .o(t_3937), .co(t_3938), .cout(t_3939));
compressor_4_2 u2_1344(.a(s_144_20), .b(s_144_19), .c(s_144_18), .d(t_3916), .cin(t_3919), .o(t_3940), .co(t_3941), .cout(t_3942));
compressor_4_2 u2_1345(.a(s_144_24), .b(s_144_23), .c(s_144_22), .d(s_144_21), .cin(t_3921), .o(t_3943), .co(t_3944), .cout(t_3945));
compressor_4_2 u2_1346(.a(s_144_29), .b(s_144_28), .c(s_144_27), .d(s_144_26), .cin(s_144_25), .o(t_3946), .co(t_3947), .cout(t_3948));
compressor_4_2 u2_1347(.a(s_144_34), .b(s_144_33), .c(s_144_32), .d(s_144_31), .cin(s_144_30), .o(t_3949), .co(t_3950), .cout(t_3951));
compressor_4_2 u2_1348(.a(s_144_39), .b(s_144_38), .c(s_144_37), .d(s_144_36), .cin(s_144_35), .o(t_3952), .co(t_3953), .cout(t_3954));
compressor_4_2 u2_1349(.a(s_144_44), .b(s_144_43), .c(s_144_42), .d(s_144_41), .cin(s_144_40), .o(t_3955), .co(t_3956), .cout(t_3957));
compressor_4_2 u2_1350(.a(s_144_49), .b(s_144_48), .c(s_144_47), .d(s_144_46), .cin(s_144_45), .o(t_3958), .co(t_3959), .cout(t_3960));
compressor_4_2 u2_1351(.a(s_144_54), .b(s_144_53), .c(s_144_52), .d(s_144_51), .cin(s_144_50), .o(t_3961), .co(t_3962), .cout(t_3963));
half_adder u0_1352(.a(s_144_56), .b(s_144_55), .o(t_3964), .cout(t_3965));
compressor_4_2 u2_1353(.a(s_145_2), .b(s_145_1), .c(s_145_0), .d(t_3924), .cin(t_3927), .o(t_3966), .co(t_3967), .cout(t_3968));
compressor_4_2 u2_1354(.a(s_145_5), .b(s_145_4), .c(s_145_3), .d(t_3930), .cin(t_3933), .o(t_3969), .co(t_3970), .cout(t_3971));
compressor_4_2 u2_1355(.a(s_145_8), .b(s_145_7), .c(s_145_6), .d(t_3936), .cin(t_3939), .o(t_3972), .co(t_3973), .cout(t_3974));
compressor_4_2 u2_1356(.a(s_145_11), .b(s_145_10), .c(s_145_9), .d(t_3942), .cin(t_3945), .o(t_3975), .co(t_3976), .cout(t_3977));
compressor_4_2 u2_1357(.a(s_145_14), .b(s_145_13), .c(s_145_12), .d(t_3948), .cin(t_3951), .o(t_3978), .co(t_3979), .cout(t_3980));
compressor_4_2 u2_1358(.a(s_145_17), .b(s_145_16), .c(s_145_15), .d(t_3954), .cin(t_3957), .o(t_3981), .co(t_3982), .cout(t_3983));
compressor_4_2 u2_1359(.a(s_145_20), .b(s_145_19), .c(s_145_18), .d(t_3960), .cin(t_3963), .o(t_3984), .co(t_3985), .cout(t_3986));
compressor_4_2 u2_1360(.a(s_145_24), .b(s_145_23), .c(s_145_22), .d(s_145_21), .cin(t_3965), .o(t_3987), .co(t_3988), .cout(t_3989));
compressor_4_2 u2_1361(.a(s_145_29), .b(s_145_28), .c(s_145_27), .d(s_145_26), .cin(s_145_25), .o(t_3990), .co(t_3991), .cout(t_3992));
compressor_4_2 u2_1362(.a(s_145_34), .b(s_145_33), .c(s_145_32), .d(s_145_31), .cin(s_145_30), .o(t_3993), .co(t_3994), .cout(t_3995));
compressor_4_2 u2_1363(.a(s_145_39), .b(s_145_38), .c(s_145_37), .d(s_145_36), .cin(s_145_35), .o(t_3996), .co(t_3997), .cout(t_3998));
compressor_4_2 u2_1364(.a(s_145_44), .b(s_145_43), .c(s_145_42), .d(s_145_41), .cin(s_145_40), .o(t_3999), .co(t_4000), .cout(t_4001));
compressor_4_2 u2_1365(.a(s_145_49), .b(s_145_48), .c(s_145_47), .d(s_145_46), .cin(s_145_45), .o(t_4002), .co(t_4003), .cout(t_4004));
compressor_4_2 u2_1366(.a(s_145_54), .b(s_145_53), .c(s_145_52), .d(s_145_51), .cin(s_145_50), .o(t_4005), .co(t_4006), .cout(t_4007));
half_adder u0_1367(.a(s_145_56), .b(s_145_55), .o(t_4008), .cout(t_4009));
compressor_4_2 u2_1368(.a(s_146_2), .b(s_146_1), .c(s_146_0), .d(t_3968), .cin(t_3971), .o(t_4010), .co(t_4011), .cout(t_4012));
compressor_4_2 u2_1369(.a(s_146_5), .b(s_146_4), .c(s_146_3), .d(t_3974), .cin(t_3977), .o(t_4013), .co(t_4014), .cout(t_4015));
compressor_4_2 u2_1370(.a(s_146_8), .b(s_146_7), .c(s_146_6), .d(t_3980), .cin(t_3983), .o(t_4016), .co(t_4017), .cout(t_4018));
compressor_4_2 u2_1371(.a(s_146_11), .b(s_146_10), .c(s_146_9), .d(t_3986), .cin(t_3989), .o(t_4019), .co(t_4020), .cout(t_4021));
compressor_4_2 u2_1372(.a(s_146_14), .b(s_146_13), .c(s_146_12), .d(t_3992), .cin(t_3995), .o(t_4022), .co(t_4023), .cout(t_4024));
compressor_4_2 u2_1373(.a(s_146_17), .b(s_146_16), .c(s_146_15), .d(t_3998), .cin(t_4001), .o(t_4025), .co(t_4026), .cout(t_4027));
compressor_4_2 u2_1374(.a(s_146_20), .b(s_146_19), .c(s_146_18), .d(t_4004), .cin(t_4007), .o(t_4028), .co(t_4029), .cout(t_4030));
compressor_4_2 u2_1375(.a(s_146_24), .b(s_146_23), .c(s_146_22), .d(s_146_21), .cin(t_4009), .o(t_4031), .co(t_4032), .cout(t_4033));
compressor_4_2 u2_1376(.a(s_146_29), .b(s_146_28), .c(s_146_27), .d(s_146_26), .cin(s_146_25), .o(t_4034), .co(t_4035), .cout(t_4036));
compressor_4_2 u2_1377(.a(s_146_34), .b(s_146_33), .c(s_146_32), .d(s_146_31), .cin(s_146_30), .o(t_4037), .co(t_4038), .cout(t_4039));
compressor_4_2 u2_1378(.a(s_146_39), .b(s_146_38), .c(s_146_37), .d(s_146_36), .cin(s_146_35), .o(t_4040), .co(t_4041), .cout(t_4042));
compressor_4_2 u2_1379(.a(s_146_44), .b(s_146_43), .c(s_146_42), .d(s_146_41), .cin(s_146_40), .o(t_4043), .co(t_4044), .cout(t_4045));
compressor_4_2 u2_1380(.a(s_146_49), .b(s_146_48), .c(s_146_47), .d(s_146_46), .cin(s_146_45), .o(t_4046), .co(t_4047), .cout(t_4048));
compressor_4_2 u2_1381(.a(s_146_54), .b(s_146_53), .c(s_146_52), .d(s_146_51), .cin(s_146_50), .o(t_4049), .co(t_4050), .cout(t_4051));
compressor_4_2 u2_1382(.a(s_147_2), .b(s_147_1), .c(s_147_0), .d(t_4012), .cin(t_4015), .o(t_4052), .co(t_4053), .cout(t_4054));
compressor_4_2 u2_1383(.a(s_147_5), .b(s_147_4), .c(s_147_3), .d(t_4018), .cin(t_4021), .o(t_4055), .co(t_4056), .cout(t_4057));
compressor_4_2 u2_1384(.a(s_147_8), .b(s_147_7), .c(s_147_6), .d(t_4024), .cin(t_4027), .o(t_4058), .co(t_4059), .cout(t_4060));
compressor_4_2 u2_1385(.a(s_147_11), .b(s_147_10), .c(s_147_9), .d(t_4030), .cin(t_4033), .o(t_4061), .co(t_4062), .cout(t_4063));
compressor_4_2 u2_1386(.a(s_147_14), .b(s_147_13), .c(s_147_12), .d(t_4036), .cin(t_4039), .o(t_4064), .co(t_4065), .cout(t_4066));
compressor_4_2 u2_1387(.a(s_147_17), .b(s_147_16), .c(s_147_15), .d(t_4042), .cin(t_4045), .o(t_4067), .co(t_4068), .cout(t_4069));
compressor_4_2 u2_1388(.a(s_147_20), .b(s_147_19), .c(s_147_18), .d(t_4048), .cin(t_4051), .o(t_4070), .co(t_4071), .cout(t_4072));
compressor_4_2 u2_1389(.a(s_147_25), .b(s_147_24), .c(s_147_23), .d(s_147_22), .cin(s_147_21), .o(t_4073), .co(t_4074), .cout(t_4075));
compressor_4_2 u2_1390(.a(s_147_30), .b(s_147_29), .c(s_147_28), .d(s_147_27), .cin(s_147_26), .o(t_4076), .co(t_4077), .cout(t_4078));
compressor_4_2 u2_1391(.a(s_147_35), .b(s_147_34), .c(s_147_33), .d(s_147_32), .cin(s_147_31), .o(t_4079), .co(t_4080), .cout(t_4081));
compressor_4_2 u2_1392(.a(s_147_40), .b(s_147_39), .c(s_147_38), .d(s_147_37), .cin(s_147_36), .o(t_4082), .co(t_4083), .cout(t_4084));
compressor_4_2 u2_1393(.a(s_147_45), .b(s_147_44), .c(s_147_43), .d(s_147_42), .cin(s_147_41), .o(t_4085), .co(t_4086), .cout(t_4087));
compressor_4_2 u2_1394(.a(s_147_50), .b(s_147_49), .c(s_147_48), .d(s_147_47), .cin(s_147_46), .o(t_4088), .co(t_4089), .cout(t_4090));
compressor_4_2 u2_1395(.a(s_147_55), .b(s_147_54), .c(s_147_53), .d(s_147_52), .cin(s_147_51), .o(t_4091), .co(t_4092), .cout(t_4093));
compressor_4_2 u2_1396(.a(s_148_2), .b(s_148_1), .c(s_148_0), .d(t_4054), .cin(t_4057), .o(t_4094), .co(t_4095), .cout(t_4096));
compressor_4_2 u2_1397(.a(s_148_5), .b(s_148_4), .c(s_148_3), .d(t_4060), .cin(t_4063), .o(t_4097), .co(t_4098), .cout(t_4099));
compressor_4_2 u2_1398(.a(s_148_8), .b(s_148_7), .c(s_148_6), .d(t_4066), .cin(t_4069), .o(t_4100), .co(t_4101), .cout(t_4102));
compressor_4_2 u2_1399(.a(s_148_11), .b(s_148_10), .c(s_148_9), .d(t_4072), .cin(t_4075), .o(t_4103), .co(t_4104), .cout(t_4105));
compressor_4_2 u2_1400(.a(s_148_14), .b(s_148_13), .c(s_148_12), .d(t_4078), .cin(t_4081), .o(t_4106), .co(t_4107), .cout(t_4108));
compressor_4_2 u2_1401(.a(s_148_17), .b(s_148_16), .c(s_148_15), .d(t_4084), .cin(t_4087), .o(t_4109), .co(t_4110), .cout(t_4111));
compressor_4_2 u2_1402(.a(s_148_20), .b(s_148_19), .c(s_148_18), .d(t_4090), .cin(t_4093), .o(t_4112), .co(t_4113), .cout(t_4114));
compressor_4_2 u2_1403(.a(s_148_25), .b(s_148_24), .c(s_148_23), .d(s_148_22), .cin(s_148_21), .o(t_4115), .co(t_4116), .cout(t_4117));
compressor_4_2 u2_1404(.a(s_148_30), .b(s_148_29), .c(s_148_28), .d(s_148_27), .cin(s_148_26), .o(t_4118), .co(t_4119), .cout(t_4120));
compressor_4_2 u2_1405(.a(s_148_35), .b(s_148_34), .c(s_148_33), .d(s_148_32), .cin(s_148_31), .o(t_4121), .co(t_4122), .cout(t_4123));
compressor_4_2 u2_1406(.a(s_148_40), .b(s_148_39), .c(s_148_38), .d(s_148_37), .cin(s_148_36), .o(t_4124), .co(t_4125), .cout(t_4126));
compressor_4_2 u2_1407(.a(s_148_45), .b(s_148_44), .c(s_148_43), .d(s_148_42), .cin(s_148_41), .o(t_4127), .co(t_4128), .cout(t_4129));
compressor_4_2 u2_1408(.a(s_148_50), .b(s_148_49), .c(s_148_48), .d(s_148_47), .cin(s_148_46), .o(t_4130), .co(t_4131), .cout(t_4132));
compressor_3_2 u1_1409(.a(s_148_53), .b(s_148_52), .cin(s_148_51), .o(t_4133), .cout(t_4134));
compressor_4_2 u2_1410(.a(s_149_2), .b(s_149_1), .c(s_149_0), .d(t_4096), .cin(t_4099), .o(t_4135), .co(t_4136), .cout(t_4137));
compressor_4_2 u2_1411(.a(s_149_5), .b(s_149_4), .c(s_149_3), .d(t_4102), .cin(t_4105), .o(t_4138), .co(t_4139), .cout(t_4140));
compressor_4_2 u2_1412(.a(s_149_8), .b(s_149_7), .c(s_149_6), .d(t_4108), .cin(t_4111), .o(t_4141), .co(t_4142), .cout(t_4143));
compressor_4_2 u2_1413(.a(s_149_11), .b(s_149_10), .c(s_149_9), .d(t_4114), .cin(t_4117), .o(t_4144), .co(t_4145), .cout(t_4146));
compressor_4_2 u2_1414(.a(s_149_14), .b(s_149_13), .c(s_149_12), .d(t_4120), .cin(t_4123), .o(t_4147), .co(t_4148), .cout(t_4149));
compressor_4_2 u2_1415(.a(s_149_17), .b(s_149_16), .c(s_149_15), .d(t_4126), .cin(t_4129), .o(t_4150), .co(t_4151), .cout(t_4152));
compressor_4_2 u2_1416(.a(s_149_20), .b(s_149_19), .c(s_149_18), .d(t_4132), .cin(t_4134), .o(t_4153), .co(t_4154), .cout(t_4155));
compressor_4_2 u2_1417(.a(s_149_25), .b(s_149_24), .c(s_149_23), .d(s_149_22), .cin(s_149_21), .o(t_4156), .co(t_4157), .cout(t_4158));
compressor_4_2 u2_1418(.a(s_149_30), .b(s_149_29), .c(s_149_28), .d(s_149_27), .cin(s_149_26), .o(t_4159), .co(t_4160), .cout(t_4161));
compressor_4_2 u2_1419(.a(s_149_35), .b(s_149_34), .c(s_149_33), .d(s_149_32), .cin(s_149_31), .o(t_4162), .co(t_4163), .cout(t_4164));
compressor_4_2 u2_1420(.a(s_149_40), .b(s_149_39), .c(s_149_38), .d(s_149_37), .cin(s_149_36), .o(t_4165), .co(t_4166), .cout(t_4167));
compressor_4_2 u2_1421(.a(s_149_45), .b(s_149_44), .c(s_149_43), .d(s_149_42), .cin(s_149_41), .o(t_4168), .co(t_4169), .cout(t_4170));
compressor_4_2 u2_1422(.a(s_149_50), .b(s_149_49), .c(s_149_48), .d(s_149_47), .cin(s_149_46), .o(t_4171), .co(t_4172), .cout(t_4173));
compressor_3_2 u1_1423(.a(s_149_53), .b(s_149_52), .cin(s_149_51), .o(t_4174), .cout(t_4175));
compressor_4_2 u2_1424(.a(s_150_2), .b(s_150_1), .c(s_150_0), .d(t_4137), .cin(t_4140), .o(t_4176), .co(t_4177), .cout(t_4178));
compressor_4_2 u2_1425(.a(s_150_5), .b(s_150_4), .c(s_150_3), .d(t_4143), .cin(t_4146), .o(t_4179), .co(t_4180), .cout(t_4181));
compressor_4_2 u2_1426(.a(s_150_8), .b(s_150_7), .c(s_150_6), .d(t_4149), .cin(t_4152), .o(t_4182), .co(t_4183), .cout(t_4184));
compressor_4_2 u2_1427(.a(s_150_11), .b(s_150_10), .c(s_150_9), .d(t_4155), .cin(t_4158), .o(t_4185), .co(t_4186), .cout(t_4187));
compressor_4_2 u2_1428(.a(s_150_14), .b(s_150_13), .c(s_150_12), .d(t_4161), .cin(t_4164), .o(t_4188), .co(t_4189), .cout(t_4190));
compressor_4_2 u2_1429(.a(s_150_17), .b(s_150_16), .c(s_150_15), .d(t_4167), .cin(t_4170), .o(t_4191), .co(t_4192), .cout(t_4193));
compressor_4_2 u2_1430(.a(s_150_20), .b(s_150_19), .c(s_150_18), .d(t_4173), .cin(t_4175), .o(t_4194), .co(t_4195), .cout(t_4196));
compressor_4_2 u2_1431(.a(s_150_25), .b(s_150_24), .c(s_150_23), .d(s_150_22), .cin(s_150_21), .o(t_4197), .co(t_4198), .cout(t_4199));
compressor_4_2 u2_1432(.a(s_150_30), .b(s_150_29), .c(s_150_28), .d(s_150_27), .cin(s_150_26), .o(t_4200), .co(t_4201), .cout(t_4202));
compressor_4_2 u2_1433(.a(s_150_35), .b(s_150_34), .c(s_150_33), .d(s_150_32), .cin(s_150_31), .o(t_4203), .co(t_4204), .cout(t_4205));
compressor_4_2 u2_1434(.a(s_150_40), .b(s_150_39), .c(s_150_38), .d(s_150_37), .cin(s_150_36), .o(t_4206), .co(t_4207), .cout(t_4208));
compressor_4_2 u2_1435(.a(s_150_45), .b(s_150_44), .c(s_150_43), .d(s_150_42), .cin(s_150_41), .o(t_4209), .co(t_4210), .cout(t_4211));
compressor_4_2 u2_1436(.a(s_150_50), .b(s_150_49), .c(s_150_48), .d(s_150_47), .cin(s_150_46), .o(t_4212), .co(t_4213), .cout(t_4214));
compressor_3_2 u1_1437(.a(s_150_53), .b(s_150_52), .cin(s_150_51), .o(t_4215), .cout(t_4216));
compressor_4_2 u2_1438(.a(s_151_2), .b(s_151_1), .c(s_151_0), .d(t_4178), .cin(t_4181), .o(t_4217), .co(t_4218), .cout(t_4219));
compressor_4_2 u2_1439(.a(s_151_5), .b(s_151_4), .c(s_151_3), .d(t_4184), .cin(t_4187), .o(t_4220), .co(t_4221), .cout(t_4222));
compressor_4_2 u2_1440(.a(s_151_8), .b(s_151_7), .c(s_151_6), .d(t_4190), .cin(t_4193), .o(t_4223), .co(t_4224), .cout(t_4225));
compressor_4_2 u2_1441(.a(s_151_11), .b(s_151_10), .c(s_151_9), .d(t_4196), .cin(t_4199), .o(t_4226), .co(t_4227), .cout(t_4228));
compressor_4_2 u2_1442(.a(s_151_14), .b(s_151_13), .c(s_151_12), .d(t_4202), .cin(t_4205), .o(t_4229), .co(t_4230), .cout(t_4231));
compressor_4_2 u2_1443(.a(s_151_17), .b(s_151_16), .c(s_151_15), .d(t_4208), .cin(t_4211), .o(t_4232), .co(t_4233), .cout(t_4234));
compressor_4_2 u2_1444(.a(s_151_20), .b(s_151_19), .c(s_151_18), .d(t_4214), .cin(t_4216), .o(t_4235), .co(t_4236), .cout(t_4237));
compressor_4_2 u2_1445(.a(s_151_25), .b(s_151_24), .c(s_151_23), .d(s_151_22), .cin(s_151_21), .o(t_4238), .co(t_4239), .cout(t_4240));
compressor_4_2 u2_1446(.a(s_151_30), .b(s_151_29), .c(s_151_28), .d(s_151_27), .cin(s_151_26), .o(t_4241), .co(t_4242), .cout(t_4243));
compressor_4_2 u2_1447(.a(s_151_35), .b(s_151_34), .c(s_151_33), .d(s_151_32), .cin(s_151_31), .o(t_4244), .co(t_4245), .cout(t_4246));
compressor_4_2 u2_1448(.a(s_151_40), .b(s_151_39), .c(s_151_38), .d(s_151_37), .cin(s_151_36), .o(t_4247), .co(t_4248), .cout(t_4249));
compressor_4_2 u2_1449(.a(s_151_45), .b(s_151_44), .c(s_151_43), .d(s_151_42), .cin(s_151_41), .o(t_4250), .co(t_4251), .cout(t_4252));
compressor_4_2 u2_1450(.a(s_151_50), .b(s_151_49), .c(s_151_48), .d(s_151_47), .cin(s_151_46), .o(t_4253), .co(t_4254), .cout(t_4255));
compressor_3_2 u1_1451(.a(s_151_53), .b(s_151_52), .cin(s_151_51), .o(t_4256), .cout(t_4257));
compressor_4_2 u2_1452(.a(s_152_2), .b(s_152_1), .c(s_152_0), .d(t_4219), .cin(t_4222), .o(t_4258), .co(t_4259), .cout(t_4260));
compressor_4_2 u2_1453(.a(s_152_5), .b(s_152_4), .c(s_152_3), .d(t_4225), .cin(t_4228), .o(t_4261), .co(t_4262), .cout(t_4263));
compressor_4_2 u2_1454(.a(s_152_8), .b(s_152_7), .c(s_152_6), .d(t_4231), .cin(t_4234), .o(t_4264), .co(t_4265), .cout(t_4266));
compressor_4_2 u2_1455(.a(s_152_11), .b(s_152_10), .c(s_152_9), .d(t_4237), .cin(t_4240), .o(t_4267), .co(t_4268), .cout(t_4269));
compressor_4_2 u2_1456(.a(s_152_14), .b(s_152_13), .c(s_152_12), .d(t_4243), .cin(t_4246), .o(t_4270), .co(t_4271), .cout(t_4272));
compressor_4_2 u2_1457(.a(s_152_17), .b(s_152_16), .c(s_152_15), .d(t_4249), .cin(t_4252), .o(t_4273), .co(t_4274), .cout(t_4275));
compressor_4_2 u2_1458(.a(s_152_20), .b(s_152_19), .c(s_152_18), .d(t_4255), .cin(t_4257), .o(t_4276), .co(t_4277), .cout(t_4278));
compressor_4_2 u2_1459(.a(s_152_25), .b(s_152_24), .c(s_152_23), .d(s_152_22), .cin(s_152_21), .o(t_4279), .co(t_4280), .cout(t_4281));
compressor_4_2 u2_1460(.a(s_152_30), .b(s_152_29), .c(s_152_28), .d(s_152_27), .cin(s_152_26), .o(t_4282), .co(t_4283), .cout(t_4284));
compressor_4_2 u2_1461(.a(s_152_35), .b(s_152_34), .c(s_152_33), .d(s_152_32), .cin(s_152_31), .o(t_4285), .co(t_4286), .cout(t_4287));
compressor_4_2 u2_1462(.a(s_152_40), .b(s_152_39), .c(s_152_38), .d(s_152_37), .cin(s_152_36), .o(t_4288), .co(t_4289), .cout(t_4290));
compressor_4_2 u2_1463(.a(s_152_45), .b(s_152_44), .c(s_152_43), .d(s_152_42), .cin(s_152_41), .o(t_4291), .co(t_4292), .cout(t_4293));
compressor_4_2 u2_1464(.a(s_152_50), .b(s_152_49), .c(s_152_48), .d(s_152_47), .cin(s_152_46), .o(t_4294), .co(t_4295), .cout(t_4296));
half_adder u0_1465(.a(s_152_52), .b(s_152_51), .o(t_4297), .cout(t_4298));
compressor_4_2 u2_1466(.a(s_153_2), .b(s_153_1), .c(s_153_0), .d(t_4260), .cin(t_4263), .o(t_4299), .co(t_4300), .cout(t_4301));
compressor_4_2 u2_1467(.a(s_153_5), .b(s_153_4), .c(s_153_3), .d(t_4266), .cin(t_4269), .o(t_4302), .co(t_4303), .cout(t_4304));
compressor_4_2 u2_1468(.a(s_153_8), .b(s_153_7), .c(s_153_6), .d(t_4272), .cin(t_4275), .o(t_4305), .co(t_4306), .cout(t_4307));
compressor_4_2 u2_1469(.a(s_153_11), .b(s_153_10), .c(s_153_9), .d(t_4278), .cin(t_4281), .o(t_4308), .co(t_4309), .cout(t_4310));
compressor_4_2 u2_1470(.a(s_153_14), .b(s_153_13), .c(s_153_12), .d(t_4284), .cin(t_4287), .o(t_4311), .co(t_4312), .cout(t_4313));
compressor_4_2 u2_1471(.a(s_153_17), .b(s_153_16), .c(s_153_15), .d(t_4290), .cin(t_4293), .o(t_4314), .co(t_4315), .cout(t_4316));
compressor_4_2 u2_1472(.a(s_153_20), .b(s_153_19), .c(s_153_18), .d(t_4296), .cin(t_4298), .o(t_4317), .co(t_4318), .cout(t_4319));
compressor_4_2 u2_1473(.a(s_153_25), .b(s_153_24), .c(s_153_23), .d(s_153_22), .cin(s_153_21), .o(t_4320), .co(t_4321), .cout(t_4322));
compressor_4_2 u2_1474(.a(s_153_30), .b(s_153_29), .c(s_153_28), .d(s_153_27), .cin(s_153_26), .o(t_4323), .co(t_4324), .cout(t_4325));
compressor_4_2 u2_1475(.a(s_153_35), .b(s_153_34), .c(s_153_33), .d(s_153_32), .cin(s_153_31), .o(t_4326), .co(t_4327), .cout(t_4328));
compressor_4_2 u2_1476(.a(s_153_40), .b(s_153_39), .c(s_153_38), .d(s_153_37), .cin(s_153_36), .o(t_4329), .co(t_4330), .cout(t_4331));
compressor_4_2 u2_1477(.a(s_153_45), .b(s_153_44), .c(s_153_43), .d(s_153_42), .cin(s_153_41), .o(t_4332), .co(t_4333), .cout(t_4334));
compressor_4_2 u2_1478(.a(s_153_50), .b(s_153_49), .c(s_153_48), .d(s_153_47), .cin(s_153_46), .o(t_4335), .co(t_4336), .cout(t_4337));
half_adder u0_1479(.a(s_153_52), .b(s_153_51), .o(t_4338), .cout(t_4339));
compressor_4_2 u2_1480(.a(s_154_2), .b(s_154_1), .c(s_154_0), .d(t_4301), .cin(t_4304), .o(t_4340), .co(t_4341), .cout(t_4342));
compressor_4_2 u2_1481(.a(s_154_5), .b(s_154_4), .c(s_154_3), .d(t_4307), .cin(t_4310), .o(t_4343), .co(t_4344), .cout(t_4345));
compressor_4_2 u2_1482(.a(s_154_8), .b(s_154_7), .c(s_154_6), .d(t_4313), .cin(t_4316), .o(t_4346), .co(t_4347), .cout(t_4348));
compressor_4_2 u2_1483(.a(s_154_11), .b(s_154_10), .c(s_154_9), .d(t_4319), .cin(t_4322), .o(t_4349), .co(t_4350), .cout(t_4351));
compressor_4_2 u2_1484(.a(s_154_14), .b(s_154_13), .c(s_154_12), .d(t_4325), .cin(t_4328), .o(t_4352), .co(t_4353), .cout(t_4354));
compressor_4_2 u2_1485(.a(s_154_17), .b(s_154_16), .c(s_154_15), .d(t_4331), .cin(t_4334), .o(t_4355), .co(t_4356), .cout(t_4357));
compressor_4_2 u2_1486(.a(s_154_20), .b(s_154_19), .c(s_154_18), .d(t_4337), .cin(t_4339), .o(t_4358), .co(t_4359), .cout(t_4360));
compressor_4_2 u2_1487(.a(s_154_25), .b(s_154_24), .c(s_154_23), .d(s_154_22), .cin(s_154_21), .o(t_4361), .co(t_4362), .cout(t_4363));
compressor_4_2 u2_1488(.a(s_154_30), .b(s_154_29), .c(s_154_28), .d(s_154_27), .cin(s_154_26), .o(t_4364), .co(t_4365), .cout(t_4366));
compressor_4_2 u2_1489(.a(s_154_35), .b(s_154_34), .c(s_154_33), .d(s_154_32), .cin(s_154_31), .o(t_4367), .co(t_4368), .cout(t_4369));
compressor_4_2 u2_1490(.a(s_154_40), .b(s_154_39), .c(s_154_38), .d(s_154_37), .cin(s_154_36), .o(t_4370), .co(t_4371), .cout(t_4372));
compressor_4_2 u2_1491(.a(s_154_45), .b(s_154_44), .c(s_154_43), .d(s_154_42), .cin(s_154_41), .o(t_4373), .co(t_4374), .cout(t_4375));
compressor_4_2 u2_1492(.a(s_154_50), .b(s_154_49), .c(s_154_48), .d(s_154_47), .cin(s_154_46), .o(t_4376), .co(t_4377), .cout(t_4378));
compressor_4_2 u2_1493(.a(s_155_2), .b(s_155_1), .c(s_155_0), .d(t_4342), .cin(t_4345), .o(t_4379), .co(t_4380), .cout(t_4381));
compressor_4_2 u2_1494(.a(s_155_5), .b(s_155_4), .c(s_155_3), .d(t_4348), .cin(t_4351), .o(t_4382), .co(t_4383), .cout(t_4384));
compressor_4_2 u2_1495(.a(s_155_8), .b(s_155_7), .c(s_155_6), .d(t_4354), .cin(t_4357), .o(t_4385), .co(t_4386), .cout(t_4387));
compressor_4_2 u2_1496(.a(s_155_11), .b(s_155_10), .c(s_155_9), .d(t_4360), .cin(t_4363), .o(t_4388), .co(t_4389), .cout(t_4390));
compressor_4_2 u2_1497(.a(s_155_14), .b(s_155_13), .c(s_155_12), .d(t_4366), .cin(t_4369), .o(t_4391), .co(t_4392), .cout(t_4393));
compressor_4_2 u2_1498(.a(s_155_17), .b(s_155_16), .c(s_155_15), .d(t_4372), .cin(t_4375), .o(t_4394), .co(t_4395), .cout(t_4396));
compressor_4_2 u2_1499(.a(s_155_21), .b(s_155_20), .c(s_155_19), .d(s_155_18), .cin(t_4378), .o(t_4397), .co(t_4398), .cout(t_4399));
compressor_4_2 u2_1500(.a(s_155_26), .b(s_155_25), .c(s_155_24), .d(s_155_23), .cin(s_155_22), .o(t_4400), .co(t_4401), .cout(t_4402));
compressor_4_2 u2_1501(.a(s_155_31), .b(s_155_30), .c(s_155_29), .d(s_155_28), .cin(s_155_27), .o(t_4403), .co(t_4404), .cout(t_4405));
compressor_4_2 u2_1502(.a(s_155_36), .b(s_155_35), .c(s_155_34), .d(s_155_33), .cin(s_155_32), .o(t_4406), .co(t_4407), .cout(t_4408));
compressor_4_2 u2_1503(.a(s_155_41), .b(s_155_40), .c(s_155_39), .d(s_155_38), .cin(s_155_37), .o(t_4409), .co(t_4410), .cout(t_4411));
compressor_4_2 u2_1504(.a(s_155_46), .b(s_155_45), .c(s_155_44), .d(s_155_43), .cin(s_155_42), .o(t_4412), .co(t_4413), .cout(t_4414));
compressor_4_2 u2_1505(.a(s_155_51), .b(s_155_50), .c(s_155_49), .d(s_155_48), .cin(s_155_47), .o(t_4415), .co(t_4416), .cout(t_4417));
compressor_4_2 u2_1506(.a(s_156_2), .b(s_156_1), .c(s_156_0), .d(t_4381), .cin(t_4384), .o(t_4418), .co(t_4419), .cout(t_4420));
compressor_4_2 u2_1507(.a(s_156_5), .b(s_156_4), .c(s_156_3), .d(t_4387), .cin(t_4390), .o(t_4421), .co(t_4422), .cout(t_4423));
compressor_4_2 u2_1508(.a(s_156_8), .b(s_156_7), .c(s_156_6), .d(t_4393), .cin(t_4396), .o(t_4424), .co(t_4425), .cout(t_4426));
compressor_4_2 u2_1509(.a(s_156_11), .b(s_156_10), .c(s_156_9), .d(t_4399), .cin(t_4402), .o(t_4427), .co(t_4428), .cout(t_4429));
compressor_4_2 u2_1510(.a(s_156_14), .b(s_156_13), .c(s_156_12), .d(t_4405), .cin(t_4408), .o(t_4430), .co(t_4431), .cout(t_4432));
compressor_4_2 u2_1511(.a(s_156_17), .b(s_156_16), .c(s_156_15), .d(t_4411), .cin(t_4414), .o(t_4433), .co(t_4434), .cout(t_4435));
compressor_4_2 u2_1512(.a(s_156_21), .b(s_156_20), .c(s_156_19), .d(s_156_18), .cin(t_4417), .o(t_4436), .co(t_4437), .cout(t_4438));
compressor_4_2 u2_1513(.a(s_156_26), .b(s_156_25), .c(s_156_24), .d(s_156_23), .cin(s_156_22), .o(t_4439), .co(t_4440), .cout(t_4441));
compressor_4_2 u2_1514(.a(s_156_31), .b(s_156_30), .c(s_156_29), .d(s_156_28), .cin(s_156_27), .o(t_4442), .co(t_4443), .cout(t_4444));
compressor_4_2 u2_1515(.a(s_156_36), .b(s_156_35), .c(s_156_34), .d(s_156_33), .cin(s_156_32), .o(t_4445), .co(t_4446), .cout(t_4447));
compressor_4_2 u2_1516(.a(s_156_41), .b(s_156_40), .c(s_156_39), .d(s_156_38), .cin(s_156_37), .o(t_4448), .co(t_4449), .cout(t_4450));
compressor_4_2 u2_1517(.a(s_156_46), .b(s_156_45), .c(s_156_44), .d(s_156_43), .cin(s_156_42), .o(t_4451), .co(t_4452), .cout(t_4453));
compressor_3_2 u1_1518(.a(s_156_49), .b(s_156_48), .cin(s_156_47), .o(t_4454), .cout(t_4455));
compressor_4_2 u2_1519(.a(s_157_2), .b(s_157_1), .c(s_157_0), .d(t_4420), .cin(t_4423), .o(t_4456), .co(t_4457), .cout(t_4458));
compressor_4_2 u2_1520(.a(s_157_5), .b(s_157_4), .c(s_157_3), .d(t_4426), .cin(t_4429), .o(t_4459), .co(t_4460), .cout(t_4461));
compressor_4_2 u2_1521(.a(s_157_8), .b(s_157_7), .c(s_157_6), .d(t_4432), .cin(t_4435), .o(t_4462), .co(t_4463), .cout(t_4464));
compressor_4_2 u2_1522(.a(s_157_11), .b(s_157_10), .c(s_157_9), .d(t_4438), .cin(t_4441), .o(t_4465), .co(t_4466), .cout(t_4467));
compressor_4_2 u2_1523(.a(s_157_14), .b(s_157_13), .c(s_157_12), .d(t_4444), .cin(t_4447), .o(t_4468), .co(t_4469), .cout(t_4470));
compressor_4_2 u2_1524(.a(s_157_17), .b(s_157_16), .c(s_157_15), .d(t_4450), .cin(t_4453), .o(t_4471), .co(t_4472), .cout(t_4473));
compressor_4_2 u2_1525(.a(s_157_21), .b(s_157_20), .c(s_157_19), .d(s_157_18), .cin(t_4455), .o(t_4474), .co(t_4475), .cout(t_4476));
compressor_4_2 u2_1526(.a(s_157_26), .b(s_157_25), .c(s_157_24), .d(s_157_23), .cin(s_157_22), .o(t_4477), .co(t_4478), .cout(t_4479));
compressor_4_2 u2_1527(.a(s_157_31), .b(s_157_30), .c(s_157_29), .d(s_157_28), .cin(s_157_27), .o(t_4480), .co(t_4481), .cout(t_4482));
compressor_4_2 u2_1528(.a(s_157_36), .b(s_157_35), .c(s_157_34), .d(s_157_33), .cin(s_157_32), .o(t_4483), .co(t_4484), .cout(t_4485));
compressor_4_2 u2_1529(.a(s_157_41), .b(s_157_40), .c(s_157_39), .d(s_157_38), .cin(s_157_37), .o(t_4486), .co(t_4487), .cout(t_4488));
compressor_4_2 u2_1530(.a(s_157_46), .b(s_157_45), .c(s_157_44), .d(s_157_43), .cin(s_157_42), .o(t_4489), .co(t_4490), .cout(t_4491));
compressor_3_2 u1_1531(.a(s_157_49), .b(s_157_48), .cin(s_157_47), .o(t_4492), .cout(t_4493));
compressor_4_2 u2_1532(.a(s_158_2), .b(s_158_1), .c(s_158_0), .d(t_4458), .cin(t_4461), .o(t_4494), .co(t_4495), .cout(t_4496));
compressor_4_2 u2_1533(.a(s_158_5), .b(s_158_4), .c(s_158_3), .d(t_4464), .cin(t_4467), .o(t_4497), .co(t_4498), .cout(t_4499));
compressor_4_2 u2_1534(.a(s_158_8), .b(s_158_7), .c(s_158_6), .d(t_4470), .cin(t_4473), .o(t_4500), .co(t_4501), .cout(t_4502));
compressor_4_2 u2_1535(.a(s_158_11), .b(s_158_10), .c(s_158_9), .d(t_4476), .cin(t_4479), .o(t_4503), .co(t_4504), .cout(t_4505));
compressor_4_2 u2_1536(.a(s_158_14), .b(s_158_13), .c(s_158_12), .d(t_4482), .cin(t_4485), .o(t_4506), .co(t_4507), .cout(t_4508));
compressor_4_2 u2_1537(.a(s_158_17), .b(s_158_16), .c(s_158_15), .d(t_4488), .cin(t_4491), .o(t_4509), .co(t_4510), .cout(t_4511));
compressor_4_2 u2_1538(.a(s_158_21), .b(s_158_20), .c(s_158_19), .d(s_158_18), .cin(t_4493), .o(t_4512), .co(t_4513), .cout(t_4514));
compressor_4_2 u2_1539(.a(s_158_26), .b(s_158_25), .c(s_158_24), .d(s_158_23), .cin(s_158_22), .o(t_4515), .co(t_4516), .cout(t_4517));
compressor_4_2 u2_1540(.a(s_158_31), .b(s_158_30), .c(s_158_29), .d(s_158_28), .cin(s_158_27), .o(t_4518), .co(t_4519), .cout(t_4520));
compressor_4_2 u2_1541(.a(s_158_36), .b(s_158_35), .c(s_158_34), .d(s_158_33), .cin(s_158_32), .o(t_4521), .co(t_4522), .cout(t_4523));
compressor_4_2 u2_1542(.a(s_158_41), .b(s_158_40), .c(s_158_39), .d(s_158_38), .cin(s_158_37), .o(t_4524), .co(t_4525), .cout(t_4526));
compressor_4_2 u2_1543(.a(s_158_46), .b(s_158_45), .c(s_158_44), .d(s_158_43), .cin(s_158_42), .o(t_4527), .co(t_4528), .cout(t_4529));
compressor_3_2 u1_1544(.a(s_158_49), .b(s_158_48), .cin(s_158_47), .o(t_4530), .cout(t_4531));
compressor_4_2 u2_1545(.a(s_159_2), .b(s_159_1), .c(s_159_0), .d(t_4496), .cin(t_4499), .o(t_4532), .co(t_4533), .cout(t_4534));
compressor_4_2 u2_1546(.a(s_159_5), .b(s_159_4), .c(s_159_3), .d(t_4502), .cin(t_4505), .o(t_4535), .co(t_4536), .cout(t_4537));
compressor_4_2 u2_1547(.a(s_159_8), .b(s_159_7), .c(s_159_6), .d(t_4508), .cin(t_4511), .o(t_4538), .co(t_4539), .cout(t_4540));
compressor_4_2 u2_1548(.a(s_159_11), .b(s_159_10), .c(s_159_9), .d(t_4514), .cin(t_4517), .o(t_4541), .co(t_4542), .cout(t_4543));
compressor_4_2 u2_1549(.a(s_159_14), .b(s_159_13), .c(s_159_12), .d(t_4520), .cin(t_4523), .o(t_4544), .co(t_4545), .cout(t_4546));
compressor_4_2 u2_1550(.a(s_159_17), .b(s_159_16), .c(s_159_15), .d(t_4526), .cin(t_4529), .o(t_4547), .co(t_4548), .cout(t_4549));
compressor_4_2 u2_1551(.a(s_159_21), .b(s_159_20), .c(s_159_19), .d(s_159_18), .cin(t_4531), .o(t_4550), .co(t_4551), .cout(t_4552));
compressor_4_2 u2_1552(.a(s_159_26), .b(s_159_25), .c(s_159_24), .d(s_159_23), .cin(s_159_22), .o(t_4553), .co(t_4554), .cout(t_4555));
compressor_4_2 u2_1553(.a(s_159_31), .b(s_159_30), .c(s_159_29), .d(s_159_28), .cin(s_159_27), .o(t_4556), .co(t_4557), .cout(t_4558));
compressor_4_2 u2_1554(.a(s_159_36), .b(s_159_35), .c(s_159_34), .d(s_159_33), .cin(s_159_32), .o(t_4559), .co(t_4560), .cout(t_4561));
compressor_4_2 u2_1555(.a(s_159_41), .b(s_159_40), .c(s_159_39), .d(s_159_38), .cin(s_159_37), .o(t_4562), .co(t_4563), .cout(t_4564));
compressor_4_2 u2_1556(.a(s_159_46), .b(s_159_45), .c(s_159_44), .d(s_159_43), .cin(s_159_42), .o(t_4565), .co(t_4566), .cout(t_4567));
compressor_3_2 u1_1557(.a(s_159_49), .b(s_159_48), .cin(s_159_47), .o(t_4568), .cout(t_4569));
compressor_4_2 u2_1558(.a(s_160_2), .b(s_160_1), .c(s_160_0), .d(t_4534), .cin(t_4537), .o(t_4570), .co(t_4571), .cout(t_4572));
compressor_4_2 u2_1559(.a(s_160_5), .b(s_160_4), .c(s_160_3), .d(t_4540), .cin(t_4543), .o(t_4573), .co(t_4574), .cout(t_4575));
compressor_4_2 u2_1560(.a(s_160_8), .b(s_160_7), .c(s_160_6), .d(t_4546), .cin(t_4549), .o(t_4576), .co(t_4577), .cout(t_4578));
compressor_4_2 u2_1561(.a(s_160_11), .b(s_160_10), .c(s_160_9), .d(t_4552), .cin(t_4555), .o(t_4579), .co(t_4580), .cout(t_4581));
compressor_4_2 u2_1562(.a(s_160_14), .b(s_160_13), .c(s_160_12), .d(t_4558), .cin(t_4561), .o(t_4582), .co(t_4583), .cout(t_4584));
compressor_4_2 u2_1563(.a(s_160_17), .b(s_160_16), .c(s_160_15), .d(t_4564), .cin(t_4567), .o(t_4585), .co(t_4586), .cout(t_4587));
compressor_4_2 u2_1564(.a(s_160_21), .b(s_160_20), .c(s_160_19), .d(s_160_18), .cin(t_4569), .o(t_4588), .co(t_4589), .cout(t_4590));
compressor_4_2 u2_1565(.a(s_160_26), .b(s_160_25), .c(s_160_24), .d(s_160_23), .cin(s_160_22), .o(t_4591), .co(t_4592), .cout(t_4593));
compressor_4_2 u2_1566(.a(s_160_31), .b(s_160_30), .c(s_160_29), .d(s_160_28), .cin(s_160_27), .o(t_4594), .co(t_4595), .cout(t_4596));
compressor_4_2 u2_1567(.a(s_160_36), .b(s_160_35), .c(s_160_34), .d(s_160_33), .cin(s_160_32), .o(t_4597), .co(t_4598), .cout(t_4599));
compressor_4_2 u2_1568(.a(s_160_41), .b(s_160_40), .c(s_160_39), .d(s_160_38), .cin(s_160_37), .o(t_4600), .co(t_4601), .cout(t_4602));
compressor_4_2 u2_1569(.a(s_160_46), .b(s_160_45), .c(s_160_44), .d(s_160_43), .cin(s_160_42), .o(t_4603), .co(t_4604), .cout(t_4605));
half_adder u0_1570(.a(s_160_48), .b(s_160_47), .o(t_4606), .cout(t_4607));
compressor_4_2 u2_1571(.a(s_161_2), .b(s_161_1), .c(s_161_0), .d(t_4572), .cin(t_4575), .o(t_4608), .co(t_4609), .cout(t_4610));
compressor_4_2 u2_1572(.a(s_161_5), .b(s_161_4), .c(s_161_3), .d(t_4578), .cin(t_4581), .o(t_4611), .co(t_4612), .cout(t_4613));
compressor_4_2 u2_1573(.a(s_161_8), .b(s_161_7), .c(s_161_6), .d(t_4584), .cin(t_4587), .o(t_4614), .co(t_4615), .cout(t_4616));
compressor_4_2 u2_1574(.a(s_161_11), .b(s_161_10), .c(s_161_9), .d(t_4590), .cin(t_4593), .o(t_4617), .co(t_4618), .cout(t_4619));
compressor_4_2 u2_1575(.a(s_161_14), .b(s_161_13), .c(s_161_12), .d(t_4596), .cin(t_4599), .o(t_4620), .co(t_4621), .cout(t_4622));
compressor_4_2 u2_1576(.a(s_161_17), .b(s_161_16), .c(s_161_15), .d(t_4602), .cin(t_4605), .o(t_4623), .co(t_4624), .cout(t_4625));
compressor_4_2 u2_1577(.a(s_161_21), .b(s_161_20), .c(s_161_19), .d(s_161_18), .cin(t_4607), .o(t_4626), .co(t_4627), .cout(t_4628));
compressor_4_2 u2_1578(.a(s_161_26), .b(s_161_25), .c(s_161_24), .d(s_161_23), .cin(s_161_22), .o(t_4629), .co(t_4630), .cout(t_4631));
compressor_4_2 u2_1579(.a(s_161_31), .b(s_161_30), .c(s_161_29), .d(s_161_28), .cin(s_161_27), .o(t_4632), .co(t_4633), .cout(t_4634));
compressor_4_2 u2_1580(.a(s_161_36), .b(s_161_35), .c(s_161_34), .d(s_161_33), .cin(s_161_32), .o(t_4635), .co(t_4636), .cout(t_4637));
compressor_4_2 u2_1581(.a(s_161_41), .b(s_161_40), .c(s_161_39), .d(s_161_38), .cin(s_161_37), .o(t_4638), .co(t_4639), .cout(t_4640));
compressor_4_2 u2_1582(.a(s_161_46), .b(s_161_45), .c(s_161_44), .d(s_161_43), .cin(s_161_42), .o(t_4641), .co(t_4642), .cout(t_4643));
half_adder u0_1583(.a(s_161_48), .b(s_161_47), .o(t_4644), .cout(t_4645));
compressor_4_2 u2_1584(.a(s_162_2), .b(s_162_1), .c(s_162_0), .d(t_4610), .cin(t_4613), .o(t_4646), .co(t_4647), .cout(t_4648));
compressor_4_2 u2_1585(.a(s_162_5), .b(s_162_4), .c(s_162_3), .d(t_4616), .cin(t_4619), .o(t_4649), .co(t_4650), .cout(t_4651));
compressor_4_2 u2_1586(.a(s_162_8), .b(s_162_7), .c(s_162_6), .d(t_4622), .cin(t_4625), .o(t_4652), .co(t_4653), .cout(t_4654));
compressor_4_2 u2_1587(.a(s_162_11), .b(s_162_10), .c(s_162_9), .d(t_4628), .cin(t_4631), .o(t_4655), .co(t_4656), .cout(t_4657));
compressor_4_2 u2_1588(.a(s_162_14), .b(s_162_13), .c(s_162_12), .d(t_4634), .cin(t_4637), .o(t_4658), .co(t_4659), .cout(t_4660));
compressor_4_2 u2_1589(.a(s_162_17), .b(s_162_16), .c(s_162_15), .d(t_4640), .cin(t_4643), .o(t_4661), .co(t_4662), .cout(t_4663));
compressor_4_2 u2_1590(.a(s_162_21), .b(s_162_20), .c(s_162_19), .d(s_162_18), .cin(t_4645), .o(t_4664), .co(t_4665), .cout(t_4666));
compressor_4_2 u2_1591(.a(s_162_26), .b(s_162_25), .c(s_162_24), .d(s_162_23), .cin(s_162_22), .o(t_4667), .co(t_4668), .cout(t_4669));
compressor_4_2 u2_1592(.a(s_162_31), .b(s_162_30), .c(s_162_29), .d(s_162_28), .cin(s_162_27), .o(t_4670), .co(t_4671), .cout(t_4672));
compressor_4_2 u2_1593(.a(s_162_36), .b(s_162_35), .c(s_162_34), .d(s_162_33), .cin(s_162_32), .o(t_4673), .co(t_4674), .cout(t_4675));
compressor_4_2 u2_1594(.a(s_162_41), .b(s_162_40), .c(s_162_39), .d(s_162_38), .cin(s_162_37), .o(t_4676), .co(t_4677), .cout(t_4678));
compressor_4_2 u2_1595(.a(s_162_46), .b(s_162_45), .c(s_162_44), .d(s_162_43), .cin(s_162_42), .o(t_4679), .co(t_4680), .cout(t_4681));
compressor_4_2 u2_1596(.a(s_163_2), .b(s_163_1), .c(s_163_0), .d(t_4648), .cin(t_4651), .o(t_4682), .co(t_4683), .cout(t_4684));
compressor_4_2 u2_1597(.a(s_163_5), .b(s_163_4), .c(s_163_3), .d(t_4654), .cin(t_4657), .o(t_4685), .co(t_4686), .cout(t_4687));
compressor_4_2 u2_1598(.a(s_163_8), .b(s_163_7), .c(s_163_6), .d(t_4660), .cin(t_4663), .o(t_4688), .co(t_4689), .cout(t_4690));
compressor_4_2 u2_1599(.a(s_163_11), .b(s_163_10), .c(s_163_9), .d(t_4666), .cin(t_4669), .o(t_4691), .co(t_4692), .cout(t_4693));
compressor_4_2 u2_1600(.a(s_163_14), .b(s_163_13), .c(s_163_12), .d(t_4672), .cin(t_4675), .o(t_4694), .co(t_4695), .cout(t_4696));
compressor_4_2 u2_1601(.a(s_163_17), .b(s_163_16), .c(s_163_15), .d(t_4678), .cin(t_4681), .o(t_4697), .co(t_4698), .cout(t_4699));
compressor_4_2 u2_1602(.a(s_163_22), .b(s_163_21), .c(s_163_20), .d(s_163_19), .cin(s_163_18), .o(t_4700), .co(t_4701), .cout(t_4702));
compressor_4_2 u2_1603(.a(s_163_27), .b(s_163_26), .c(s_163_25), .d(s_163_24), .cin(s_163_23), .o(t_4703), .co(t_4704), .cout(t_4705));
compressor_4_2 u2_1604(.a(s_163_32), .b(s_163_31), .c(s_163_30), .d(s_163_29), .cin(s_163_28), .o(t_4706), .co(t_4707), .cout(t_4708));
compressor_4_2 u2_1605(.a(s_163_37), .b(s_163_36), .c(s_163_35), .d(s_163_34), .cin(s_163_33), .o(t_4709), .co(t_4710), .cout(t_4711));
compressor_4_2 u2_1606(.a(s_163_42), .b(s_163_41), .c(s_163_40), .d(s_163_39), .cin(s_163_38), .o(t_4712), .co(t_4713), .cout(t_4714));
compressor_4_2 u2_1607(.a(s_163_47), .b(s_163_46), .c(s_163_45), .d(s_163_44), .cin(s_163_43), .o(t_4715), .co(t_4716), .cout(t_4717));
compressor_4_2 u2_1608(.a(s_164_2), .b(s_164_1), .c(s_164_0), .d(t_4684), .cin(t_4687), .o(t_4718), .co(t_4719), .cout(t_4720));
compressor_4_2 u2_1609(.a(s_164_5), .b(s_164_4), .c(s_164_3), .d(t_4690), .cin(t_4693), .o(t_4721), .co(t_4722), .cout(t_4723));
compressor_4_2 u2_1610(.a(s_164_8), .b(s_164_7), .c(s_164_6), .d(t_4696), .cin(t_4699), .o(t_4724), .co(t_4725), .cout(t_4726));
compressor_4_2 u2_1611(.a(s_164_11), .b(s_164_10), .c(s_164_9), .d(t_4702), .cin(t_4705), .o(t_4727), .co(t_4728), .cout(t_4729));
compressor_4_2 u2_1612(.a(s_164_14), .b(s_164_13), .c(s_164_12), .d(t_4708), .cin(t_4711), .o(t_4730), .co(t_4731), .cout(t_4732));
compressor_4_2 u2_1613(.a(s_164_17), .b(s_164_16), .c(s_164_15), .d(t_4714), .cin(t_4717), .o(t_4733), .co(t_4734), .cout(t_4735));
compressor_4_2 u2_1614(.a(s_164_22), .b(s_164_21), .c(s_164_20), .d(s_164_19), .cin(s_164_18), .o(t_4736), .co(t_4737), .cout(t_4738));
compressor_4_2 u2_1615(.a(s_164_27), .b(s_164_26), .c(s_164_25), .d(s_164_24), .cin(s_164_23), .o(t_4739), .co(t_4740), .cout(t_4741));
compressor_4_2 u2_1616(.a(s_164_32), .b(s_164_31), .c(s_164_30), .d(s_164_29), .cin(s_164_28), .o(t_4742), .co(t_4743), .cout(t_4744));
compressor_4_2 u2_1617(.a(s_164_37), .b(s_164_36), .c(s_164_35), .d(s_164_34), .cin(s_164_33), .o(t_4745), .co(t_4746), .cout(t_4747));
compressor_4_2 u2_1618(.a(s_164_42), .b(s_164_41), .c(s_164_40), .d(s_164_39), .cin(s_164_38), .o(t_4748), .co(t_4749), .cout(t_4750));
compressor_3_2 u1_1619(.a(s_164_45), .b(s_164_44), .cin(s_164_43), .o(t_4751), .cout(t_4752));
compressor_4_2 u2_1620(.a(s_165_2), .b(s_165_1), .c(s_165_0), .d(t_4720), .cin(t_4723), .o(t_4753), .co(t_4754), .cout(t_4755));
compressor_4_2 u2_1621(.a(s_165_5), .b(s_165_4), .c(s_165_3), .d(t_4726), .cin(t_4729), .o(t_4756), .co(t_4757), .cout(t_4758));
compressor_4_2 u2_1622(.a(s_165_8), .b(s_165_7), .c(s_165_6), .d(t_4732), .cin(t_4735), .o(t_4759), .co(t_4760), .cout(t_4761));
compressor_4_2 u2_1623(.a(s_165_11), .b(s_165_10), .c(s_165_9), .d(t_4738), .cin(t_4741), .o(t_4762), .co(t_4763), .cout(t_4764));
compressor_4_2 u2_1624(.a(s_165_14), .b(s_165_13), .c(s_165_12), .d(t_4744), .cin(t_4747), .o(t_4765), .co(t_4766), .cout(t_4767));
compressor_4_2 u2_1625(.a(s_165_17), .b(s_165_16), .c(s_165_15), .d(t_4750), .cin(t_4752), .o(t_4768), .co(t_4769), .cout(t_4770));
compressor_4_2 u2_1626(.a(s_165_22), .b(s_165_21), .c(s_165_20), .d(s_165_19), .cin(s_165_18), .o(t_4771), .co(t_4772), .cout(t_4773));
compressor_4_2 u2_1627(.a(s_165_27), .b(s_165_26), .c(s_165_25), .d(s_165_24), .cin(s_165_23), .o(t_4774), .co(t_4775), .cout(t_4776));
compressor_4_2 u2_1628(.a(s_165_32), .b(s_165_31), .c(s_165_30), .d(s_165_29), .cin(s_165_28), .o(t_4777), .co(t_4778), .cout(t_4779));
compressor_4_2 u2_1629(.a(s_165_37), .b(s_165_36), .c(s_165_35), .d(s_165_34), .cin(s_165_33), .o(t_4780), .co(t_4781), .cout(t_4782));
compressor_4_2 u2_1630(.a(s_165_42), .b(s_165_41), .c(s_165_40), .d(s_165_39), .cin(s_165_38), .o(t_4783), .co(t_4784), .cout(t_4785));
compressor_3_2 u1_1631(.a(s_165_45), .b(s_165_44), .cin(s_165_43), .o(t_4786), .cout(t_4787));
compressor_4_2 u2_1632(.a(s_166_2), .b(s_166_1), .c(s_166_0), .d(t_4755), .cin(t_4758), .o(t_4788), .co(t_4789), .cout(t_4790));
compressor_4_2 u2_1633(.a(s_166_5), .b(s_166_4), .c(s_166_3), .d(t_4761), .cin(t_4764), .o(t_4791), .co(t_4792), .cout(t_4793));
compressor_4_2 u2_1634(.a(s_166_8), .b(s_166_7), .c(s_166_6), .d(t_4767), .cin(t_4770), .o(t_4794), .co(t_4795), .cout(t_4796));
compressor_4_2 u2_1635(.a(s_166_11), .b(s_166_10), .c(s_166_9), .d(t_4773), .cin(t_4776), .o(t_4797), .co(t_4798), .cout(t_4799));
compressor_4_2 u2_1636(.a(s_166_14), .b(s_166_13), .c(s_166_12), .d(t_4779), .cin(t_4782), .o(t_4800), .co(t_4801), .cout(t_4802));
compressor_4_2 u2_1637(.a(s_166_17), .b(s_166_16), .c(s_166_15), .d(t_4785), .cin(t_4787), .o(t_4803), .co(t_4804), .cout(t_4805));
compressor_4_2 u2_1638(.a(s_166_22), .b(s_166_21), .c(s_166_20), .d(s_166_19), .cin(s_166_18), .o(t_4806), .co(t_4807), .cout(t_4808));
compressor_4_2 u2_1639(.a(s_166_27), .b(s_166_26), .c(s_166_25), .d(s_166_24), .cin(s_166_23), .o(t_4809), .co(t_4810), .cout(t_4811));
compressor_4_2 u2_1640(.a(s_166_32), .b(s_166_31), .c(s_166_30), .d(s_166_29), .cin(s_166_28), .o(t_4812), .co(t_4813), .cout(t_4814));
compressor_4_2 u2_1641(.a(s_166_37), .b(s_166_36), .c(s_166_35), .d(s_166_34), .cin(s_166_33), .o(t_4815), .co(t_4816), .cout(t_4817));
compressor_4_2 u2_1642(.a(s_166_42), .b(s_166_41), .c(s_166_40), .d(s_166_39), .cin(s_166_38), .o(t_4818), .co(t_4819), .cout(t_4820));
compressor_3_2 u1_1643(.a(s_166_45), .b(s_166_44), .cin(s_166_43), .o(t_4821), .cout(t_4822));
compressor_4_2 u2_1644(.a(s_167_2), .b(s_167_1), .c(s_167_0), .d(t_4790), .cin(t_4793), .o(t_4823), .co(t_4824), .cout(t_4825));
compressor_4_2 u2_1645(.a(s_167_5), .b(s_167_4), .c(s_167_3), .d(t_4796), .cin(t_4799), .o(t_4826), .co(t_4827), .cout(t_4828));
compressor_4_2 u2_1646(.a(s_167_8), .b(s_167_7), .c(s_167_6), .d(t_4802), .cin(t_4805), .o(t_4829), .co(t_4830), .cout(t_4831));
compressor_4_2 u2_1647(.a(s_167_11), .b(s_167_10), .c(s_167_9), .d(t_4808), .cin(t_4811), .o(t_4832), .co(t_4833), .cout(t_4834));
compressor_4_2 u2_1648(.a(s_167_14), .b(s_167_13), .c(s_167_12), .d(t_4814), .cin(t_4817), .o(t_4835), .co(t_4836), .cout(t_4837));
compressor_4_2 u2_1649(.a(s_167_17), .b(s_167_16), .c(s_167_15), .d(t_4820), .cin(t_4822), .o(t_4838), .co(t_4839), .cout(t_4840));
compressor_4_2 u2_1650(.a(s_167_22), .b(s_167_21), .c(s_167_20), .d(s_167_19), .cin(s_167_18), .o(t_4841), .co(t_4842), .cout(t_4843));
compressor_4_2 u2_1651(.a(s_167_27), .b(s_167_26), .c(s_167_25), .d(s_167_24), .cin(s_167_23), .o(t_4844), .co(t_4845), .cout(t_4846));
compressor_4_2 u2_1652(.a(s_167_32), .b(s_167_31), .c(s_167_30), .d(s_167_29), .cin(s_167_28), .o(t_4847), .co(t_4848), .cout(t_4849));
compressor_4_2 u2_1653(.a(s_167_37), .b(s_167_36), .c(s_167_35), .d(s_167_34), .cin(s_167_33), .o(t_4850), .co(t_4851), .cout(t_4852));
compressor_4_2 u2_1654(.a(s_167_42), .b(s_167_41), .c(s_167_40), .d(s_167_39), .cin(s_167_38), .o(t_4853), .co(t_4854), .cout(t_4855));
compressor_3_2 u1_1655(.a(s_167_45), .b(s_167_44), .cin(s_167_43), .o(t_4856), .cout(t_4857));
compressor_4_2 u2_1656(.a(s_168_2), .b(s_168_1), .c(s_168_0), .d(t_4825), .cin(t_4828), .o(t_4858), .co(t_4859), .cout(t_4860));
compressor_4_2 u2_1657(.a(s_168_5), .b(s_168_4), .c(s_168_3), .d(t_4831), .cin(t_4834), .o(t_4861), .co(t_4862), .cout(t_4863));
compressor_4_2 u2_1658(.a(s_168_8), .b(s_168_7), .c(s_168_6), .d(t_4837), .cin(t_4840), .o(t_4864), .co(t_4865), .cout(t_4866));
compressor_4_2 u2_1659(.a(s_168_11), .b(s_168_10), .c(s_168_9), .d(t_4843), .cin(t_4846), .o(t_4867), .co(t_4868), .cout(t_4869));
compressor_4_2 u2_1660(.a(s_168_14), .b(s_168_13), .c(s_168_12), .d(t_4849), .cin(t_4852), .o(t_4870), .co(t_4871), .cout(t_4872));
compressor_4_2 u2_1661(.a(s_168_17), .b(s_168_16), .c(s_168_15), .d(t_4855), .cin(t_4857), .o(t_4873), .co(t_4874), .cout(t_4875));
compressor_4_2 u2_1662(.a(s_168_22), .b(s_168_21), .c(s_168_20), .d(s_168_19), .cin(s_168_18), .o(t_4876), .co(t_4877), .cout(t_4878));
compressor_4_2 u2_1663(.a(s_168_27), .b(s_168_26), .c(s_168_25), .d(s_168_24), .cin(s_168_23), .o(t_4879), .co(t_4880), .cout(t_4881));
compressor_4_2 u2_1664(.a(s_168_32), .b(s_168_31), .c(s_168_30), .d(s_168_29), .cin(s_168_28), .o(t_4882), .co(t_4883), .cout(t_4884));
compressor_4_2 u2_1665(.a(s_168_37), .b(s_168_36), .c(s_168_35), .d(s_168_34), .cin(s_168_33), .o(t_4885), .co(t_4886), .cout(t_4887));
compressor_4_2 u2_1666(.a(s_168_42), .b(s_168_41), .c(s_168_40), .d(s_168_39), .cin(s_168_38), .o(t_4888), .co(t_4889), .cout(t_4890));
half_adder u0_1667(.a(s_168_44), .b(s_168_43), .o(t_4891), .cout(t_4892));
compressor_4_2 u2_1668(.a(s_169_2), .b(s_169_1), .c(s_169_0), .d(t_4860), .cin(t_4863), .o(t_4893), .co(t_4894), .cout(t_4895));
compressor_4_2 u2_1669(.a(s_169_5), .b(s_169_4), .c(s_169_3), .d(t_4866), .cin(t_4869), .o(t_4896), .co(t_4897), .cout(t_4898));
compressor_4_2 u2_1670(.a(s_169_8), .b(s_169_7), .c(s_169_6), .d(t_4872), .cin(t_4875), .o(t_4899), .co(t_4900), .cout(t_4901));
compressor_4_2 u2_1671(.a(s_169_11), .b(s_169_10), .c(s_169_9), .d(t_4878), .cin(t_4881), .o(t_4902), .co(t_4903), .cout(t_4904));
compressor_4_2 u2_1672(.a(s_169_14), .b(s_169_13), .c(s_169_12), .d(t_4884), .cin(t_4887), .o(t_4905), .co(t_4906), .cout(t_4907));
compressor_4_2 u2_1673(.a(s_169_17), .b(s_169_16), .c(s_169_15), .d(t_4890), .cin(t_4892), .o(t_4908), .co(t_4909), .cout(t_4910));
compressor_4_2 u2_1674(.a(s_169_22), .b(s_169_21), .c(s_169_20), .d(s_169_19), .cin(s_169_18), .o(t_4911), .co(t_4912), .cout(t_4913));
compressor_4_2 u2_1675(.a(s_169_27), .b(s_169_26), .c(s_169_25), .d(s_169_24), .cin(s_169_23), .o(t_4914), .co(t_4915), .cout(t_4916));
compressor_4_2 u2_1676(.a(s_169_32), .b(s_169_31), .c(s_169_30), .d(s_169_29), .cin(s_169_28), .o(t_4917), .co(t_4918), .cout(t_4919));
compressor_4_2 u2_1677(.a(s_169_37), .b(s_169_36), .c(s_169_35), .d(s_169_34), .cin(s_169_33), .o(t_4920), .co(t_4921), .cout(t_4922));
compressor_4_2 u2_1678(.a(s_169_42), .b(s_169_41), .c(s_169_40), .d(s_169_39), .cin(s_169_38), .o(t_4923), .co(t_4924), .cout(t_4925));
half_adder u0_1679(.a(s_169_44), .b(s_169_43), .o(t_4926), .cout(t_4927));
compressor_4_2 u2_1680(.a(s_170_2), .b(s_170_1), .c(s_170_0), .d(t_4895), .cin(t_4898), .o(t_4928), .co(t_4929), .cout(t_4930));
compressor_4_2 u2_1681(.a(s_170_5), .b(s_170_4), .c(s_170_3), .d(t_4901), .cin(t_4904), .o(t_4931), .co(t_4932), .cout(t_4933));
compressor_4_2 u2_1682(.a(s_170_8), .b(s_170_7), .c(s_170_6), .d(t_4907), .cin(t_4910), .o(t_4934), .co(t_4935), .cout(t_4936));
compressor_4_2 u2_1683(.a(s_170_11), .b(s_170_10), .c(s_170_9), .d(t_4913), .cin(t_4916), .o(t_4937), .co(t_4938), .cout(t_4939));
compressor_4_2 u2_1684(.a(s_170_14), .b(s_170_13), .c(s_170_12), .d(t_4919), .cin(t_4922), .o(t_4940), .co(t_4941), .cout(t_4942));
compressor_4_2 u2_1685(.a(s_170_17), .b(s_170_16), .c(s_170_15), .d(t_4925), .cin(t_4927), .o(t_4943), .co(t_4944), .cout(t_4945));
compressor_4_2 u2_1686(.a(s_170_22), .b(s_170_21), .c(s_170_20), .d(s_170_19), .cin(s_170_18), .o(t_4946), .co(t_4947), .cout(t_4948));
compressor_4_2 u2_1687(.a(s_170_27), .b(s_170_26), .c(s_170_25), .d(s_170_24), .cin(s_170_23), .o(t_4949), .co(t_4950), .cout(t_4951));
compressor_4_2 u2_1688(.a(s_170_32), .b(s_170_31), .c(s_170_30), .d(s_170_29), .cin(s_170_28), .o(t_4952), .co(t_4953), .cout(t_4954));
compressor_4_2 u2_1689(.a(s_170_37), .b(s_170_36), .c(s_170_35), .d(s_170_34), .cin(s_170_33), .o(t_4955), .co(t_4956), .cout(t_4957));
compressor_4_2 u2_1690(.a(s_170_42), .b(s_170_41), .c(s_170_40), .d(s_170_39), .cin(s_170_38), .o(t_4958), .co(t_4959), .cout(t_4960));
compressor_4_2 u2_1691(.a(s_171_2), .b(s_171_1), .c(s_171_0), .d(t_4930), .cin(t_4933), .o(t_4961), .co(t_4962), .cout(t_4963));
compressor_4_2 u2_1692(.a(s_171_5), .b(s_171_4), .c(s_171_3), .d(t_4936), .cin(t_4939), .o(t_4964), .co(t_4965), .cout(t_4966));
compressor_4_2 u2_1693(.a(s_171_8), .b(s_171_7), .c(s_171_6), .d(t_4942), .cin(t_4945), .o(t_4967), .co(t_4968), .cout(t_4969));
compressor_4_2 u2_1694(.a(s_171_11), .b(s_171_10), .c(s_171_9), .d(t_4948), .cin(t_4951), .o(t_4970), .co(t_4971), .cout(t_4972));
compressor_4_2 u2_1695(.a(s_171_14), .b(s_171_13), .c(s_171_12), .d(t_4954), .cin(t_4957), .o(t_4973), .co(t_4974), .cout(t_4975));
compressor_4_2 u2_1696(.a(s_171_18), .b(s_171_17), .c(s_171_16), .d(s_171_15), .cin(t_4960), .o(t_4976), .co(t_4977), .cout(t_4978));
compressor_4_2 u2_1697(.a(s_171_23), .b(s_171_22), .c(s_171_21), .d(s_171_20), .cin(s_171_19), .o(t_4979), .co(t_4980), .cout(t_4981));
compressor_4_2 u2_1698(.a(s_171_28), .b(s_171_27), .c(s_171_26), .d(s_171_25), .cin(s_171_24), .o(t_4982), .co(t_4983), .cout(t_4984));
compressor_4_2 u2_1699(.a(s_171_33), .b(s_171_32), .c(s_171_31), .d(s_171_30), .cin(s_171_29), .o(t_4985), .co(t_4986), .cout(t_4987));
compressor_4_2 u2_1700(.a(s_171_38), .b(s_171_37), .c(s_171_36), .d(s_171_35), .cin(s_171_34), .o(t_4988), .co(t_4989), .cout(t_4990));
compressor_4_2 u2_1701(.a(s_171_43), .b(s_171_42), .c(s_171_41), .d(s_171_40), .cin(s_171_39), .o(t_4991), .co(t_4992), .cout(t_4993));
compressor_4_2 u2_1702(.a(s_172_2), .b(s_172_1), .c(s_172_0), .d(t_4963), .cin(t_4966), .o(t_4994), .co(t_4995), .cout(t_4996));
compressor_4_2 u2_1703(.a(s_172_5), .b(s_172_4), .c(s_172_3), .d(t_4969), .cin(t_4972), .o(t_4997), .co(t_4998), .cout(t_4999));
compressor_4_2 u2_1704(.a(s_172_8), .b(s_172_7), .c(s_172_6), .d(t_4975), .cin(t_4978), .o(t_5000), .co(t_5001), .cout(t_5002));
compressor_4_2 u2_1705(.a(s_172_11), .b(s_172_10), .c(s_172_9), .d(t_4981), .cin(t_4984), .o(t_5003), .co(t_5004), .cout(t_5005));
compressor_4_2 u2_1706(.a(s_172_14), .b(s_172_13), .c(s_172_12), .d(t_4987), .cin(t_4990), .o(t_5006), .co(t_5007), .cout(t_5008));
compressor_4_2 u2_1707(.a(s_172_18), .b(s_172_17), .c(s_172_16), .d(s_172_15), .cin(t_4993), .o(t_5009), .co(t_5010), .cout(t_5011));
compressor_4_2 u2_1708(.a(s_172_23), .b(s_172_22), .c(s_172_21), .d(s_172_20), .cin(s_172_19), .o(t_5012), .co(t_5013), .cout(t_5014));
compressor_4_2 u2_1709(.a(s_172_28), .b(s_172_27), .c(s_172_26), .d(s_172_25), .cin(s_172_24), .o(t_5015), .co(t_5016), .cout(t_5017));
compressor_4_2 u2_1710(.a(s_172_33), .b(s_172_32), .c(s_172_31), .d(s_172_30), .cin(s_172_29), .o(t_5018), .co(t_5019), .cout(t_5020));
compressor_4_2 u2_1711(.a(s_172_38), .b(s_172_37), .c(s_172_36), .d(s_172_35), .cin(s_172_34), .o(t_5021), .co(t_5022), .cout(t_5023));
compressor_3_2 u1_1712(.a(s_172_41), .b(s_172_40), .cin(s_172_39), .o(t_5024), .cout(t_5025));
compressor_4_2 u2_1713(.a(s_173_2), .b(s_173_1), .c(s_173_0), .d(t_4996), .cin(t_4999), .o(t_5026), .co(t_5027), .cout(t_5028));
compressor_4_2 u2_1714(.a(s_173_5), .b(s_173_4), .c(s_173_3), .d(t_5002), .cin(t_5005), .o(t_5029), .co(t_5030), .cout(t_5031));
compressor_4_2 u2_1715(.a(s_173_8), .b(s_173_7), .c(s_173_6), .d(t_5008), .cin(t_5011), .o(t_5032), .co(t_5033), .cout(t_5034));
compressor_4_2 u2_1716(.a(s_173_11), .b(s_173_10), .c(s_173_9), .d(t_5014), .cin(t_5017), .o(t_5035), .co(t_5036), .cout(t_5037));
compressor_4_2 u2_1717(.a(s_173_14), .b(s_173_13), .c(s_173_12), .d(t_5020), .cin(t_5023), .o(t_5038), .co(t_5039), .cout(t_5040));
compressor_4_2 u2_1718(.a(s_173_18), .b(s_173_17), .c(s_173_16), .d(s_173_15), .cin(t_5025), .o(t_5041), .co(t_5042), .cout(t_5043));
compressor_4_2 u2_1719(.a(s_173_23), .b(s_173_22), .c(s_173_21), .d(s_173_20), .cin(s_173_19), .o(t_5044), .co(t_5045), .cout(t_5046));
compressor_4_2 u2_1720(.a(s_173_28), .b(s_173_27), .c(s_173_26), .d(s_173_25), .cin(s_173_24), .o(t_5047), .co(t_5048), .cout(t_5049));
compressor_4_2 u2_1721(.a(s_173_33), .b(s_173_32), .c(s_173_31), .d(s_173_30), .cin(s_173_29), .o(t_5050), .co(t_5051), .cout(t_5052));
compressor_4_2 u2_1722(.a(s_173_38), .b(s_173_37), .c(s_173_36), .d(s_173_35), .cin(s_173_34), .o(t_5053), .co(t_5054), .cout(t_5055));
compressor_3_2 u1_1723(.a(s_173_41), .b(s_173_40), .cin(s_173_39), .o(t_5056), .cout(t_5057));
compressor_4_2 u2_1724(.a(s_174_2), .b(s_174_1), .c(s_174_0), .d(t_5028), .cin(t_5031), .o(t_5058), .co(t_5059), .cout(t_5060));
compressor_4_2 u2_1725(.a(s_174_5), .b(s_174_4), .c(s_174_3), .d(t_5034), .cin(t_5037), .o(t_5061), .co(t_5062), .cout(t_5063));
compressor_4_2 u2_1726(.a(s_174_8), .b(s_174_7), .c(s_174_6), .d(t_5040), .cin(t_5043), .o(t_5064), .co(t_5065), .cout(t_5066));
compressor_4_2 u2_1727(.a(s_174_11), .b(s_174_10), .c(s_174_9), .d(t_5046), .cin(t_5049), .o(t_5067), .co(t_5068), .cout(t_5069));
compressor_4_2 u2_1728(.a(s_174_14), .b(s_174_13), .c(s_174_12), .d(t_5052), .cin(t_5055), .o(t_5070), .co(t_5071), .cout(t_5072));
compressor_4_2 u2_1729(.a(s_174_18), .b(s_174_17), .c(s_174_16), .d(s_174_15), .cin(t_5057), .o(t_5073), .co(t_5074), .cout(t_5075));
compressor_4_2 u2_1730(.a(s_174_23), .b(s_174_22), .c(s_174_21), .d(s_174_20), .cin(s_174_19), .o(t_5076), .co(t_5077), .cout(t_5078));
compressor_4_2 u2_1731(.a(s_174_28), .b(s_174_27), .c(s_174_26), .d(s_174_25), .cin(s_174_24), .o(t_5079), .co(t_5080), .cout(t_5081));
compressor_4_2 u2_1732(.a(s_174_33), .b(s_174_32), .c(s_174_31), .d(s_174_30), .cin(s_174_29), .o(t_5082), .co(t_5083), .cout(t_5084));
compressor_4_2 u2_1733(.a(s_174_38), .b(s_174_37), .c(s_174_36), .d(s_174_35), .cin(s_174_34), .o(t_5085), .co(t_5086), .cout(t_5087));
compressor_3_2 u1_1734(.a(s_174_41), .b(s_174_40), .cin(s_174_39), .o(t_5088), .cout(t_5089));
compressor_4_2 u2_1735(.a(s_175_2), .b(s_175_1), .c(s_175_0), .d(t_5060), .cin(t_5063), .o(t_5090), .co(t_5091), .cout(t_5092));
compressor_4_2 u2_1736(.a(s_175_5), .b(s_175_4), .c(s_175_3), .d(t_5066), .cin(t_5069), .o(t_5093), .co(t_5094), .cout(t_5095));
compressor_4_2 u2_1737(.a(s_175_8), .b(s_175_7), .c(s_175_6), .d(t_5072), .cin(t_5075), .o(t_5096), .co(t_5097), .cout(t_5098));
compressor_4_2 u2_1738(.a(s_175_11), .b(s_175_10), .c(s_175_9), .d(t_5078), .cin(t_5081), .o(t_5099), .co(t_5100), .cout(t_5101));
compressor_4_2 u2_1739(.a(s_175_14), .b(s_175_13), .c(s_175_12), .d(t_5084), .cin(t_5087), .o(t_5102), .co(t_5103), .cout(t_5104));
compressor_4_2 u2_1740(.a(s_175_18), .b(s_175_17), .c(s_175_16), .d(s_175_15), .cin(t_5089), .o(t_5105), .co(t_5106), .cout(t_5107));
compressor_4_2 u2_1741(.a(s_175_23), .b(s_175_22), .c(s_175_21), .d(s_175_20), .cin(s_175_19), .o(t_5108), .co(t_5109), .cout(t_5110));
compressor_4_2 u2_1742(.a(s_175_28), .b(s_175_27), .c(s_175_26), .d(s_175_25), .cin(s_175_24), .o(t_5111), .co(t_5112), .cout(t_5113));
compressor_4_2 u2_1743(.a(s_175_33), .b(s_175_32), .c(s_175_31), .d(s_175_30), .cin(s_175_29), .o(t_5114), .co(t_5115), .cout(t_5116));
compressor_4_2 u2_1744(.a(s_175_38), .b(s_175_37), .c(s_175_36), .d(s_175_35), .cin(s_175_34), .o(t_5117), .co(t_5118), .cout(t_5119));
compressor_3_2 u1_1745(.a(s_175_41), .b(s_175_40), .cin(s_175_39), .o(t_5120), .cout(t_5121));
compressor_4_2 u2_1746(.a(s_176_2), .b(s_176_1), .c(s_176_0), .d(t_5092), .cin(t_5095), .o(t_5122), .co(t_5123), .cout(t_5124));
compressor_4_2 u2_1747(.a(s_176_5), .b(s_176_4), .c(s_176_3), .d(t_5098), .cin(t_5101), .o(t_5125), .co(t_5126), .cout(t_5127));
compressor_4_2 u2_1748(.a(s_176_8), .b(s_176_7), .c(s_176_6), .d(t_5104), .cin(t_5107), .o(t_5128), .co(t_5129), .cout(t_5130));
compressor_4_2 u2_1749(.a(s_176_11), .b(s_176_10), .c(s_176_9), .d(t_5110), .cin(t_5113), .o(t_5131), .co(t_5132), .cout(t_5133));
compressor_4_2 u2_1750(.a(s_176_14), .b(s_176_13), .c(s_176_12), .d(t_5116), .cin(t_5119), .o(t_5134), .co(t_5135), .cout(t_5136));
compressor_4_2 u2_1751(.a(s_176_18), .b(s_176_17), .c(s_176_16), .d(s_176_15), .cin(t_5121), .o(t_5137), .co(t_5138), .cout(t_5139));
compressor_4_2 u2_1752(.a(s_176_23), .b(s_176_22), .c(s_176_21), .d(s_176_20), .cin(s_176_19), .o(t_5140), .co(t_5141), .cout(t_5142));
compressor_4_2 u2_1753(.a(s_176_28), .b(s_176_27), .c(s_176_26), .d(s_176_25), .cin(s_176_24), .o(t_5143), .co(t_5144), .cout(t_5145));
compressor_4_2 u2_1754(.a(s_176_33), .b(s_176_32), .c(s_176_31), .d(s_176_30), .cin(s_176_29), .o(t_5146), .co(t_5147), .cout(t_5148));
compressor_4_2 u2_1755(.a(s_176_38), .b(s_176_37), .c(s_176_36), .d(s_176_35), .cin(s_176_34), .o(t_5149), .co(t_5150), .cout(t_5151));
half_adder u0_1756(.a(s_176_40), .b(s_176_39), .o(t_5152), .cout(t_5153));
compressor_4_2 u2_1757(.a(s_177_2), .b(s_177_1), .c(s_177_0), .d(t_5124), .cin(t_5127), .o(t_5154), .co(t_5155), .cout(t_5156));
compressor_4_2 u2_1758(.a(s_177_5), .b(s_177_4), .c(s_177_3), .d(t_5130), .cin(t_5133), .o(t_5157), .co(t_5158), .cout(t_5159));
compressor_4_2 u2_1759(.a(s_177_8), .b(s_177_7), .c(s_177_6), .d(t_5136), .cin(t_5139), .o(t_5160), .co(t_5161), .cout(t_5162));
compressor_4_2 u2_1760(.a(s_177_11), .b(s_177_10), .c(s_177_9), .d(t_5142), .cin(t_5145), .o(t_5163), .co(t_5164), .cout(t_5165));
compressor_4_2 u2_1761(.a(s_177_14), .b(s_177_13), .c(s_177_12), .d(t_5148), .cin(t_5151), .o(t_5166), .co(t_5167), .cout(t_5168));
compressor_4_2 u2_1762(.a(s_177_18), .b(s_177_17), .c(s_177_16), .d(s_177_15), .cin(t_5153), .o(t_5169), .co(t_5170), .cout(t_5171));
compressor_4_2 u2_1763(.a(s_177_23), .b(s_177_22), .c(s_177_21), .d(s_177_20), .cin(s_177_19), .o(t_5172), .co(t_5173), .cout(t_5174));
compressor_4_2 u2_1764(.a(s_177_28), .b(s_177_27), .c(s_177_26), .d(s_177_25), .cin(s_177_24), .o(t_5175), .co(t_5176), .cout(t_5177));
compressor_4_2 u2_1765(.a(s_177_33), .b(s_177_32), .c(s_177_31), .d(s_177_30), .cin(s_177_29), .o(t_5178), .co(t_5179), .cout(t_5180));
compressor_4_2 u2_1766(.a(s_177_38), .b(s_177_37), .c(s_177_36), .d(s_177_35), .cin(s_177_34), .o(t_5181), .co(t_5182), .cout(t_5183));
half_adder u0_1767(.a(s_177_40), .b(s_177_39), .o(t_5184), .cout(t_5185));
compressor_4_2 u2_1768(.a(s_178_2), .b(s_178_1), .c(s_178_0), .d(t_5156), .cin(t_5159), .o(t_5186), .co(t_5187), .cout(t_5188));
compressor_4_2 u2_1769(.a(s_178_5), .b(s_178_4), .c(s_178_3), .d(t_5162), .cin(t_5165), .o(t_5189), .co(t_5190), .cout(t_5191));
compressor_4_2 u2_1770(.a(s_178_8), .b(s_178_7), .c(s_178_6), .d(t_5168), .cin(t_5171), .o(t_5192), .co(t_5193), .cout(t_5194));
compressor_4_2 u2_1771(.a(s_178_11), .b(s_178_10), .c(s_178_9), .d(t_5174), .cin(t_5177), .o(t_5195), .co(t_5196), .cout(t_5197));
compressor_4_2 u2_1772(.a(s_178_14), .b(s_178_13), .c(s_178_12), .d(t_5180), .cin(t_5183), .o(t_5198), .co(t_5199), .cout(t_5200));
compressor_4_2 u2_1773(.a(s_178_18), .b(s_178_17), .c(s_178_16), .d(s_178_15), .cin(t_5185), .o(t_5201), .co(t_5202), .cout(t_5203));
compressor_4_2 u2_1774(.a(s_178_23), .b(s_178_22), .c(s_178_21), .d(s_178_20), .cin(s_178_19), .o(t_5204), .co(t_5205), .cout(t_5206));
compressor_4_2 u2_1775(.a(s_178_28), .b(s_178_27), .c(s_178_26), .d(s_178_25), .cin(s_178_24), .o(t_5207), .co(t_5208), .cout(t_5209));
compressor_4_2 u2_1776(.a(s_178_33), .b(s_178_32), .c(s_178_31), .d(s_178_30), .cin(s_178_29), .o(t_5210), .co(t_5211), .cout(t_5212));
compressor_4_2 u2_1777(.a(s_178_38), .b(s_178_37), .c(s_178_36), .d(s_178_35), .cin(s_178_34), .o(t_5213), .co(t_5214), .cout(t_5215));
compressor_4_2 u2_1778(.a(s_179_2), .b(s_179_1), .c(s_179_0), .d(t_5188), .cin(t_5191), .o(t_5216), .co(t_5217), .cout(t_5218));
compressor_4_2 u2_1779(.a(s_179_5), .b(s_179_4), .c(s_179_3), .d(t_5194), .cin(t_5197), .o(t_5219), .co(t_5220), .cout(t_5221));
compressor_4_2 u2_1780(.a(s_179_8), .b(s_179_7), .c(s_179_6), .d(t_5200), .cin(t_5203), .o(t_5222), .co(t_5223), .cout(t_5224));
compressor_4_2 u2_1781(.a(s_179_11), .b(s_179_10), .c(s_179_9), .d(t_5206), .cin(t_5209), .o(t_5225), .co(t_5226), .cout(t_5227));
compressor_4_2 u2_1782(.a(s_179_14), .b(s_179_13), .c(s_179_12), .d(t_5212), .cin(t_5215), .o(t_5228), .co(t_5229), .cout(t_5230));
compressor_4_2 u2_1783(.a(s_179_19), .b(s_179_18), .c(s_179_17), .d(s_179_16), .cin(s_179_15), .o(t_5231), .co(t_5232), .cout(t_5233));
compressor_4_2 u2_1784(.a(s_179_24), .b(s_179_23), .c(s_179_22), .d(s_179_21), .cin(s_179_20), .o(t_5234), .co(t_5235), .cout(t_5236));
compressor_4_2 u2_1785(.a(s_179_29), .b(s_179_28), .c(s_179_27), .d(s_179_26), .cin(s_179_25), .o(t_5237), .co(t_5238), .cout(t_5239));
compressor_4_2 u2_1786(.a(s_179_34), .b(s_179_33), .c(s_179_32), .d(s_179_31), .cin(s_179_30), .o(t_5240), .co(t_5241), .cout(t_5242));
compressor_4_2 u2_1787(.a(s_179_39), .b(s_179_38), .c(s_179_37), .d(s_179_36), .cin(s_179_35), .o(t_5243), .co(t_5244), .cout(t_5245));
compressor_4_2 u2_1788(.a(s_180_2), .b(s_180_1), .c(s_180_0), .d(t_5218), .cin(t_5221), .o(t_5246), .co(t_5247), .cout(t_5248));
compressor_4_2 u2_1789(.a(s_180_5), .b(s_180_4), .c(s_180_3), .d(t_5224), .cin(t_5227), .o(t_5249), .co(t_5250), .cout(t_5251));
compressor_4_2 u2_1790(.a(s_180_8), .b(s_180_7), .c(s_180_6), .d(t_5230), .cin(t_5233), .o(t_5252), .co(t_5253), .cout(t_5254));
compressor_4_2 u2_1791(.a(s_180_11), .b(s_180_10), .c(s_180_9), .d(t_5236), .cin(t_5239), .o(t_5255), .co(t_5256), .cout(t_5257));
compressor_4_2 u2_1792(.a(s_180_14), .b(s_180_13), .c(s_180_12), .d(t_5242), .cin(t_5245), .o(t_5258), .co(t_5259), .cout(t_5260));
compressor_4_2 u2_1793(.a(s_180_19), .b(s_180_18), .c(s_180_17), .d(s_180_16), .cin(s_180_15), .o(t_5261), .co(t_5262), .cout(t_5263));
compressor_4_2 u2_1794(.a(s_180_24), .b(s_180_23), .c(s_180_22), .d(s_180_21), .cin(s_180_20), .o(t_5264), .co(t_5265), .cout(t_5266));
compressor_4_2 u2_1795(.a(s_180_29), .b(s_180_28), .c(s_180_27), .d(s_180_26), .cin(s_180_25), .o(t_5267), .co(t_5268), .cout(t_5269));
compressor_4_2 u2_1796(.a(s_180_34), .b(s_180_33), .c(s_180_32), .d(s_180_31), .cin(s_180_30), .o(t_5270), .co(t_5271), .cout(t_5272));
compressor_3_2 u1_1797(.a(s_180_37), .b(s_180_36), .cin(s_180_35), .o(t_5273), .cout(t_5274));
compressor_4_2 u2_1798(.a(s_181_2), .b(s_181_1), .c(s_181_0), .d(t_5248), .cin(t_5251), .o(t_5275), .co(t_5276), .cout(t_5277));
compressor_4_2 u2_1799(.a(s_181_5), .b(s_181_4), .c(s_181_3), .d(t_5254), .cin(t_5257), .o(t_5278), .co(t_5279), .cout(t_5280));
compressor_4_2 u2_1800(.a(s_181_8), .b(s_181_7), .c(s_181_6), .d(t_5260), .cin(t_5263), .o(t_5281), .co(t_5282), .cout(t_5283));
compressor_4_2 u2_1801(.a(s_181_11), .b(s_181_10), .c(s_181_9), .d(t_5266), .cin(t_5269), .o(t_5284), .co(t_5285), .cout(t_5286));
compressor_4_2 u2_1802(.a(s_181_14), .b(s_181_13), .c(s_181_12), .d(t_5272), .cin(t_5274), .o(t_5287), .co(t_5288), .cout(t_5289));
compressor_4_2 u2_1803(.a(s_181_19), .b(s_181_18), .c(s_181_17), .d(s_181_16), .cin(s_181_15), .o(t_5290), .co(t_5291), .cout(t_5292));
compressor_4_2 u2_1804(.a(s_181_24), .b(s_181_23), .c(s_181_22), .d(s_181_21), .cin(s_181_20), .o(t_5293), .co(t_5294), .cout(t_5295));
compressor_4_2 u2_1805(.a(s_181_29), .b(s_181_28), .c(s_181_27), .d(s_181_26), .cin(s_181_25), .o(t_5296), .co(t_5297), .cout(t_5298));
compressor_4_2 u2_1806(.a(s_181_34), .b(s_181_33), .c(s_181_32), .d(s_181_31), .cin(s_181_30), .o(t_5299), .co(t_5300), .cout(t_5301));
compressor_3_2 u1_1807(.a(s_181_37), .b(s_181_36), .cin(s_181_35), .o(t_5302), .cout(t_5303));
compressor_4_2 u2_1808(.a(s_182_2), .b(s_182_1), .c(s_182_0), .d(t_5277), .cin(t_5280), .o(t_5304), .co(t_5305), .cout(t_5306));
compressor_4_2 u2_1809(.a(s_182_5), .b(s_182_4), .c(s_182_3), .d(t_5283), .cin(t_5286), .o(t_5307), .co(t_5308), .cout(t_5309));
compressor_4_2 u2_1810(.a(s_182_8), .b(s_182_7), .c(s_182_6), .d(t_5289), .cin(t_5292), .o(t_5310), .co(t_5311), .cout(t_5312));
compressor_4_2 u2_1811(.a(s_182_11), .b(s_182_10), .c(s_182_9), .d(t_5295), .cin(t_5298), .o(t_5313), .co(t_5314), .cout(t_5315));
compressor_4_2 u2_1812(.a(s_182_14), .b(s_182_13), .c(s_182_12), .d(t_5301), .cin(t_5303), .o(t_5316), .co(t_5317), .cout(t_5318));
compressor_4_2 u2_1813(.a(s_182_19), .b(s_182_18), .c(s_182_17), .d(s_182_16), .cin(s_182_15), .o(t_5319), .co(t_5320), .cout(t_5321));
compressor_4_2 u2_1814(.a(s_182_24), .b(s_182_23), .c(s_182_22), .d(s_182_21), .cin(s_182_20), .o(t_5322), .co(t_5323), .cout(t_5324));
compressor_4_2 u2_1815(.a(s_182_29), .b(s_182_28), .c(s_182_27), .d(s_182_26), .cin(s_182_25), .o(t_5325), .co(t_5326), .cout(t_5327));
compressor_4_2 u2_1816(.a(s_182_34), .b(s_182_33), .c(s_182_32), .d(s_182_31), .cin(s_182_30), .o(t_5328), .co(t_5329), .cout(t_5330));
compressor_3_2 u1_1817(.a(s_182_37), .b(s_182_36), .cin(s_182_35), .o(t_5331), .cout(t_5332));
compressor_4_2 u2_1818(.a(s_183_2), .b(s_183_1), .c(s_183_0), .d(t_5306), .cin(t_5309), .o(t_5333), .co(t_5334), .cout(t_5335));
compressor_4_2 u2_1819(.a(s_183_5), .b(s_183_4), .c(s_183_3), .d(t_5312), .cin(t_5315), .o(t_5336), .co(t_5337), .cout(t_5338));
compressor_4_2 u2_1820(.a(s_183_8), .b(s_183_7), .c(s_183_6), .d(t_5318), .cin(t_5321), .o(t_5339), .co(t_5340), .cout(t_5341));
compressor_4_2 u2_1821(.a(s_183_11), .b(s_183_10), .c(s_183_9), .d(t_5324), .cin(t_5327), .o(t_5342), .co(t_5343), .cout(t_5344));
compressor_4_2 u2_1822(.a(s_183_14), .b(s_183_13), .c(s_183_12), .d(t_5330), .cin(t_5332), .o(t_5345), .co(t_5346), .cout(t_5347));
compressor_4_2 u2_1823(.a(s_183_19), .b(s_183_18), .c(s_183_17), .d(s_183_16), .cin(s_183_15), .o(t_5348), .co(t_5349), .cout(t_5350));
compressor_4_2 u2_1824(.a(s_183_24), .b(s_183_23), .c(s_183_22), .d(s_183_21), .cin(s_183_20), .o(t_5351), .co(t_5352), .cout(t_5353));
compressor_4_2 u2_1825(.a(s_183_29), .b(s_183_28), .c(s_183_27), .d(s_183_26), .cin(s_183_25), .o(t_5354), .co(t_5355), .cout(t_5356));
compressor_4_2 u2_1826(.a(s_183_34), .b(s_183_33), .c(s_183_32), .d(s_183_31), .cin(s_183_30), .o(t_5357), .co(t_5358), .cout(t_5359));
compressor_3_2 u1_1827(.a(s_183_37), .b(s_183_36), .cin(s_183_35), .o(t_5360), .cout(t_5361));
compressor_4_2 u2_1828(.a(s_184_2), .b(s_184_1), .c(s_184_0), .d(t_5335), .cin(t_5338), .o(t_5362), .co(t_5363), .cout(t_5364));
compressor_4_2 u2_1829(.a(s_184_5), .b(s_184_4), .c(s_184_3), .d(t_5341), .cin(t_5344), .o(t_5365), .co(t_5366), .cout(t_5367));
compressor_4_2 u2_1830(.a(s_184_8), .b(s_184_7), .c(s_184_6), .d(t_5347), .cin(t_5350), .o(t_5368), .co(t_5369), .cout(t_5370));
compressor_4_2 u2_1831(.a(s_184_11), .b(s_184_10), .c(s_184_9), .d(t_5353), .cin(t_5356), .o(t_5371), .co(t_5372), .cout(t_5373));
compressor_4_2 u2_1832(.a(s_184_14), .b(s_184_13), .c(s_184_12), .d(t_5359), .cin(t_5361), .o(t_5374), .co(t_5375), .cout(t_5376));
compressor_4_2 u2_1833(.a(s_184_19), .b(s_184_18), .c(s_184_17), .d(s_184_16), .cin(s_184_15), .o(t_5377), .co(t_5378), .cout(t_5379));
compressor_4_2 u2_1834(.a(s_184_24), .b(s_184_23), .c(s_184_22), .d(s_184_21), .cin(s_184_20), .o(t_5380), .co(t_5381), .cout(t_5382));
compressor_4_2 u2_1835(.a(s_184_29), .b(s_184_28), .c(s_184_27), .d(s_184_26), .cin(s_184_25), .o(t_5383), .co(t_5384), .cout(t_5385));
compressor_4_2 u2_1836(.a(s_184_34), .b(s_184_33), .c(s_184_32), .d(s_184_31), .cin(s_184_30), .o(t_5386), .co(t_5387), .cout(t_5388));
half_adder u0_1837(.a(s_184_36), .b(s_184_35), .o(t_5389), .cout(t_5390));
compressor_4_2 u2_1838(.a(s_185_2), .b(s_185_1), .c(s_185_0), .d(t_5364), .cin(t_5367), .o(t_5391), .co(t_5392), .cout(t_5393));
compressor_4_2 u2_1839(.a(s_185_5), .b(s_185_4), .c(s_185_3), .d(t_5370), .cin(t_5373), .o(t_5394), .co(t_5395), .cout(t_5396));
compressor_4_2 u2_1840(.a(s_185_8), .b(s_185_7), .c(s_185_6), .d(t_5376), .cin(t_5379), .o(t_5397), .co(t_5398), .cout(t_5399));
compressor_4_2 u2_1841(.a(s_185_11), .b(s_185_10), .c(s_185_9), .d(t_5382), .cin(t_5385), .o(t_5400), .co(t_5401), .cout(t_5402));
compressor_4_2 u2_1842(.a(s_185_14), .b(s_185_13), .c(s_185_12), .d(t_5388), .cin(t_5390), .o(t_5403), .co(t_5404), .cout(t_5405));
compressor_4_2 u2_1843(.a(s_185_19), .b(s_185_18), .c(s_185_17), .d(s_185_16), .cin(s_185_15), .o(t_5406), .co(t_5407), .cout(t_5408));
compressor_4_2 u2_1844(.a(s_185_24), .b(s_185_23), .c(s_185_22), .d(s_185_21), .cin(s_185_20), .o(t_5409), .co(t_5410), .cout(t_5411));
compressor_4_2 u2_1845(.a(s_185_29), .b(s_185_28), .c(s_185_27), .d(s_185_26), .cin(s_185_25), .o(t_5412), .co(t_5413), .cout(t_5414));
compressor_4_2 u2_1846(.a(s_185_34), .b(s_185_33), .c(s_185_32), .d(s_185_31), .cin(s_185_30), .o(t_5415), .co(t_5416), .cout(t_5417));
half_adder u0_1847(.a(s_185_36), .b(s_185_35), .o(t_5418), .cout(t_5419));
compressor_4_2 u2_1848(.a(s_186_2), .b(s_186_1), .c(s_186_0), .d(t_5393), .cin(t_5396), .o(t_5420), .co(t_5421), .cout(t_5422));
compressor_4_2 u2_1849(.a(s_186_5), .b(s_186_4), .c(s_186_3), .d(t_5399), .cin(t_5402), .o(t_5423), .co(t_5424), .cout(t_5425));
compressor_4_2 u2_1850(.a(s_186_8), .b(s_186_7), .c(s_186_6), .d(t_5405), .cin(t_5408), .o(t_5426), .co(t_5427), .cout(t_5428));
compressor_4_2 u2_1851(.a(s_186_11), .b(s_186_10), .c(s_186_9), .d(t_5411), .cin(t_5414), .o(t_5429), .co(t_5430), .cout(t_5431));
compressor_4_2 u2_1852(.a(s_186_14), .b(s_186_13), .c(s_186_12), .d(t_5417), .cin(t_5419), .o(t_5432), .co(t_5433), .cout(t_5434));
compressor_4_2 u2_1853(.a(s_186_19), .b(s_186_18), .c(s_186_17), .d(s_186_16), .cin(s_186_15), .o(t_5435), .co(t_5436), .cout(t_5437));
compressor_4_2 u2_1854(.a(s_186_24), .b(s_186_23), .c(s_186_22), .d(s_186_21), .cin(s_186_20), .o(t_5438), .co(t_5439), .cout(t_5440));
compressor_4_2 u2_1855(.a(s_186_29), .b(s_186_28), .c(s_186_27), .d(s_186_26), .cin(s_186_25), .o(t_5441), .co(t_5442), .cout(t_5443));
compressor_4_2 u2_1856(.a(s_186_34), .b(s_186_33), .c(s_186_32), .d(s_186_31), .cin(s_186_30), .o(t_5444), .co(t_5445), .cout(t_5446));
compressor_4_2 u2_1857(.a(s_187_2), .b(s_187_1), .c(s_187_0), .d(t_5422), .cin(t_5425), .o(t_5447), .co(t_5448), .cout(t_5449));
compressor_4_2 u2_1858(.a(s_187_5), .b(s_187_4), .c(s_187_3), .d(t_5428), .cin(t_5431), .o(t_5450), .co(t_5451), .cout(t_5452));
compressor_4_2 u2_1859(.a(s_187_8), .b(s_187_7), .c(s_187_6), .d(t_5434), .cin(t_5437), .o(t_5453), .co(t_5454), .cout(t_5455));
compressor_4_2 u2_1860(.a(s_187_11), .b(s_187_10), .c(s_187_9), .d(t_5440), .cin(t_5443), .o(t_5456), .co(t_5457), .cout(t_5458));
compressor_4_2 u2_1861(.a(s_187_15), .b(s_187_14), .c(s_187_13), .d(s_187_12), .cin(t_5446), .o(t_5459), .co(t_5460), .cout(t_5461));
compressor_4_2 u2_1862(.a(s_187_20), .b(s_187_19), .c(s_187_18), .d(s_187_17), .cin(s_187_16), .o(t_5462), .co(t_5463), .cout(t_5464));
compressor_4_2 u2_1863(.a(s_187_25), .b(s_187_24), .c(s_187_23), .d(s_187_22), .cin(s_187_21), .o(t_5465), .co(t_5466), .cout(t_5467));
compressor_4_2 u2_1864(.a(s_187_30), .b(s_187_29), .c(s_187_28), .d(s_187_27), .cin(s_187_26), .o(t_5468), .co(t_5469), .cout(t_5470));
compressor_4_2 u2_1865(.a(s_187_35), .b(s_187_34), .c(s_187_33), .d(s_187_32), .cin(s_187_31), .o(t_5471), .co(t_5472), .cout(t_5473));
compressor_4_2 u2_1866(.a(s_188_2), .b(s_188_1), .c(s_188_0), .d(t_5449), .cin(t_5452), .o(t_5474), .co(t_5475), .cout(t_5476));
compressor_4_2 u2_1867(.a(s_188_5), .b(s_188_4), .c(s_188_3), .d(t_5455), .cin(t_5458), .o(t_5477), .co(t_5478), .cout(t_5479));
compressor_4_2 u2_1868(.a(s_188_8), .b(s_188_7), .c(s_188_6), .d(t_5461), .cin(t_5464), .o(t_5480), .co(t_5481), .cout(t_5482));
compressor_4_2 u2_1869(.a(s_188_11), .b(s_188_10), .c(s_188_9), .d(t_5467), .cin(t_5470), .o(t_5483), .co(t_5484), .cout(t_5485));
compressor_4_2 u2_1870(.a(s_188_15), .b(s_188_14), .c(s_188_13), .d(s_188_12), .cin(t_5473), .o(t_5486), .co(t_5487), .cout(t_5488));
compressor_4_2 u2_1871(.a(s_188_20), .b(s_188_19), .c(s_188_18), .d(s_188_17), .cin(s_188_16), .o(t_5489), .co(t_5490), .cout(t_5491));
compressor_4_2 u2_1872(.a(s_188_25), .b(s_188_24), .c(s_188_23), .d(s_188_22), .cin(s_188_21), .o(t_5492), .co(t_5493), .cout(t_5494));
compressor_4_2 u2_1873(.a(s_188_30), .b(s_188_29), .c(s_188_28), .d(s_188_27), .cin(s_188_26), .o(t_5495), .co(t_5496), .cout(t_5497));
compressor_3_2 u1_1874(.a(s_188_33), .b(s_188_32), .cin(s_188_31), .o(t_5498), .cout(t_5499));
compressor_4_2 u2_1875(.a(s_189_2), .b(s_189_1), .c(s_189_0), .d(t_5476), .cin(t_5479), .o(t_5500), .co(t_5501), .cout(t_5502));
compressor_4_2 u2_1876(.a(s_189_5), .b(s_189_4), .c(s_189_3), .d(t_5482), .cin(t_5485), .o(t_5503), .co(t_5504), .cout(t_5505));
compressor_4_2 u2_1877(.a(s_189_8), .b(s_189_7), .c(s_189_6), .d(t_5488), .cin(t_5491), .o(t_5506), .co(t_5507), .cout(t_5508));
compressor_4_2 u2_1878(.a(s_189_11), .b(s_189_10), .c(s_189_9), .d(t_5494), .cin(t_5497), .o(t_5509), .co(t_5510), .cout(t_5511));
compressor_4_2 u2_1879(.a(s_189_15), .b(s_189_14), .c(s_189_13), .d(s_189_12), .cin(t_5499), .o(t_5512), .co(t_5513), .cout(t_5514));
compressor_4_2 u2_1880(.a(s_189_20), .b(s_189_19), .c(s_189_18), .d(s_189_17), .cin(s_189_16), .o(t_5515), .co(t_5516), .cout(t_5517));
compressor_4_2 u2_1881(.a(s_189_25), .b(s_189_24), .c(s_189_23), .d(s_189_22), .cin(s_189_21), .o(t_5518), .co(t_5519), .cout(t_5520));
compressor_4_2 u2_1882(.a(s_189_30), .b(s_189_29), .c(s_189_28), .d(s_189_27), .cin(s_189_26), .o(t_5521), .co(t_5522), .cout(t_5523));
compressor_3_2 u1_1883(.a(s_189_33), .b(s_189_32), .cin(s_189_31), .o(t_5524), .cout(t_5525));
compressor_4_2 u2_1884(.a(s_190_2), .b(s_190_1), .c(s_190_0), .d(t_5502), .cin(t_5505), .o(t_5526), .co(t_5527), .cout(t_5528));
compressor_4_2 u2_1885(.a(s_190_5), .b(s_190_4), .c(s_190_3), .d(t_5508), .cin(t_5511), .o(t_5529), .co(t_5530), .cout(t_5531));
compressor_4_2 u2_1886(.a(s_190_8), .b(s_190_7), .c(s_190_6), .d(t_5514), .cin(t_5517), .o(t_5532), .co(t_5533), .cout(t_5534));
compressor_4_2 u2_1887(.a(s_190_11), .b(s_190_10), .c(s_190_9), .d(t_5520), .cin(t_5523), .o(t_5535), .co(t_5536), .cout(t_5537));
compressor_4_2 u2_1888(.a(s_190_15), .b(s_190_14), .c(s_190_13), .d(s_190_12), .cin(t_5525), .o(t_5538), .co(t_5539), .cout(t_5540));
compressor_4_2 u2_1889(.a(s_190_20), .b(s_190_19), .c(s_190_18), .d(s_190_17), .cin(s_190_16), .o(t_5541), .co(t_5542), .cout(t_5543));
compressor_4_2 u2_1890(.a(s_190_25), .b(s_190_24), .c(s_190_23), .d(s_190_22), .cin(s_190_21), .o(t_5544), .co(t_5545), .cout(t_5546));
compressor_4_2 u2_1891(.a(s_190_30), .b(s_190_29), .c(s_190_28), .d(s_190_27), .cin(s_190_26), .o(t_5547), .co(t_5548), .cout(t_5549));
compressor_3_2 u1_1892(.a(s_190_33), .b(s_190_32), .cin(s_190_31), .o(t_5550), .cout(t_5551));
compressor_4_2 u2_1893(.a(s_191_2), .b(s_191_1), .c(s_191_0), .d(t_5528), .cin(t_5531), .o(t_5552), .co(t_5553), .cout(t_5554));
compressor_4_2 u2_1894(.a(s_191_5), .b(s_191_4), .c(s_191_3), .d(t_5534), .cin(t_5537), .o(t_5555), .co(t_5556), .cout(t_5557));
compressor_4_2 u2_1895(.a(s_191_8), .b(s_191_7), .c(s_191_6), .d(t_5540), .cin(t_5543), .o(t_5558), .co(t_5559), .cout(t_5560));
compressor_4_2 u2_1896(.a(s_191_11), .b(s_191_10), .c(s_191_9), .d(t_5546), .cin(t_5549), .o(t_5561), .co(t_5562), .cout(t_5563));
compressor_4_2 u2_1897(.a(s_191_15), .b(s_191_14), .c(s_191_13), .d(s_191_12), .cin(t_5551), .o(t_5564), .co(t_5565), .cout(t_5566));
compressor_4_2 u2_1898(.a(s_191_20), .b(s_191_19), .c(s_191_18), .d(s_191_17), .cin(s_191_16), .o(t_5567), .co(t_5568), .cout(t_5569));
compressor_4_2 u2_1899(.a(s_191_25), .b(s_191_24), .c(s_191_23), .d(s_191_22), .cin(s_191_21), .o(t_5570), .co(t_5571), .cout(t_5572));
compressor_4_2 u2_1900(.a(s_191_30), .b(s_191_29), .c(s_191_28), .d(s_191_27), .cin(s_191_26), .o(t_5573), .co(t_5574), .cout(t_5575));
compressor_3_2 u1_1901(.a(s_191_33), .b(s_191_32), .cin(s_191_31), .o(t_5576), .cout(t_5577));
compressor_4_2 u2_1902(.a(s_192_2), .b(s_192_1), .c(s_192_0), .d(t_5554), .cin(t_5557), .o(t_5578), .co(t_5579), .cout(t_5580));
compressor_4_2 u2_1903(.a(s_192_5), .b(s_192_4), .c(s_192_3), .d(t_5560), .cin(t_5563), .o(t_5581), .co(t_5582), .cout(t_5583));
compressor_4_2 u2_1904(.a(s_192_8), .b(s_192_7), .c(s_192_6), .d(t_5566), .cin(t_5569), .o(t_5584), .co(t_5585), .cout(t_5586));
compressor_4_2 u2_1905(.a(s_192_11), .b(s_192_10), .c(s_192_9), .d(t_5572), .cin(t_5575), .o(t_5587), .co(t_5588), .cout(t_5589));
compressor_4_2 u2_1906(.a(s_192_15), .b(s_192_14), .c(s_192_13), .d(s_192_12), .cin(t_5577), .o(t_5590), .co(t_5591), .cout(t_5592));
compressor_4_2 u2_1907(.a(s_192_20), .b(s_192_19), .c(s_192_18), .d(s_192_17), .cin(s_192_16), .o(t_5593), .co(t_5594), .cout(t_5595));
compressor_4_2 u2_1908(.a(s_192_25), .b(s_192_24), .c(s_192_23), .d(s_192_22), .cin(s_192_21), .o(t_5596), .co(t_5597), .cout(t_5598));
compressor_4_2 u2_1909(.a(s_192_30), .b(s_192_29), .c(s_192_28), .d(s_192_27), .cin(s_192_26), .o(t_5599), .co(t_5600), .cout(t_5601));
half_adder u0_1910(.a(s_192_32), .b(s_192_31), .o(t_5602), .cout(t_5603));
compressor_4_2 u2_1911(.a(s_193_2), .b(s_193_1), .c(s_193_0), .d(t_5580), .cin(t_5583), .o(t_5604), .co(t_5605), .cout(t_5606));
compressor_4_2 u2_1912(.a(s_193_5), .b(s_193_4), .c(s_193_3), .d(t_5586), .cin(t_5589), .o(t_5607), .co(t_5608), .cout(t_5609));
compressor_4_2 u2_1913(.a(s_193_8), .b(s_193_7), .c(s_193_6), .d(t_5592), .cin(t_5595), .o(t_5610), .co(t_5611), .cout(t_5612));
compressor_4_2 u2_1914(.a(s_193_11), .b(s_193_10), .c(s_193_9), .d(t_5598), .cin(t_5601), .o(t_5613), .co(t_5614), .cout(t_5615));
compressor_4_2 u2_1915(.a(s_193_15), .b(s_193_14), .c(s_193_13), .d(s_193_12), .cin(t_5603), .o(t_5616), .co(t_5617), .cout(t_5618));
compressor_4_2 u2_1916(.a(s_193_20), .b(s_193_19), .c(s_193_18), .d(s_193_17), .cin(s_193_16), .o(t_5619), .co(t_5620), .cout(t_5621));
compressor_4_2 u2_1917(.a(s_193_25), .b(s_193_24), .c(s_193_23), .d(s_193_22), .cin(s_193_21), .o(t_5622), .co(t_5623), .cout(t_5624));
compressor_4_2 u2_1918(.a(s_193_30), .b(s_193_29), .c(s_193_28), .d(s_193_27), .cin(s_193_26), .o(t_5625), .co(t_5626), .cout(t_5627));
half_adder u0_1919(.a(s_193_32), .b(s_193_31), .o(t_5628), .cout(t_5629));
compressor_4_2 u2_1920(.a(s_194_2), .b(s_194_1), .c(s_194_0), .d(t_5606), .cin(t_5609), .o(t_5630), .co(t_5631), .cout(t_5632));
compressor_4_2 u2_1921(.a(s_194_5), .b(s_194_4), .c(s_194_3), .d(t_5612), .cin(t_5615), .o(t_5633), .co(t_5634), .cout(t_5635));
compressor_4_2 u2_1922(.a(s_194_8), .b(s_194_7), .c(s_194_6), .d(t_5618), .cin(t_5621), .o(t_5636), .co(t_5637), .cout(t_5638));
compressor_4_2 u2_1923(.a(s_194_11), .b(s_194_10), .c(s_194_9), .d(t_5624), .cin(t_5627), .o(t_5639), .co(t_5640), .cout(t_5641));
compressor_4_2 u2_1924(.a(s_194_15), .b(s_194_14), .c(s_194_13), .d(s_194_12), .cin(t_5629), .o(t_5642), .co(t_5643), .cout(t_5644));
compressor_4_2 u2_1925(.a(s_194_20), .b(s_194_19), .c(s_194_18), .d(s_194_17), .cin(s_194_16), .o(t_5645), .co(t_5646), .cout(t_5647));
compressor_4_2 u2_1926(.a(s_194_25), .b(s_194_24), .c(s_194_23), .d(s_194_22), .cin(s_194_21), .o(t_5648), .co(t_5649), .cout(t_5650));
compressor_4_2 u2_1927(.a(s_194_30), .b(s_194_29), .c(s_194_28), .d(s_194_27), .cin(s_194_26), .o(t_5651), .co(t_5652), .cout(t_5653));
compressor_4_2 u2_1928(.a(s_195_2), .b(s_195_1), .c(s_195_0), .d(t_5632), .cin(t_5635), .o(t_5654), .co(t_5655), .cout(t_5656));
compressor_4_2 u2_1929(.a(s_195_5), .b(s_195_4), .c(s_195_3), .d(t_5638), .cin(t_5641), .o(t_5657), .co(t_5658), .cout(t_5659));
compressor_4_2 u2_1930(.a(s_195_8), .b(s_195_7), .c(s_195_6), .d(t_5644), .cin(t_5647), .o(t_5660), .co(t_5661), .cout(t_5662));
compressor_4_2 u2_1931(.a(s_195_11), .b(s_195_10), .c(s_195_9), .d(t_5650), .cin(t_5653), .o(t_5663), .co(t_5664), .cout(t_5665));
compressor_4_2 u2_1932(.a(s_195_16), .b(s_195_15), .c(s_195_14), .d(s_195_13), .cin(s_195_12), .o(t_5666), .co(t_5667), .cout(t_5668));
compressor_4_2 u2_1933(.a(s_195_21), .b(s_195_20), .c(s_195_19), .d(s_195_18), .cin(s_195_17), .o(t_5669), .co(t_5670), .cout(t_5671));
compressor_4_2 u2_1934(.a(s_195_26), .b(s_195_25), .c(s_195_24), .d(s_195_23), .cin(s_195_22), .o(t_5672), .co(t_5673), .cout(t_5674));
compressor_4_2 u2_1935(.a(s_195_31), .b(s_195_30), .c(s_195_29), .d(s_195_28), .cin(s_195_27), .o(t_5675), .co(t_5676), .cout(t_5677));
compressor_4_2 u2_1936(.a(s_196_2), .b(s_196_1), .c(s_196_0), .d(t_5656), .cin(t_5659), .o(t_5678), .co(t_5679), .cout(t_5680));
compressor_4_2 u2_1937(.a(s_196_5), .b(s_196_4), .c(s_196_3), .d(t_5662), .cin(t_5665), .o(t_5681), .co(t_5682), .cout(t_5683));
compressor_4_2 u2_1938(.a(s_196_8), .b(s_196_7), .c(s_196_6), .d(t_5668), .cin(t_5671), .o(t_5684), .co(t_5685), .cout(t_5686));
compressor_4_2 u2_1939(.a(s_196_11), .b(s_196_10), .c(s_196_9), .d(t_5674), .cin(t_5677), .o(t_5687), .co(t_5688), .cout(t_5689));
compressor_4_2 u2_1940(.a(s_196_16), .b(s_196_15), .c(s_196_14), .d(s_196_13), .cin(s_196_12), .o(t_5690), .co(t_5691), .cout(t_5692));
compressor_4_2 u2_1941(.a(s_196_21), .b(s_196_20), .c(s_196_19), .d(s_196_18), .cin(s_196_17), .o(t_5693), .co(t_5694), .cout(t_5695));
compressor_4_2 u2_1942(.a(s_196_26), .b(s_196_25), .c(s_196_24), .d(s_196_23), .cin(s_196_22), .o(t_5696), .co(t_5697), .cout(t_5698));
compressor_3_2 u1_1943(.a(s_196_29), .b(s_196_28), .cin(s_196_27), .o(t_5699), .cout(t_5700));
compressor_4_2 u2_1944(.a(s_197_2), .b(s_197_1), .c(s_197_0), .d(t_5680), .cin(t_5683), .o(t_5701), .co(t_5702), .cout(t_5703));
compressor_4_2 u2_1945(.a(s_197_5), .b(s_197_4), .c(s_197_3), .d(t_5686), .cin(t_5689), .o(t_5704), .co(t_5705), .cout(t_5706));
compressor_4_2 u2_1946(.a(s_197_8), .b(s_197_7), .c(s_197_6), .d(t_5692), .cin(t_5695), .o(t_5707), .co(t_5708), .cout(t_5709));
compressor_4_2 u2_1947(.a(s_197_11), .b(s_197_10), .c(s_197_9), .d(t_5698), .cin(t_5700), .o(t_5710), .co(t_5711), .cout(t_5712));
compressor_4_2 u2_1948(.a(s_197_16), .b(s_197_15), .c(s_197_14), .d(s_197_13), .cin(s_197_12), .o(t_5713), .co(t_5714), .cout(t_5715));
compressor_4_2 u2_1949(.a(s_197_21), .b(s_197_20), .c(s_197_19), .d(s_197_18), .cin(s_197_17), .o(t_5716), .co(t_5717), .cout(t_5718));
compressor_4_2 u2_1950(.a(s_197_26), .b(s_197_25), .c(s_197_24), .d(s_197_23), .cin(s_197_22), .o(t_5719), .co(t_5720), .cout(t_5721));
compressor_3_2 u1_1951(.a(s_197_29), .b(s_197_28), .cin(s_197_27), .o(t_5722), .cout(t_5723));
compressor_4_2 u2_1952(.a(s_198_2), .b(s_198_1), .c(s_198_0), .d(t_5703), .cin(t_5706), .o(t_5724), .co(t_5725), .cout(t_5726));
compressor_4_2 u2_1953(.a(s_198_5), .b(s_198_4), .c(s_198_3), .d(t_5709), .cin(t_5712), .o(t_5727), .co(t_5728), .cout(t_5729));
compressor_4_2 u2_1954(.a(s_198_8), .b(s_198_7), .c(s_198_6), .d(t_5715), .cin(t_5718), .o(t_5730), .co(t_5731), .cout(t_5732));
compressor_4_2 u2_1955(.a(s_198_11), .b(s_198_10), .c(s_198_9), .d(t_5721), .cin(t_5723), .o(t_5733), .co(t_5734), .cout(t_5735));
compressor_4_2 u2_1956(.a(s_198_16), .b(s_198_15), .c(s_198_14), .d(s_198_13), .cin(s_198_12), .o(t_5736), .co(t_5737), .cout(t_5738));
compressor_4_2 u2_1957(.a(s_198_21), .b(s_198_20), .c(s_198_19), .d(s_198_18), .cin(s_198_17), .o(t_5739), .co(t_5740), .cout(t_5741));
compressor_4_2 u2_1958(.a(s_198_26), .b(s_198_25), .c(s_198_24), .d(s_198_23), .cin(s_198_22), .o(t_5742), .co(t_5743), .cout(t_5744));
compressor_3_2 u1_1959(.a(s_198_29), .b(s_198_28), .cin(s_198_27), .o(t_5745), .cout(t_5746));
compressor_4_2 u2_1960(.a(s_199_2), .b(s_199_1), .c(s_199_0), .d(t_5726), .cin(t_5729), .o(t_5747), .co(t_5748), .cout(t_5749));
compressor_4_2 u2_1961(.a(s_199_5), .b(s_199_4), .c(s_199_3), .d(t_5732), .cin(t_5735), .o(t_5750), .co(t_5751), .cout(t_5752));
compressor_4_2 u2_1962(.a(s_199_8), .b(s_199_7), .c(s_199_6), .d(t_5738), .cin(t_5741), .o(t_5753), .co(t_5754), .cout(t_5755));
compressor_4_2 u2_1963(.a(s_199_11), .b(s_199_10), .c(s_199_9), .d(t_5744), .cin(t_5746), .o(t_5756), .co(t_5757), .cout(t_5758));
compressor_4_2 u2_1964(.a(s_199_16), .b(s_199_15), .c(s_199_14), .d(s_199_13), .cin(s_199_12), .o(t_5759), .co(t_5760), .cout(t_5761));
compressor_4_2 u2_1965(.a(s_199_21), .b(s_199_20), .c(s_199_19), .d(s_199_18), .cin(s_199_17), .o(t_5762), .co(t_5763), .cout(t_5764));
compressor_4_2 u2_1966(.a(s_199_26), .b(s_199_25), .c(s_199_24), .d(s_199_23), .cin(s_199_22), .o(t_5765), .co(t_5766), .cout(t_5767));
compressor_3_2 u1_1967(.a(s_199_29), .b(s_199_28), .cin(s_199_27), .o(t_5768), .cout(t_5769));
compressor_4_2 u2_1968(.a(s_200_2), .b(s_200_1), .c(s_200_0), .d(t_5749), .cin(t_5752), .o(t_5770), .co(t_5771), .cout(t_5772));
compressor_4_2 u2_1969(.a(s_200_5), .b(s_200_4), .c(s_200_3), .d(t_5755), .cin(t_5758), .o(t_5773), .co(t_5774), .cout(t_5775));
compressor_4_2 u2_1970(.a(s_200_8), .b(s_200_7), .c(s_200_6), .d(t_5761), .cin(t_5764), .o(t_5776), .co(t_5777), .cout(t_5778));
compressor_4_2 u2_1971(.a(s_200_11), .b(s_200_10), .c(s_200_9), .d(t_5767), .cin(t_5769), .o(t_5779), .co(t_5780), .cout(t_5781));
compressor_4_2 u2_1972(.a(s_200_16), .b(s_200_15), .c(s_200_14), .d(s_200_13), .cin(s_200_12), .o(t_5782), .co(t_5783), .cout(t_5784));
compressor_4_2 u2_1973(.a(s_200_21), .b(s_200_20), .c(s_200_19), .d(s_200_18), .cin(s_200_17), .o(t_5785), .co(t_5786), .cout(t_5787));
compressor_4_2 u2_1974(.a(s_200_26), .b(s_200_25), .c(s_200_24), .d(s_200_23), .cin(s_200_22), .o(t_5788), .co(t_5789), .cout(t_5790));
half_adder u0_1975(.a(s_200_28), .b(s_200_27), .o(t_5791), .cout(t_5792));
compressor_4_2 u2_1976(.a(s_201_2), .b(s_201_1), .c(s_201_0), .d(t_5772), .cin(t_5775), .o(t_5793), .co(t_5794), .cout(t_5795));
compressor_4_2 u2_1977(.a(s_201_5), .b(s_201_4), .c(s_201_3), .d(t_5778), .cin(t_5781), .o(t_5796), .co(t_5797), .cout(t_5798));
compressor_4_2 u2_1978(.a(s_201_8), .b(s_201_7), .c(s_201_6), .d(t_5784), .cin(t_5787), .o(t_5799), .co(t_5800), .cout(t_5801));
compressor_4_2 u2_1979(.a(s_201_11), .b(s_201_10), .c(s_201_9), .d(t_5790), .cin(t_5792), .o(t_5802), .co(t_5803), .cout(t_5804));
compressor_4_2 u2_1980(.a(s_201_16), .b(s_201_15), .c(s_201_14), .d(s_201_13), .cin(s_201_12), .o(t_5805), .co(t_5806), .cout(t_5807));
compressor_4_2 u2_1981(.a(s_201_21), .b(s_201_20), .c(s_201_19), .d(s_201_18), .cin(s_201_17), .o(t_5808), .co(t_5809), .cout(t_5810));
compressor_4_2 u2_1982(.a(s_201_26), .b(s_201_25), .c(s_201_24), .d(s_201_23), .cin(s_201_22), .o(t_5811), .co(t_5812), .cout(t_5813));
half_adder u0_1983(.a(s_201_28), .b(s_201_27), .o(t_5814), .cout(t_5815));
compressor_4_2 u2_1984(.a(s_202_2), .b(s_202_1), .c(s_202_0), .d(t_5795), .cin(t_5798), .o(t_5816), .co(t_5817), .cout(t_5818));
compressor_4_2 u2_1985(.a(s_202_5), .b(s_202_4), .c(s_202_3), .d(t_5801), .cin(t_5804), .o(t_5819), .co(t_5820), .cout(t_5821));
compressor_4_2 u2_1986(.a(s_202_8), .b(s_202_7), .c(s_202_6), .d(t_5807), .cin(t_5810), .o(t_5822), .co(t_5823), .cout(t_5824));
compressor_4_2 u2_1987(.a(s_202_11), .b(s_202_10), .c(s_202_9), .d(t_5813), .cin(t_5815), .o(t_5825), .co(t_5826), .cout(t_5827));
compressor_4_2 u2_1988(.a(s_202_16), .b(s_202_15), .c(s_202_14), .d(s_202_13), .cin(s_202_12), .o(t_5828), .co(t_5829), .cout(t_5830));
compressor_4_2 u2_1989(.a(s_202_21), .b(s_202_20), .c(s_202_19), .d(s_202_18), .cin(s_202_17), .o(t_5831), .co(t_5832), .cout(t_5833));
compressor_4_2 u2_1990(.a(s_202_26), .b(s_202_25), .c(s_202_24), .d(s_202_23), .cin(s_202_22), .o(t_5834), .co(t_5835), .cout(t_5836));
compressor_4_2 u2_1991(.a(s_203_2), .b(s_203_1), .c(s_203_0), .d(t_5818), .cin(t_5821), .o(t_5837), .co(t_5838), .cout(t_5839));
compressor_4_2 u2_1992(.a(s_203_5), .b(s_203_4), .c(s_203_3), .d(t_5824), .cin(t_5827), .o(t_5840), .co(t_5841), .cout(t_5842));
compressor_4_2 u2_1993(.a(s_203_8), .b(s_203_7), .c(s_203_6), .d(t_5830), .cin(t_5833), .o(t_5843), .co(t_5844), .cout(t_5845));
compressor_4_2 u2_1994(.a(s_203_12), .b(s_203_11), .c(s_203_10), .d(s_203_9), .cin(t_5836), .o(t_5846), .co(t_5847), .cout(t_5848));
compressor_4_2 u2_1995(.a(s_203_17), .b(s_203_16), .c(s_203_15), .d(s_203_14), .cin(s_203_13), .o(t_5849), .co(t_5850), .cout(t_5851));
compressor_4_2 u2_1996(.a(s_203_22), .b(s_203_21), .c(s_203_20), .d(s_203_19), .cin(s_203_18), .o(t_5852), .co(t_5853), .cout(t_5854));
compressor_4_2 u2_1997(.a(s_203_27), .b(s_203_26), .c(s_203_25), .d(s_203_24), .cin(s_203_23), .o(t_5855), .co(t_5856), .cout(t_5857));
compressor_4_2 u2_1998(.a(s_204_2), .b(s_204_1), .c(s_204_0), .d(t_5839), .cin(t_5842), .o(t_5858), .co(t_5859), .cout(t_5860));
compressor_4_2 u2_1999(.a(s_204_5), .b(s_204_4), .c(s_204_3), .d(t_5845), .cin(t_5848), .o(t_5861), .co(t_5862), .cout(t_5863));
compressor_4_2 u2_2000(.a(s_204_8), .b(s_204_7), .c(s_204_6), .d(t_5851), .cin(t_5854), .o(t_5864), .co(t_5865), .cout(t_5866));
compressor_4_2 u2_2001(.a(s_204_12), .b(s_204_11), .c(s_204_10), .d(s_204_9), .cin(t_5857), .o(t_5867), .co(t_5868), .cout(t_5869));
compressor_4_2 u2_2002(.a(s_204_17), .b(s_204_16), .c(s_204_15), .d(s_204_14), .cin(s_204_13), .o(t_5870), .co(t_5871), .cout(t_5872));
compressor_4_2 u2_2003(.a(s_204_22), .b(s_204_21), .c(s_204_20), .d(s_204_19), .cin(s_204_18), .o(t_5873), .co(t_5874), .cout(t_5875));
compressor_3_2 u1_2004(.a(s_204_25), .b(s_204_24), .cin(s_204_23), .o(t_5876), .cout(t_5877));
compressor_4_2 u2_2005(.a(s_205_2), .b(s_205_1), .c(s_205_0), .d(t_5860), .cin(t_5863), .o(t_5878), .co(t_5879), .cout(t_5880));
compressor_4_2 u2_2006(.a(s_205_5), .b(s_205_4), .c(s_205_3), .d(t_5866), .cin(t_5869), .o(t_5881), .co(t_5882), .cout(t_5883));
compressor_4_2 u2_2007(.a(s_205_8), .b(s_205_7), .c(s_205_6), .d(t_5872), .cin(t_5875), .o(t_5884), .co(t_5885), .cout(t_5886));
compressor_4_2 u2_2008(.a(s_205_12), .b(s_205_11), .c(s_205_10), .d(s_205_9), .cin(t_5877), .o(t_5887), .co(t_5888), .cout(t_5889));
compressor_4_2 u2_2009(.a(s_205_17), .b(s_205_16), .c(s_205_15), .d(s_205_14), .cin(s_205_13), .o(t_5890), .co(t_5891), .cout(t_5892));
compressor_4_2 u2_2010(.a(s_205_22), .b(s_205_21), .c(s_205_20), .d(s_205_19), .cin(s_205_18), .o(t_5893), .co(t_5894), .cout(t_5895));
compressor_3_2 u1_2011(.a(s_205_25), .b(s_205_24), .cin(s_205_23), .o(t_5896), .cout(t_5897));
compressor_4_2 u2_2012(.a(s_206_2), .b(s_206_1), .c(s_206_0), .d(t_5880), .cin(t_5883), .o(t_5898), .co(t_5899), .cout(t_5900));
compressor_4_2 u2_2013(.a(s_206_5), .b(s_206_4), .c(s_206_3), .d(t_5886), .cin(t_5889), .o(t_5901), .co(t_5902), .cout(t_5903));
compressor_4_2 u2_2014(.a(s_206_8), .b(s_206_7), .c(s_206_6), .d(t_5892), .cin(t_5895), .o(t_5904), .co(t_5905), .cout(t_5906));
compressor_4_2 u2_2015(.a(s_206_12), .b(s_206_11), .c(s_206_10), .d(s_206_9), .cin(t_5897), .o(t_5907), .co(t_5908), .cout(t_5909));
compressor_4_2 u2_2016(.a(s_206_17), .b(s_206_16), .c(s_206_15), .d(s_206_14), .cin(s_206_13), .o(t_5910), .co(t_5911), .cout(t_5912));
compressor_4_2 u2_2017(.a(s_206_22), .b(s_206_21), .c(s_206_20), .d(s_206_19), .cin(s_206_18), .o(t_5913), .co(t_5914), .cout(t_5915));
compressor_3_2 u1_2018(.a(s_206_25), .b(s_206_24), .cin(s_206_23), .o(t_5916), .cout(t_5917));
compressor_4_2 u2_2019(.a(s_207_2), .b(s_207_1), .c(s_207_0), .d(t_5900), .cin(t_5903), .o(t_5918), .co(t_5919), .cout(t_5920));
compressor_4_2 u2_2020(.a(s_207_5), .b(s_207_4), .c(s_207_3), .d(t_5906), .cin(t_5909), .o(t_5921), .co(t_5922), .cout(t_5923));
compressor_4_2 u2_2021(.a(s_207_8), .b(s_207_7), .c(s_207_6), .d(t_5912), .cin(t_5915), .o(t_5924), .co(t_5925), .cout(t_5926));
compressor_4_2 u2_2022(.a(s_207_12), .b(s_207_11), .c(s_207_10), .d(s_207_9), .cin(t_5917), .o(t_5927), .co(t_5928), .cout(t_5929));
compressor_4_2 u2_2023(.a(s_207_17), .b(s_207_16), .c(s_207_15), .d(s_207_14), .cin(s_207_13), .o(t_5930), .co(t_5931), .cout(t_5932));
compressor_4_2 u2_2024(.a(s_207_22), .b(s_207_21), .c(s_207_20), .d(s_207_19), .cin(s_207_18), .o(t_5933), .co(t_5934), .cout(t_5935));
compressor_3_2 u1_2025(.a(s_207_25), .b(s_207_24), .cin(s_207_23), .o(t_5936), .cout(t_5937));
compressor_4_2 u2_2026(.a(s_208_2), .b(s_208_1), .c(s_208_0), .d(t_5920), .cin(t_5923), .o(t_5938), .co(t_5939), .cout(t_5940));
compressor_4_2 u2_2027(.a(s_208_5), .b(s_208_4), .c(s_208_3), .d(t_5926), .cin(t_5929), .o(t_5941), .co(t_5942), .cout(t_5943));
compressor_4_2 u2_2028(.a(s_208_8), .b(s_208_7), .c(s_208_6), .d(t_5932), .cin(t_5935), .o(t_5944), .co(t_5945), .cout(t_5946));
compressor_4_2 u2_2029(.a(s_208_12), .b(s_208_11), .c(s_208_10), .d(s_208_9), .cin(t_5937), .o(t_5947), .co(t_5948), .cout(t_5949));
compressor_4_2 u2_2030(.a(s_208_17), .b(s_208_16), .c(s_208_15), .d(s_208_14), .cin(s_208_13), .o(t_5950), .co(t_5951), .cout(t_5952));
compressor_4_2 u2_2031(.a(s_208_22), .b(s_208_21), .c(s_208_20), .d(s_208_19), .cin(s_208_18), .o(t_5953), .co(t_5954), .cout(t_5955));
half_adder u0_2032(.a(s_208_24), .b(s_208_23), .o(t_5956), .cout(t_5957));
compressor_4_2 u2_2033(.a(s_209_2), .b(s_209_1), .c(s_209_0), .d(t_5940), .cin(t_5943), .o(t_5958), .co(t_5959), .cout(t_5960));
compressor_4_2 u2_2034(.a(s_209_5), .b(s_209_4), .c(s_209_3), .d(t_5946), .cin(t_5949), .o(t_5961), .co(t_5962), .cout(t_5963));
compressor_4_2 u2_2035(.a(s_209_8), .b(s_209_7), .c(s_209_6), .d(t_5952), .cin(t_5955), .o(t_5964), .co(t_5965), .cout(t_5966));
compressor_4_2 u2_2036(.a(s_209_12), .b(s_209_11), .c(s_209_10), .d(s_209_9), .cin(t_5957), .o(t_5967), .co(t_5968), .cout(t_5969));
compressor_4_2 u2_2037(.a(s_209_17), .b(s_209_16), .c(s_209_15), .d(s_209_14), .cin(s_209_13), .o(t_5970), .co(t_5971), .cout(t_5972));
compressor_4_2 u2_2038(.a(s_209_22), .b(s_209_21), .c(s_209_20), .d(s_209_19), .cin(s_209_18), .o(t_5973), .co(t_5974), .cout(t_5975));
half_adder u0_2039(.a(s_209_24), .b(s_209_23), .o(t_5976), .cout(t_5977));
compressor_4_2 u2_2040(.a(s_210_2), .b(s_210_1), .c(s_210_0), .d(t_5960), .cin(t_5963), .o(t_5978), .co(t_5979), .cout(t_5980));
compressor_4_2 u2_2041(.a(s_210_5), .b(s_210_4), .c(s_210_3), .d(t_5966), .cin(t_5969), .o(t_5981), .co(t_5982), .cout(t_5983));
compressor_4_2 u2_2042(.a(s_210_8), .b(s_210_7), .c(s_210_6), .d(t_5972), .cin(t_5975), .o(t_5984), .co(t_5985), .cout(t_5986));
compressor_4_2 u2_2043(.a(s_210_12), .b(s_210_11), .c(s_210_10), .d(s_210_9), .cin(t_5977), .o(t_5987), .co(t_5988), .cout(t_5989));
compressor_4_2 u2_2044(.a(s_210_17), .b(s_210_16), .c(s_210_15), .d(s_210_14), .cin(s_210_13), .o(t_5990), .co(t_5991), .cout(t_5992));
compressor_4_2 u2_2045(.a(s_210_22), .b(s_210_21), .c(s_210_20), .d(s_210_19), .cin(s_210_18), .o(t_5993), .co(t_5994), .cout(t_5995));
compressor_4_2 u2_2046(.a(s_211_2), .b(s_211_1), .c(s_211_0), .d(t_5980), .cin(t_5983), .o(t_5996), .co(t_5997), .cout(t_5998));
compressor_4_2 u2_2047(.a(s_211_5), .b(s_211_4), .c(s_211_3), .d(t_5986), .cin(t_5989), .o(t_5999), .co(t_6000), .cout(t_6001));
compressor_4_2 u2_2048(.a(s_211_8), .b(s_211_7), .c(s_211_6), .d(t_5992), .cin(t_5995), .o(t_6002), .co(t_6003), .cout(t_6004));
compressor_4_2 u2_2049(.a(s_211_13), .b(s_211_12), .c(s_211_11), .d(s_211_10), .cin(s_211_9), .o(t_6005), .co(t_6006), .cout(t_6007));
compressor_4_2 u2_2050(.a(s_211_18), .b(s_211_17), .c(s_211_16), .d(s_211_15), .cin(s_211_14), .o(t_6008), .co(t_6009), .cout(t_6010));
compressor_4_2 u2_2051(.a(s_211_23), .b(s_211_22), .c(s_211_21), .d(s_211_20), .cin(s_211_19), .o(t_6011), .co(t_6012), .cout(t_6013));
compressor_4_2 u2_2052(.a(s_212_2), .b(s_212_1), .c(s_212_0), .d(t_5998), .cin(t_6001), .o(t_6014), .co(t_6015), .cout(t_6016));
compressor_4_2 u2_2053(.a(s_212_5), .b(s_212_4), .c(s_212_3), .d(t_6004), .cin(t_6007), .o(t_6017), .co(t_6018), .cout(t_6019));
compressor_4_2 u2_2054(.a(s_212_8), .b(s_212_7), .c(s_212_6), .d(t_6010), .cin(t_6013), .o(t_6020), .co(t_6021), .cout(t_6022));
compressor_4_2 u2_2055(.a(s_212_13), .b(s_212_12), .c(s_212_11), .d(s_212_10), .cin(s_212_9), .o(t_6023), .co(t_6024), .cout(t_6025));
compressor_4_2 u2_2056(.a(s_212_18), .b(s_212_17), .c(s_212_16), .d(s_212_15), .cin(s_212_14), .o(t_6026), .co(t_6027), .cout(t_6028));
compressor_3_2 u1_2057(.a(s_212_21), .b(s_212_20), .cin(s_212_19), .o(t_6029), .cout(t_6030));
compressor_4_2 u2_2058(.a(s_213_2), .b(s_213_1), .c(s_213_0), .d(t_6016), .cin(t_6019), .o(t_6031), .co(t_6032), .cout(t_6033));
compressor_4_2 u2_2059(.a(s_213_5), .b(s_213_4), .c(s_213_3), .d(t_6022), .cin(t_6025), .o(t_6034), .co(t_6035), .cout(t_6036));
compressor_4_2 u2_2060(.a(s_213_8), .b(s_213_7), .c(s_213_6), .d(t_6028), .cin(t_6030), .o(t_6037), .co(t_6038), .cout(t_6039));
compressor_4_2 u2_2061(.a(s_213_13), .b(s_213_12), .c(s_213_11), .d(s_213_10), .cin(s_213_9), .o(t_6040), .co(t_6041), .cout(t_6042));
compressor_4_2 u2_2062(.a(s_213_18), .b(s_213_17), .c(s_213_16), .d(s_213_15), .cin(s_213_14), .o(t_6043), .co(t_6044), .cout(t_6045));
compressor_3_2 u1_2063(.a(s_213_21), .b(s_213_20), .cin(s_213_19), .o(t_6046), .cout(t_6047));
compressor_4_2 u2_2064(.a(s_214_2), .b(s_214_1), .c(s_214_0), .d(t_6033), .cin(t_6036), .o(t_6048), .co(t_6049), .cout(t_6050));
compressor_4_2 u2_2065(.a(s_214_5), .b(s_214_4), .c(s_214_3), .d(t_6039), .cin(t_6042), .o(t_6051), .co(t_6052), .cout(t_6053));
compressor_4_2 u2_2066(.a(s_214_8), .b(s_214_7), .c(s_214_6), .d(t_6045), .cin(t_6047), .o(t_6054), .co(t_6055), .cout(t_6056));
compressor_4_2 u2_2067(.a(s_214_13), .b(s_214_12), .c(s_214_11), .d(s_214_10), .cin(s_214_9), .o(t_6057), .co(t_6058), .cout(t_6059));
compressor_4_2 u2_2068(.a(s_214_18), .b(s_214_17), .c(s_214_16), .d(s_214_15), .cin(s_214_14), .o(t_6060), .co(t_6061), .cout(t_6062));
compressor_3_2 u1_2069(.a(s_214_21), .b(s_214_20), .cin(s_214_19), .o(t_6063), .cout(t_6064));
compressor_4_2 u2_2070(.a(s_215_2), .b(s_215_1), .c(s_215_0), .d(t_6050), .cin(t_6053), .o(t_6065), .co(t_6066), .cout(t_6067));
compressor_4_2 u2_2071(.a(s_215_5), .b(s_215_4), .c(s_215_3), .d(t_6056), .cin(t_6059), .o(t_6068), .co(t_6069), .cout(t_6070));
compressor_4_2 u2_2072(.a(s_215_8), .b(s_215_7), .c(s_215_6), .d(t_6062), .cin(t_6064), .o(t_6071), .co(t_6072), .cout(t_6073));
compressor_4_2 u2_2073(.a(s_215_13), .b(s_215_12), .c(s_215_11), .d(s_215_10), .cin(s_215_9), .o(t_6074), .co(t_6075), .cout(t_6076));
compressor_4_2 u2_2074(.a(s_215_18), .b(s_215_17), .c(s_215_16), .d(s_215_15), .cin(s_215_14), .o(t_6077), .co(t_6078), .cout(t_6079));
compressor_3_2 u1_2075(.a(s_215_21), .b(s_215_20), .cin(s_215_19), .o(t_6080), .cout(t_6081));
compressor_4_2 u2_2076(.a(s_216_2), .b(s_216_1), .c(s_216_0), .d(t_6067), .cin(t_6070), .o(t_6082), .co(t_6083), .cout(t_6084));
compressor_4_2 u2_2077(.a(s_216_5), .b(s_216_4), .c(s_216_3), .d(t_6073), .cin(t_6076), .o(t_6085), .co(t_6086), .cout(t_6087));
compressor_4_2 u2_2078(.a(s_216_8), .b(s_216_7), .c(s_216_6), .d(t_6079), .cin(t_6081), .o(t_6088), .co(t_6089), .cout(t_6090));
compressor_4_2 u2_2079(.a(s_216_13), .b(s_216_12), .c(s_216_11), .d(s_216_10), .cin(s_216_9), .o(t_6091), .co(t_6092), .cout(t_6093));
compressor_4_2 u2_2080(.a(s_216_18), .b(s_216_17), .c(s_216_16), .d(s_216_15), .cin(s_216_14), .o(t_6094), .co(t_6095), .cout(t_6096));
half_adder u0_2081(.a(s_216_20), .b(s_216_19), .o(t_6097), .cout(t_6098));
compressor_4_2 u2_2082(.a(s_217_2), .b(s_217_1), .c(s_217_0), .d(t_6084), .cin(t_6087), .o(t_6099), .co(t_6100), .cout(t_6101));
compressor_4_2 u2_2083(.a(s_217_5), .b(s_217_4), .c(s_217_3), .d(t_6090), .cin(t_6093), .o(t_6102), .co(t_6103), .cout(t_6104));
compressor_4_2 u2_2084(.a(s_217_8), .b(s_217_7), .c(s_217_6), .d(t_6096), .cin(t_6098), .o(t_6105), .co(t_6106), .cout(t_6107));
compressor_4_2 u2_2085(.a(s_217_13), .b(s_217_12), .c(s_217_11), .d(s_217_10), .cin(s_217_9), .o(t_6108), .co(t_6109), .cout(t_6110));
compressor_4_2 u2_2086(.a(s_217_18), .b(s_217_17), .c(s_217_16), .d(s_217_15), .cin(s_217_14), .o(t_6111), .co(t_6112), .cout(t_6113));
half_adder u0_2087(.a(s_217_20), .b(s_217_19), .o(t_6114), .cout(t_6115));
compressor_4_2 u2_2088(.a(s_218_2), .b(s_218_1), .c(s_218_0), .d(t_6101), .cin(t_6104), .o(t_6116), .co(t_6117), .cout(t_6118));
compressor_4_2 u2_2089(.a(s_218_5), .b(s_218_4), .c(s_218_3), .d(t_6107), .cin(t_6110), .o(t_6119), .co(t_6120), .cout(t_6121));
compressor_4_2 u2_2090(.a(s_218_8), .b(s_218_7), .c(s_218_6), .d(t_6113), .cin(t_6115), .o(t_6122), .co(t_6123), .cout(t_6124));
compressor_4_2 u2_2091(.a(s_218_13), .b(s_218_12), .c(s_218_11), .d(s_218_10), .cin(s_218_9), .o(t_6125), .co(t_6126), .cout(t_6127));
compressor_4_2 u2_2092(.a(s_218_18), .b(s_218_17), .c(s_218_16), .d(s_218_15), .cin(s_218_14), .o(t_6128), .co(t_6129), .cout(t_6130));
compressor_4_2 u2_2093(.a(s_219_2), .b(s_219_1), .c(s_219_0), .d(t_6118), .cin(t_6121), .o(t_6131), .co(t_6132), .cout(t_6133));
compressor_4_2 u2_2094(.a(s_219_5), .b(s_219_4), .c(s_219_3), .d(t_6124), .cin(t_6127), .o(t_6134), .co(t_6135), .cout(t_6136));
compressor_4_2 u2_2095(.a(s_219_9), .b(s_219_8), .c(s_219_7), .d(s_219_6), .cin(t_6130), .o(t_6137), .co(t_6138), .cout(t_6139));
compressor_4_2 u2_2096(.a(s_219_14), .b(s_219_13), .c(s_219_12), .d(s_219_11), .cin(s_219_10), .o(t_6140), .co(t_6141), .cout(t_6142));
compressor_4_2 u2_2097(.a(s_219_19), .b(s_219_18), .c(s_219_17), .d(s_219_16), .cin(s_219_15), .o(t_6143), .co(t_6144), .cout(t_6145));
compressor_4_2 u2_2098(.a(s_220_2), .b(s_220_1), .c(s_220_0), .d(t_6133), .cin(t_6136), .o(t_6146), .co(t_6147), .cout(t_6148));
compressor_4_2 u2_2099(.a(s_220_5), .b(s_220_4), .c(s_220_3), .d(t_6139), .cin(t_6142), .o(t_6149), .co(t_6150), .cout(t_6151));
compressor_4_2 u2_2100(.a(s_220_9), .b(s_220_8), .c(s_220_7), .d(s_220_6), .cin(t_6145), .o(t_6152), .co(t_6153), .cout(t_6154));
compressor_4_2 u2_2101(.a(s_220_14), .b(s_220_13), .c(s_220_12), .d(s_220_11), .cin(s_220_10), .o(t_6155), .co(t_6156), .cout(t_6157));
compressor_3_2 u1_2102(.a(s_220_17), .b(s_220_16), .cin(s_220_15), .o(t_6158), .cout(t_6159));
compressor_4_2 u2_2103(.a(s_221_2), .b(s_221_1), .c(s_221_0), .d(t_6148), .cin(t_6151), .o(t_6160), .co(t_6161), .cout(t_6162));
compressor_4_2 u2_2104(.a(s_221_5), .b(s_221_4), .c(s_221_3), .d(t_6154), .cin(t_6157), .o(t_6163), .co(t_6164), .cout(t_6165));
compressor_4_2 u2_2105(.a(s_221_9), .b(s_221_8), .c(s_221_7), .d(s_221_6), .cin(t_6159), .o(t_6166), .co(t_6167), .cout(t_6168));
compressor_4_2 u2_2106(.a(s_221_14), .b(s_221_13), .c(s_221_12), .d(s_221_11), .cin(s_221_10), .o(t_6169), .co(t_6170), .cout(t_6171));
compressor_3_2 u1_2107(.a(s_221_17), .b(s_221_16), .cin(s_221_15), .o(t_6172), .cout(t_6173));
compressor_4_2 u2_2108(.a(s_222_2), .b(s_222_1), .c(s_222_0), .d(t_6162), .cin(t_6165), .o(t_6174), .co(t_6175), .cout(t_6176));
compressor_4_2 u2_2109(.a(s_222_5), .b(s_222_4), .c(s_222_3), .d(t_6168), .cin(t_6171), .o(t_6177), .co(t_6178), .cout(t_6179));
compressor_4_2 u2_2110(.a(s_222_9), .b(s_222_8), .c(s_222_7), .d(s_222_6), .cin(t_6173), .o(t_6180), .co(t_6181), .cout(t_6182));
compressor_4_2 u2_2111(.a(s_222_14), .b(s_222_13), .c(s_222_12), .d(s_222_11), .cin(s_222_10), .o(t_6183), .co(t_6184), .cout(t_6185));
compressor_3_2 u1_2112(.a(s_222_17), .b(s_222_16), .cin(s_222_15), .o(t_6186), .cout(t_6187));
compressor_4_2 u2_2113(.a(s_223_2), .b(s_223_1), .c(s_223_0), .d(t_6176), .cin(t_6179), .o(t_6188), .co(t_6189), .cout(t_6190));
compressor_4_2 u2_2114(.a(s_223_5), .b(s_223_4), .c(s_223_3), .d(t_6182), .cin(t_6185), .o(t_6191), .co(t_6192), .cout(t_6193));
compressor_4_2 u2_2115(.a(s_223_9), .b(s_223_8), .c(s_223_7), .d(s_223_6), .cin(t_6187), .o(t_6194), .co(t_6195), .cout(t_6196));
compressor_4_2 u2_2116(.a(s_223_14), .b(s_223_13), .c(s_223_12), .d(s_223_11), .cin(s_223_10), .o(t_6197), .co(t_6198), .cout(t_6199));
compressor_3_2 u1_2117(.a(s_223_17), .b(s_223_16), .cin(s_223_15), .o(t_6200), .cout(t_6201));
compressor_4_2 u2_2118(.a(s_224_2), .b(s_224_1), .c(s_224_0), .d(t_6190), .cin(t_6193), .o(t_6202), .co(t_6203), .cout(t_6204));
compressor_4_2 u2_2119(.a(s_224_5), .b(s_224_4), .c(s_224_3), .d(t_6196), .cin(t_6199), .o(t_6205), .co(t_6206), .cout(t_6207));
compressor_4_2 u2_2120(.a(s_224_9), .b(s_224_8), .c(s_224_7), .d(s_224_6), .cin(t_6201), .o(t_6208), .co(t_6209), .cout(t_6210));
compressor_4_2 u2_2121(.a(s_224_14), .b(s_224_13), .c(s_224_12), .d(s_224_11), .cin(s_224_10), .o(t_6211), .co(t_6212), .cout(t_6213));
half_adder u0_2122(.a(s_224_16), .b(s_224_15), .o(t_6214), .cout(t_6215));
compressor_4_2 u2_2123(.a(s_225_2), .b(s_225_1), .c(s_225_0), .d(t_6204), .cin(t_6207), .o(t_6216), .co(t_6217), .cout(t_6218));
compressor_4_2 u2_2124(.a(s_225_5), .b(s_225_4), .c(s_225_3), .d(t_6210), .cin(t_6213), .o(t_6219), .co(t_6220), .cout(t_6221));
compressor_4_2 u2_2125(.a(s_225_9), .b(s_225_8), .c(s_225_7), .d(s_225_6), .cin(t_6215), .o(t_6222), .co(t_6223), .cout(t_6224));
compressor_4_2 u2_2126(.a(s_225_14), .b(s_225_13), .c(s_225_12), .d(s_225_11), .cin(s_225_10), .o(t_6225), .co(t_6226), .cout(t_6227));
half_adder u0_2127(.a(s_225_16), .b(s_225_15), .o(t_6228), .cout(t_6229));
compressor_4_2 u2_2128(.a(s_226_2), .b(s_226_1), .c(s_226_0), .d(t_6218), .cin(t_6221), .o(t_6230), .co(t_6231), .cout(t_6232));
compressor_4_2 u2_2129(.a(s_226_5), .b(s_226_4), .c(s_226_3), .d(t_6224), .cin(t_6227), .o(t_6233), .co(t_6234), .cout(t_6235));
compressor_4_2 u2_2130(.a(s_226_9), .b(s_226_8), .c(s_226_7), .d(s_226_6), .cin(t_6229), .o(t_6236), .co(t_6237), .cout(t_6238));
compressor_4_2 u2_2131(.a(s_226_14), .b(s_226_13), .c(s_226_12), .d(s_226_11), .cin(s_226_10), .o(t_6239), .co(t_6240), .cout(t_6241));
compressor_4_2 u2_2132(.a(s_227_2), .b(s_227_1), .c(s_227_0), .d(t_6232), .cin(t_6235), .o(t_6242), .co(t_6243), .cout(t_6244));
compressor_4_2 u2_2133(.a(s_227_5), .b(s_227_4), .c(s_227_3), .d(t_6238), .cin(t_6241), .o(t_6245), .co(t_6246), .cout(t_6247));
compressor_4_2 u2_2134(.a(s_227_10), .b(s_227_9), .c(s_227_8), .d(s_227_7), .cin(s_227_6), .o(t_6248), .co(t_6249), .cout(t_6250));
compressor_4_2 u2_2135(.a(s_227_15), .b(s_227_14), .c(s_227_13), .d(s_227_12), .cin(s_227_11), .o(t_6251), .co(t_6252), .cout(t_6253));
compressor_4_2 u2_2136(.a(s_228_2), .b(s_228_1), .c(s_228_0), .d(t_6244), .cin(t_6247), .o(t_6254), .co(t_6255), .cout(t_6256));
compressor_4_2 u2_2137(.a(s_228_5), .b(s_228_4), .c(s_228_3), .d(t_6250), .cin(t_6253), .o(t_6257), .co(t_6258), .cout(t_6259));
compressor_4_2 u2_2138(.a(s_228_10), .b(s_228_9), .c(s_228_8), .d(s_228_7), .cin(s_228_6), .o(t_6260), .co(t_6261), .cout(t_6262));
compressor_3_2 u1_2139(.a(s_228_13), .b(s_228_12), .cin(s_228_11), .o(t_6263), .cout(t_6264));
compressor_4_2 u2_2140(.a(s_229_2), .b(s_229_1), .c(s_229_0), .d(t_6256), .cin(t_6259), .o(t_6265), .co(t_6266), .cout(t_6267));
compressor_4_2 u2_2141(.a(s_229_5), .b(s_229_4), .c(s_229_3), .d(t_6262), .cin(t_6264), .o(t_6268), .co(t_6269), .cout(t_6270));
compressor_4_2 u2_2142(.a(s_229_10), .b(s_229_9), .c(s_229_8), .d(s_229_7), .cin(s_229_6), .o(t_6271), .co(t_6272), .cout(t_6273));
compressor_3_2 u1_2143(.a(s_229_13), .b(s_229_12), .cin(s_229_11), .o(t_6274), .cout(t_6275));
compressor_4_2 u2_2144(.a(s_230_2), .b(s_230_1), .c(s_230_0), .d(t_6267), .cin(t_6270), .o(t_6276), .co(t_6277), .cout(t_6278));
compressor_4_2 u2_2145(.a(s_230_5), .b(s_230_4), .c(s_230_3), .d(t_6273), .cin(t_6275), .o(t_6279), .co(t_6280), .cout(t_6281));
compressor_4_2 u2_2146(.a(s_230_10), .b(s_230_9), .c(s_230_8), .d(s_230_7), .cin(s_230_6), .o(t_6282), .co(t_6283), .cout(t_6284));
compressor_3_2 u1_2147(.a(s_230_13), .b(s_230_12), .cin(s_230_11), .o(t_6285), .cout(t_6286));
compressor_4_2 u2_2148(.a(s_231_2), .b(s_231_1), .c(s_231_0), .d(t_6278), .cin(t_6281), .o(t_6287), .co(t_6288), .cout(t_6289));
compressor_4_2 u2_2149(.a(s_231_5), .b(s_231_4), .c(s_231_3), .d(t_6284), .cin(t_6286), .o(t_6290), .co(t_6291), .cout(t_6292));
compressor_4_2 u2_2150(.a(s_231_10), .b(s_231_9), .c(s_231_8), .d(s_231_7), .cin(s_231_6), .o(t_6293), .co(t_6294), .cout(t_6295));
compressor_3_2 u1_2151(.a(s_231_13), .b(s_231_12), .cin(s_231_11), .o(t_6296), .cout(t_6297));
compressor_4_2 u2_2152(.a(s_232_2), .b(s_232_1), .c(s_232_0), .d(t_6289), .cin(t_6292), .o(t_6298), .co(t_6299), .cout(t_6300));
compressor_4_2 u2_2153(.a(s_232_5), .b(s_232_4), .c(s_232_3), .d(t_6295), .cin(t_6297), .o(t_6301), .co(t_6302), .cout(t_6303));
compressor_4_2 u2_2154(.a(s_232_10), .b(s_232_9), .c(s_232_8), .d(s_232_7), .cin(s_232_6), .o(t_6304), .co(t_6305), .cout(t_6306));
half_adder u0_2155(.a(s_232_12), .b(s_232_11), .o(t_6307), .cout(t_6308));
compressor_4_2 u2_2156(.a(s_233_2), .b(s_233_1), .c(s_233_0), .d(t_6300), .cin(t_6303), .o(t_6309), .co(t_6310), .cout(t_6311));
compressor_4_2 u2_2157(.a(s_233_5), .b(s_233_4), .c(s_233_3), .d(t_6306), .cin(t_6308), .o(t_6312), .co(t_6313), .cout(t_6314));
compressor_4_2 u2_2158(.a(s_233_10), .b(s_233_9), .c(s_233_8), .d(s_233_7), .cin(s_233_6), .o(t_6315), .co(t_6316), .cout(t_6317));
half_adder u0_2159(.a(s_233_12), .b(s_233_11), .o(t_6318), .cout(t_6319));
compressor_4_2 u2_2160(.a(s_234_2), .b(s_234_1), .c(s_234_0), .d(t_6311), .cin(t_6314), .o(t_6320), .co(t_6321), .cout(t_6322));
compressor_4_2 u2_2161(.a(s_234_5), .b(s_234_4), .c(s_234_3), .d(t_6317), .cin(t_6319), .o(t_6323), .co(t_6324), .cout(t_6325));
compressor_4_2 u2_2162(.a(s_234_10), .b(s_234_9), .c(s_234_8), .d(s_234_7), .cin(s_234_6), .o(t_6326), .co(t_6327), .cout(t_6328));
compressor_4_2 u2_2163(.a(s_235_2), .b(s_235_1), .c(s_235_0), .d(t_6322), .cin(t_6325), .o(t_6329), .co(t_6330), .cout(t_6331));
compressor_4_2 u2_2164(.a(s_235_6), .b(s_235_5), .c(s_235_4), .d(s_235_3), .cin(t_6328), .o(t_6332), .co(t_6333), .cout(t_6334));
compressor_4_2 u2_2165(.a(s_235_11), .b(s_235_10), .c(s_235_9), .d(s_235_8), .cin(s_235_7), .o(t_6335), .co(t_6336), .cout(t_6337));
compressor_4_2 u2_2166(.a(s_236_2), .b(s_236_1), .c(s_236_0), .d(t_6331), .cin(t_6334), .o(t_6338), .co(t_6339), .cout(t_6340));
compressor_4_2 u2_2167(.a(s_236_6), .b(s_236_5), .c(s_236_4), .d(s_236_3), .cin(t_6337), .o(t_6341), .co(t_6342), .cout(t_6343));
compressor_3_2 u1_2168(.a(s_236_9), .b(s_236_8), .cin(s_236_7), .o(t_6344), .cout(t_6345));
compressor_4_2 u2_2169(.a(s_237_2), .b(s_237_1), .c(s_237_0), .d(t_6340), .cin(t_6343), .o(t_6346), .co(t_6347), .cout(t_6348));
compressor_4_2 u2_2170(.a(s_237_6), .b(s_237_5), .c(s_237_4), .d(s_237_3), .cin(t_6345), .o(t_6349), .co(t_6350), .cout(t_6351));
compressor_3_2 u1_2171(.a(s_237_9), .b(s_237_8), .cin(s_237_7), .o(t_6352), .cout(t_6353));
compressor_4_2 u2_2172(.a(s_238_2), .b(s_238_1), .c(s_238_0), .d(t_6348), .cin(t_6351), .o(t_6354), .co(t_6355), .cout(t_6356));
compressor_4_2 u2_2173(.a(s_238_6), .b(s_238_5), .c(s_238_4), .d(s_238_3), .cin(t_6353), .o(t_6357), .co(t_6358), .cout(t_6359));
compressor_3_2 u1_2174(.a(s_238_9), .b(s_238_8), .cin(s_238_7), .o(t_6360), .cout(t_6361));
compressor_4_2 u2_2175(.a(s_239_2), .b(s_239_1), .c(s_239_0), .d(t_6356), .cin(t_6359), .o(t_6362), .co(t_6363), .cout(t_6364));
compressor_4_2 u2_2176(.a(s_239_6), .b(s_239_5), .c(s_239_4), .d(s_239_3), .cin(t_6361), .o(t_6365), .co(t_6366), .cout(t_6367));
compressor_3_2 u1_2177(.a(s_239_9), .b(s_239_8), .cin(s_239_7), .o(t_6368), .cout(t_6369));
compressor_4_2 u2_2178(.a(s_240_2), .b(s_240_1), .c(s_240_0), .d(t_6364), .cin(t_6367), .o(t_6370), .co(t_6371), .cout(t_6372));
compressor_4_2 u2_2179(.a(s_240_6), .b(s_240_5), .c(s_240_4), .d(s_240_3), .cin(t_6369), .o(t_6373), .co(t_6374), .cout(t_6375));
half_adder u0_2180(.a(s_240_8), .b(s_240_7), .o(t_6376), .cout(t_6377));
compressor_4_2 u2_2181(.a(s_241_2), .b(s_241_1), .c(s_241_0), .d(t_6372), .cin(t_6375), .o(t_6378), .co(t_6379), .cout(t_6380));
compressor_4_2 u2_2182(.a(s_241_6), .b(s_241_5), .c(s_241_4), .d(s_241_3), .cin(t_6377), .o(t_6381), .co(t_6382), .cout(t_6383));
half_adder u0_2183(.a(s_241_8), .b(s_241_7), .o(t_6384), .cout(t_6385));
compressor_4_2 u2_2184(.a(s_242_2), .b(s_242_1), .c(s_242_0), .d(t_6380), .cin(t_6383), .o(t_6386), .co(t_6387), .cout(t_6388));
compressor_4_2 u2_2185(.a(s_242_6), .b(s_242_5), .c(s_242_4), .d(s_242_3), .cin(t_6385), .o(t_6389), .co(t_6390), .cout(t_6391));
compressor_4_2 u2_2186(.a(s_243_2), .b(s_243_1), .c(s_243_0), .d(t_6388), .cin(t_6391), .o(t_6392), .co(t_6393), .cout(t_6394));
compressor_4_2 u2_2187(.a(s_243_7), .b(s_243_6), .c(s_243_5), .d(s_243_4), .cin(s_243_3), .o(t_6395), .co(t_6396), .cout(t_6397));
compressor_4_2 u2_2188(.a(s_244_2), .b(s_244_1), .c(s_244_0), .d(t_6394), .cin(t_6397), .o(t_6398), .co(t_6399), .cout(t_6400));
compressor_3_2 u1_2189(.a(s_244_5), .b(s_244_4), .cin(s_244_3), .o(t_6401), .cout(t_6402));
compressor_4_2 u2_2190(.a(s_245_2), .b(s_245_1), .c(s_245_0), .d(t_6400), .cin(t_6402), .o(t_6403), .co(t_6404), .cout(t_6405));
compressor_3_2 u1_2191(.a(s_245_5), .b(s_245_4), .cin(s_245_3), .o(t_6406), .cout(t_6407));
compressor_4_2 u2_2192(.a(s_246_2), .b(s_246_1), .c(s_246_0), .d(t_6405), .cin(t_6407), .o(t_6408), .co(t_6409), .cout(t_6410));
compressor_3_2 u1_2193(.a(s_246_5), .b(s_246_4), .cin(s_246_3), .o(t_6411), .cout(t_6412));
compressor_4_2 u2_2194(.a(s_247_2), .b(s_247_1), .c(s_247_0), .d(t_6410), .cin(t_6412), .o(t_6413), .co(t_6414), .cout(t_6415));
compressor_3_2 u1_2195(.a(s_247_5), .b(s_247_4), .cin(s_247_3), .o(t_6416), .cout(t_6417));
compressor_4_2 u2_2196(.a(s_248_2), .b(s_248_1), .c(s_248_0), .d(t_6415), .cin(t_6417), .o(t_6418), .co(t_6419), .cout(t_6420));
half_adder u0_2197(.a(s_248_4), .b(s_248_3), .o(t_6421), .cout(t_6422));
compressor_4_2 u2_2198(.a(s_249_2), .b(s_249_1), .c(s_249_0), .d(t_6420), .cin(t_6422), .o(t_6423), .co(t_6424), .cout(t_6425));
half_adder u0_2199(.a(s_249_4), .b(s_249_3), .o(t_6426), .cout(t_6427));
compressor_4_2 u2_2200(.a(s_250_2), .b(s_250_1), .c(s_250_0), .d(t_6425), .cin(t_6427), .o(t_6428), .co(t_6429), .cout(t_6430));
compressor_4_2 u2_2201(.a(s_251_3), .b(s_251_2), .c(s_251_1), .d(s_251_0), .cin(t_6430), .o(t_6431), .co(t_6432), .cout(t_6433));
compressor_3_2 u1_2202(.a(s_252_1), .b(s_252_0), .cin(t_6433), .o(t_6434), .cout(t_6435));
compressor_3_2 u1_2203(.a(s_253_2), .b(s_253_1), .cin(s_253_0), .o(t_6436), .cout(t_6437));
half_adder u0_2204(.a(s_254_1), .b(s_254_0), .o(t_6438), .cout(t_6439));
half_adder u0_2205(.a(s_255_1), .b(s_255_0), .o(t_6440), .cout());

/* u0_2206 Output nets */
wire t_6441,   t_6442;
/* u0_2207 Output nets */
wire t_6443,   t_6444;
/* u1_2208 Output nets */
wire t_6445,   t_6446;
/* u0_2209 Output nets */
wire t_6447,   t_6448;
/* u0_2210 Output nets */
wire t_6449,   t_6450;
/* u1_2211 Output nets */
wire t_6451,   t_6452;
/* u1_2212 Output nets */
wire t_6453,   t_6454;
/* u2_2213 Output nets */
wire t_6455,   t_6456,   t_6457;
/* u1_2214 Output nets */
wire t_6458,   t_6459;
/* u1_2215 Output nets */
wire t_6460,   t_6461;
/* u2_2216 Output nets */
wire t_6462,   t_6463,   t_6464;
/* u2_2217 Output nets */
wire t_6465,   t_6466,   t_6467;
/* u2_2218 Output nets */
wire t_6468,   t_6469,   t_6470;
/* u2_2219 Output nets */
wire t_6471,   t_6472,   t_6473;
/* u2_2220 Output nets */
wire t_6474,   t_6475,   t_6476;
/* u2_2221 Output nets */
wire t_6477,   t_6478,   t_6479;
/* u0_2222 Output nets */
wire t_6480,   t_6481;
/* u2_2223 Output nets */
wire t_6482,   t_6483,   t_6484;
/* u0_2224 Output nets */
wire t_6485,   t_6486;
/* u2_2225 Output nets */
wire t_6487,   t_6488,   t_6489;
/* u0_2226 Output nets */
wire t_6490,   t_6491;
/* u2_2227 Output nets */
wire t_6492,   t_6493,   t_6494;
/* u1_2228 Output nets */
wire t_6495,   t_6496;
/* u2_2229 Output nets */
wire t_6497,   t_6498,   t_6499;
/* u1_2230 Output nets */
wire t_6500,   t_6501;
/* u2_2231 Output nets */
wire t_6502,   t_6503,   t_6504;
/* u1_2232 Output nets */
wire t_6505,   t_6506;
/* u2_2233 Output nets */
wire t_6507,   t_6508,   t_6509;
/* u1_2234 Output nets */
wire t_6510,   t_6511;
/* u2_2235 Output nets */
wire t_6512,   t_6513,   t_6514;
/* u1_2236 Output nets */
wire t_6515,   t_6516;
/* u2_2237 Output nets */
wire t_6517,   t_6518,   t_6519;
/* u2_2238 Output nets */
wire t_6520,   t_6521,   t_6522;
/* u2_2239 Output nets */
wire t_6523,   t_6524,   t_6525;
/* u1_2240 Output nets */
wire t_6526,   t_6527;
/* u2_2241 Output nets */
wire t_6528,   t_6529,   t_6530;
/* u1_2242 Output nets */
wire t_6531,   t_6532;
/* u2_2243 Output nets */
wire t_6533,   t_6534,   t_6535;
/* u2_2244 Output nets */
wire t_6536,   t_6537,   t_6538;
/* u2_2245 Output nets */
wire t_6539,   t_6540,   t_6541;
/* u2_2246 Output nets */
wire t_6542,   t_6543,   t_6544;
/* u2_2247 Output nets */
wire t_6545,   t_6546,   t_6547;
/* u2_2248 Output nets */
wire t_6548,   t_6549,   t_6550;
/* u2_2249 Output nets */
wire t_6551,   t_6552,   t_6553;
/* u2_2250 Output nets */
wire t_6554,   t_6555,   t_6556;
/* u2_2251 Output nets */
wire t_6557,   t_6558,   t_6559;
/* u2_2252 Output nets */
wire t_6560,   t_6561,   t_6562;
/* u2_2253 Output nets */
wire t_6563,   t_6564,   t_6565;
/* u2_2254 Output nets */
wire t_6566,   t_6567,   t_6568;
/* u0_2255 Output nets */
wire t_6569,   t_6570;
/* u2_2256 Output nets */
wire t_6571,   t_6572,   t_6573;
/* u2_2257 Output nets */
wire t_6574,   t_6575,   t_6576;
/* u0_2258 Output nets */
wire t_6577,   t_6578;
/* u2_2259 Output nets */
wire t_6579,   t_6580,   t_6581;
/* u2_2260 Output nets */
wire t_6582,   t_6583,   t_6584;
/* u0_2261 Output nets */
wire t_6585,   t_6586;
/* u2_2262 Output nets */
wire t_6587,   t_6588,   t_6589;
/* u2_2263 Output nets */
wire t_6590,   t_6591,   t_6592;
/* u1_2264 Output nets */
wire t_6593,   t_6594;
/* u2_2265 Output nets */
wire t_6595,   t_6596,   t_6597;
/* u2_2266 Output nets */
wire t_6598,   t_6599,   t_6600;
/* u1_2267 Output nets */
wire t_6601,   t_6602;
/* u2_2268 Output nets */
wire t_6603,   t_6604,   t_6605;
/* u2_2269 Output nets */
wire t_6606,   t_6607,   t_6608;
/* u1_2270 Output nets */
wire t_6609,   t_6610;
/* u2_2271 Output nets */
wire t_6611,   t_6612,   t_6613;
/* u2_2272 Output nets */
wire t_6614,   t_6615,   t_6616;
/* u1_2273 Output nets */
wire t_6617,   t_6618;
/* u2_2274 Output nets */
wire t_6619,   t_6620,   t_6621;
/* u2_2275 Output nets */
wire t_6622,   t_6623,   t_6624;
/* u1_2276 Output nets */
wire t_6625,   t_6626;
/* u2_2277 Output nets */
wire t_6627,   t_6628,   t_6629;
/* u2_2278 Output nets */
wire t_6630,   t_6631,   t_6632;
/* u2_2279 Output nets */
wire t_6633,   t_6634,   t_6635;
/* u2_2280 Output nets */
wire t_6636,   t_6637,   t_6638;
/* u2_2281 Output nets */
wire t_6639,   t_6640,   t_6641;
/* u1_2282 Output nets */
wire t_6642,   t_6643;
/* u2_2283 Output nets */
wire t_6644,   t_6645,   t_6646;
/* u2_2284 Output nets */
wire t_6647,   t_6648,   t_6649;
/* u1_2285 Output nets */
wire t_6650,   t_6651;
/* u2_2286 Output nets */
wire t_6652,   t_6653,   t_6654;
/* u2_2287 Output nets */
wire t_6655,   t_6656,   t_6657;
/* u2_2288 Output nets */
wire t_6658,   t_6659,   t_6660;
/* u2_2289 Output nets */
wire t_6661,   t_6662,   t_6663;
/* u2_2290 Output nets */
wire t_6664,   t_6665,   t_6666;
/* u2_2291 Output nets */
wire t_6667,   t_6668,   t_6669;
/* u2_2292 Output nets */
wire t_6670,   t_6671,   t_6672;
/* u2_2293 Output nets */
wire t_6673,   t_6674,   t_6675;
/* u2_2294 Output nets */
wire t_6676,   t_6677,   t_6678;
/* u2_2295 Output nets */
wire t_6679,   t_6680,   t_6681;
/* u2_2296 Output nets */
wire t_6682,   t_6683,   t_6684;
/* u2_2297 Output nets */
wire t_6685,   t_6686,   t_6687;
/* u2_2298 Output nets */
wire t_6688,   t_6689,   t_6690;
/* u2_2299 Output nets */
wire t_6691,   t_6692,   t_6693;
/* u2_2300 Output nets */
wire t_6694,   t_6695,   t_6696;
/* u2_2301 Output nets */
wire t_6697,   t_6698,   t_6699;
/* u2_2302 Output nets */
wire t_6700,   t_6701,   t_6702;
/* u2_2303 Output nets */
wire t_6703,   t_6704,   t_6705;
/* u0_2304 Output nets */
wire t_6706,   t_6707;
/* u2_2305 Output nets */
wire t_6708,   t_6709,   t_6710;
/* u2_2306 Output nets */
wire t_6711,   t_6712,   t_6713;
/* u2_2307 Output nets */
wire t_6714,   t_6715,   t_6716;
/* u0_2308 Output nets */
wire t_6717,   t_6718;
/* u2_2309 Output nets */
wire t_6719,   t_6720,   t_6721;
/* u2_2310 Output nets */
wire t_6722,   t_6723,   t_6724;
/* u2_2311 Output nets */
wire t_6725,   t_6726,   t_6727;
/* u0_2312 Output nets */
wire t_6728,   t_6729;
/* u2_2313 Output nets */
wire t_6730,   t_6731,   t_6732;
/* u2_2314 Output nets */
wire t_6733,   t_6734,   t_6735;
/* u2_2315 Output nets */
wire t_6736,   t_6737,   t_6738;
/* u1_2316 Output nets */
wire t_6739,   t_6740;
/* u2_2317 Output nets */
wire t_6741,   t_6742,   t_6743;
/* u2_2318 Output nets */
wire t_6744,   t_6745,   t_6746;
/* u2_2319 Output nets */
wire t_6747,   t_6748,   t_6749;
/* u1_2320 Output nets */
wire t_6750,   t_6751;
/* u2_2321 Output nets */
wire t_6752,   t_6753,   t_6754;
/* u2_2322 Output nets */
wire t_6755,   t_6756,   t_6757;
/* u2_2323 Output nets */
wire t_6758,   t_6759,   t_6760;
/* u1_2324 Output nets */
wire t_6761,   t_6762;
/* u2_2325 Output nets */
wire t_6763,   t_6764,   t_6765;
/* u2_2326 Output nets */
wire t_6766,   t_6767,   t_6768;
/* u2_2327 Output nets */
wire t_6769,   t_6770,   t_6771;
/* u1_2328 Output nets */
wire t_6772,   t_6773;
/* u2_2329 Output nets */
wire t_6774,   t_6775,   t_6776;
/* u2_2330 Output nets */
wire t_6777,   t_6778,   t_6779;
/* u2_2331 Output nets */
wire t_6780,   t_6781,   t_6782;
/* u1_2332 Output nets */
wire t_6783,   t_6784;
/* u2_2333 Output nets */
wire t_6785,   t_6786,   t_6787;
/* u2_2334 Output nets */
wire t_6788,   t_6789,   t_6790;
/* u2_2335 Output nets */
wire t_6791,   t_6792,   t_6793;
/* u2_2336 Output nets */
wire t_6794,   t_6795,   t_6796;
/* u2_2337 Output nets */
wire t_6797,   t_6798,   t_6799;
/* u2_2338 Output nets */
wire t_6800,   t_6801,   t_6802;
/* u2_2339 Output nets */
wire t_6803,   t_6804,   t_6805;
/* u1_2340 Output nets */
wire t_6806,   t_6807;
/* u2_2341 Output nets */
wire t_6808,   t_6809,   t_6810;
/* u2_2342 Output nets */
wire t_6811,   t_6812,   t_6813;
/* u2_2343 Output nets */
wire t_6814,   t_6815,   t_6816;
/* u1_2344 Output nets */
wire t_6817,   t_6818;
/* u2_2345 Output nets */
wire t_6819,   t_6820,   t_6821;
/* u2_2346 Output nets */
wire t_6822,   t_6823,   t_6824;
/* u2_2347 Output nets */
wire t_6825,   t_6826,   t_6827;
/* u2_2348 Output nets */
wire t_6828,   t_6829,   t_6830;
/* u2_2349 Output nets */
wire t_6831,   t_6832,   t_6833;
/* u2_2350 Output nets */
wire t_6834,   t_6835,   t_6836;
/* u2_2351 Output nets */
wire t_6837,   t_6838,   t_6839;
/* u2_2352 Output nets */
wire t_6840,   t_6841,   t_6842;
/* u2_2353 Output nets */
wire t_6843,   t_6844,   t_6845;
/* u2_2354 Output nets */
wire t_6846,   t_6847,   t_6848;
/* u2_2355 Output nets */
wire t_6849,   t_6850,   t_6851;
/* u2_2356 Output nets */
wire t_6852,   t_6853,   t_6854;
/* u2_2357 Output nets */
wire t_6855,   t_6856,   t_6857;
/* u2_2358 Output nets */
wire t_6858,   t_6859,   t_6860;
/* u2_2359 Output nets */
wire t_6861,   t_6862,   t_6863;
/* u2_2360 Output nets */
wire t_6864,   t_6865,   t_6866;
/* u2_2361 Output nets */
wire t_6867,   t_6868,   t_6869;
/* u2_2362 Output nets */
wire t_6870,   t_6871,   t_6872;
/* u2_2363 Output nets */
wire t_6873,   t_6874,   t_6875;
/* u2_2364 Output nets */
wire t_6876,   t_6877,   t_6878;
/* u2_2365 Output nets */
wire t_6879,   t_6880,   t_6881;
/* u2_2366 Output nets */
wire t_6882,   t_6883,   t_6884;
/* u2_2367 Output nets */
wire t_6885,   t_6886,   t_6887;
/* u2_2368 Output nets */
wire t_6888,   t_6889,   t_6890;
/* u0_2369 Output nets */
wire t_6891,   t_6892;
/* u2_2370 Output nets */
wire t_6893,   t_6894,   t_6895;
/* u2_2371 Output nets */
wire t_6896,   t_6897,   t_6898;
/* u2_2372 Output nets */
wire t_6899,   t_6900,   t_6901;
/* u2_2373 Output nets */
wire t_6902,   t_6903,   t_6904;
/* u0_2374 Output nets */
wire t_6905,   t_6906;
/* u2_2375 Output nets */
wire t_6907,   t_6908,   t_6909;
/* u2_2376 Output nets */
wire t_6910,   t_6911,   t_6912;
/* u2_2377 Output nets */
wire t_6913,   t_6914,   t_6915;
/* u2_2378 Output nets */
wire t_6916,   t_6917,   t_6918;
/* u0_2379 Output nets */
wire t_6919,   t_6920;
/* u2_2380 Output nets */
wire t_6921,   t_6922,   t_6923;
/* u2_2381 Output nets */
wire t_6924,   t_6925,   t_6926;
/* u2_2382 Output nets */
wire t_6927,   t_6928,   t_6929;
/* u2_2383 Output nets */
wire t_6930,   t_6931,   t_6932;
/* u1_2384 Output nets */
wire t_6933,   t_6934;
/* u2_2385 Output nets */
wire t_6935,   t_6936,   t_6937;
/* u2_2386 Output nets */
wire t_6938,   t_6939,   t_6940;
/* u2_2387 Output nets */
wire t_6941,   t_6942,   t_6943;
/* u2_2388 Output nets */
wire t_6944,   t_6945,   t_6946;
/* u1_2389 Output nets */
wire t_6947,   t_6948;
/* u2_2390 Output nets */
wire t_6949,   t_6950,   t_6951;
/* u2_2391 Output nets */
wire t_6952,   t_6953,   t_6954;
/* u2_2392 Output nets */
wire t_6955,   t_6956,   t_6957;
/* u2_2393 Output nets */
wire t_6958,   t_6959,   t_6960;
/* u1_2394 Output nets */
wire t_6961,   t_6962;
/* u2_2395 Output nets */
wire t_6963,   t_6964,   t_6965;
/* u2_2396 Output nets */
wire t_6966,   t_6967,   t_6968;
/* u2_2397 Output nets */
wire t_6969,   t_6970,   t_6971;
/* u2_2398 Output nets */
wire t_6972,   t_6973,   t_6974;
/* u1_2399 Output nets */
wire t_6975,   t_6976;
/* u2_2400 Output nets */
wire t_6977,   t_6978,   t_6979;
/* u2_2401 Output nets */
wire t_6980,   t_6981,   t_6982;
/* u2_2402 Output nets */
wire t_6983,   t_6984,   t_6985;
/* u2_2403 Output nets */
wire t_6986,   t_6987,   t_6988;
/* u1_2404 Output nets */
wire t_6989,   t_6990;
/* u2_2405 Output nets */
wire t_6991,   t_6992,   t_6993;
/* u2_2406 Output nets */
wire t_6994,   t_6995,   t_6996;
/* u2_2407 Output nets */
wire t_6997,   t_6998,   t_6999;
/* u2_2408 Output nets */
wire t_7000,   t_7001,   t_7002;
/* u2_2409 Output nets */
wire t_7003,   t_7004,   t_7005;
/* u2_2410 Output nets */
wire t_7006,   t_7007,   t_7008;
/* u2_2411 Output nets */
wire t_7009,   t_7010,   t_7011;
/* u2_2412 Output nets */
wire t_7012,   t_7013,   t_7014;
/* u2_2413 Output nets */
wire t_7015,   t_7016,   t_7017;
/* u1_2414 Output nets */
wire t_7018,   t_7019;
/* u2_2415 Output nets */
wire t_7020,   t_7021,   t_7022;
/* u2_2416 Output nets */
wire t_7023,   t_7024,   t_7025;
/* u2_2417 Output nets */
wire t_7026,   t_7027,   t_7028;
/* u2_2418 Output nets */
wire t_7029,   t_7030,   t_7031;
/* u1_2419 Output nets */
wire t_7032,   t_7033;
/* u2_2420 Output nets */
wire t_7034,   t_7035,   t_7036;
/* u2_2421 Output nets */
wire t_7037,   t_7038,   t_7039;
/* u2_2422 Output nets */
wire t_7040,   t_7041,   t_7042;
/* u2_2423 Output nets */
wire t_7043,   t_7044,   t_7045;
/* u2_2424 Output nets */
wire t_7046,   t_7047,   t_7048;
/* u2_2425 Output nets */
wire t_7049,   t_7050,   t_7051;
/* u2_2426 Output nets */
wire t_7052,   t_7053,   t_7054;
/* u2_2427 Output nets */
wire t_7055,   t_7056,   t_7057;
/* u2_2428 Output nets */
wire t_7058,   t_7059,   t_7060;
/* u2_2429 Output nets */
wire t_7061,   t_7062,   t_7063;
/* u2_2430 Output nets */
wire t_7064,   t_7065,   t_7066;
/* u2_2431 Output nets */
wire t_7067,   t_7068,   t_7069;
/* u2_2432 Output nets */
wire t_7070,   t_7071,   t_7072;
/* u2_2433 Output nets */
wire t_7073,   t_7074,   t_7075;
/* u2_2434 Output nets */
wire t_7076,   t_7077,   t_7078;
/* u2_2435 Output nets */
wire t_7079,   t_7080,   t_7081;
/* u2_2436 Output nets */
wire t_7082,   t_7083,   t_7084;
/* u2_2437 Output nets */
wire t_7085,   t_7086,   t_7087;
/* u2_2438 Output nets */
wire t_7088,   t_7089,   t_7090;
/* u2_2439 Output nets */
wire t_7091,   t_7092,   t_7093;
/* u2_2440 Output nets */
wire t_7094,   t_7095,   t_7096;
/* u2_2441 Output nets */
wire t_7097,   t_7098,   t_7099;
/* u2_2442 Output nets */
wire t_7100,   t_7101,   t_7102;
/* u2_2443 Output nets */
wire t_7103,   t_7104,   t_7105;
/* u2_2444 Output nets */
wire t_7106,   t_7107,   t_7108;
/* u2_2445 Output nets */
wire t_7109,   t_7110,   t_7111;
/* u2_2446 Output nets */
wire t_7112,   t_7113,   t_7114;
/* u2_2447 Output nets */
wire t_7115,   t_7116,   t_7117;
/* u2_2448 Output nets */
wire t_7118,   t_7119,   t_7120;
/* u2_2449 Output nets */
wire t_7121,   t_7122,   t_7123;
/* u0_2450 Output nets */
wire t_7124,   t_7125;
/* u2_2451 Output nets */
wire t_7126,   t_7127,   t_7128;
/* u2_2452 Output nets */
wire t_7129,   t_7130,   t_7131;
/* u2_2453 Output nets */
wire t_7132,   t_7133,   t_7134;
/* u2_2454 Output nets */
wire t_7135,   t_7136,   t_7137;
/* u2_2455 Output nets */
wire t_7138,   t_7139,   t_7140;
/* u0_2456 Output nets */
wire t_7141,   t_7142;
/* u2_2457 Output nets */
wire t_7143,   t_7144,   t_7145;
/* u2_2458 Output nets */
wire t_7146,   t_7147,   t_7148;
/* u2_2459 Output nets */
wire t_7149,   t_7150,   t_7151;
/* u2_2460 Output nets */
wire t_7152,   t_7153,   t_7154;
/* u2_2461 Output nets */
wire t_7155,   t_7156,   t_7157;
/* u0_2462 Output nets */
wire t_7158,   t_7159;
/* u2_2463 Output nets */
wire t_7160,   t_7161,   t_7162;
/* u2_2464 Output nets */
wire t_7163,   t_7164,   t_7165;
/* u2_2465 Output nets */
wire t_7166,   t_7167,   t_7168;
/* u2_2466 Output nets */
wire t_7169,   t_7170,   t_7171;
/* u2_2467 Output nets */
wire t_7172,   t_7173,   t_7174;
/* u1_2468 Output nets */
wire t_7175,   t_7176;
/* u2_2469 Output nets */
wire t_7177,   t_7178,   t_7179;
/* u2_2470 Output nets */
wire t_7180,   t_7181,   t_7182;
/* u2_2471 Output nets */
wire t_7183,   t_7184,   t_7185;
/* u2_2472 Output nets */
wire t_7186,   t_7187,   t_7188;
/* u2_2473 Output nets */
wire t_7189,   t_7190,   t_7191;
/* u1_2474 Output nets */
wire t_7192,   t_7193;
/* u2_2475 Output nets */
wire t_7194,   t_7195,   t_7196;
/* u2_2476 Output nets */
wire t_7197,   t_7198,   t_7199;
/* u2_2477 Output nets */
wire t_7200,   t_7201,   t_7202;
/* u2_2478 Output nets */
wire t_7203,   t_7204,   t_7205;
/* u2_2479 Output nets */
wire t_7206,   t_7207,   t_7208;
/* u1_2480 Output nets */
wire t_7209,   t_7210;
/* u2_2481 Output nets */
wire t_7211,   t_7212,   t_7213;
/* u2_2482 Output nets */
wire t_7214,   t_7215,   t_7216;
/* u2_2483 Output nets */
wire t_7217,   t_7218,   t_7219;
/* u2_2484 Output nets */
wire t_7220,   t_7221,   t_7222;
/* u2_2485 Output nets */
wire t_7223,   t_7224,   t_7225;
/* u1_2486 Output nets */
wire t_7226,   t_7227;
/* u2_2487 Output nets */
wire t_7228,   t_7229,   t_7230;
/* u2_2488 Output nets */
wire t_7231,   t_7232,   t_7233;
/* u2_2489 Output nets */
wire t_7234,   t_7235,   t_7236;
/* u2_2490 Output nets */
wire t_7237,   t_7238,   t_7239;
/* u2_2491 Output nets */
wire t_7240,   t_7241,   t_7242;
/* u1_2492 Output nets */
wire t_7243,   t_7244;
/* u2_2493 Output nets */
wire t_7245,   t_7246,   t_7247;
/* u2_2494 Output nets */
wire t_7248,   t_7249,   t_7250;
/* u2_2495 Output nets */
wire t_7251,   t_7252,   t_7253;
/* u2_2496 Output nets */
wire t_7254,   t_7255,   t_7256;
/* u2_2497 Output nets */
wire t_7257,   t_7258,   t_7259;
/* u2_2498 Output nets */
wire t_7260,   t_7261,   t_7262;
/* u2_2499 Output nets */
wire t_7263,   t_7264,   t_7265;
/* u2_2500 Output nets */
wire t_7266,   t_7267,   t_7268;
/* u2_2501 Output nets */
wire t_7269,   t_7270,   t_7271;
/* u2_2502 Output nets */
wire t_7272,   t_7273,   t_7274;
/* u2_2503 Output nets */
wire t_7275,   t_7276,   t_7277;
/* u1_2504 Output nets */
wire t_7278,   t_7279;
/* u2_2505 Output nets */
wire t_7280,   t_7281,   t_7282;
/* u2_2506 Output nets */
wire t_7283,   t_7284,   t_7285;
/* u2_2507 Output nets */
wire t_7286,   t_7287,   t_7288;
/* u2_2508 Output nets */
wire t_7289,   t_7290,   t_7291;
/* u2_2509 Output nets */
wire t_7292,   t_7293,   t_7294;
/* u1_2510 Output nets */
wire t_7295,   t_7296;
/* u2_2511 Output nets */
wire t_7297,   t_7298,   t_7299;
/* u2_2512 Output nets */
wire t_7300,   t_7301,   t_7302;
/* u2_2513 Output nets */
wire t_7303,   t_7304,   t_7305;
/* u2_2514 Output nets */
wire t_7306,   t_7307,   t_7308;
/* u2_2515 Output nets */
wire t_7309,   t_7310,   t_7311;
/* u2_2516 Output nets */
wire t_7312,   t_7313,   t_7314;
/* u2_2517 Output nets */
wire t_7315,   t_7316,   t_7317;
/* u2_2518 Output nets */
wire t_7318,   t_7319,   t_7320;
/* u2_2519 Output nets */
wire t_7321,   t_7322,   t_7323;
/* u2_2520 Output nets */
wire t_7324,   t_7325,   t_7326;
/* u2_2521 Output nets */
wire t_7327,   t_7328,   t_7329;
/* u2_2522 Output nets */
wire t_7330,   t_7331,   t_7332;
/* u2_2523 Output nets */
wire t_7333,   t_7334,   t_7335;
/* u2_2524 Output nets */
wire t_7336,   t_7337,   t_7338;
/* u2_2525 Output nets */
wire t_7339,   t_7340,   t_7341;
/* u2_2526 Output nets */
wire t_7342,   t_7343,   t_7344;
/* u2_2527 Output nets */
wire t_7345,   t_7346,   t_7347;
/* u2_2528 Output nets */
wire t_7348,   t_7349,   t_7350;
/* u2_2529 Output nets */
wire t_7351,   t_7352,   t_7353;
/* u2_2530 Output nets */
wire t_7354,   t_7355,   t_7356;
/* u2_2531 Output nets */
wire t_7357,   t_7358,   t_7359;
/* u2_2532 Output nets */
wire t_7360,   t_7361,   t_7362;
/* u2_2533 Output nets */
wire t_7363,   t_7364,   t_7365;
/* u2_2534 Output nets */
wire t_7366,   t_7367,   t_7368;
/* u2_2535 Output nets */
wire t_7369,   t_7370,   t_7371;
/* u2_2536 Output nets */
wire t_7372,   t_7373,   t_7374;
/* u2_2537 Output nets */
wire t_7375,   t_7376,   t_7377;
/* u2_2538 Output nets */
wire t_7378,   t_7379,   t_7380;
/* u2_2539 Output nets */
wire t_7381,   t_7382,   t_7383;
/* u2_2540 Output nets */
wire t_7384,   t_7385,   t_7386;
/* u2_2541 Output nets */
wire t_7387,   t_7388,   t_7389;
/* u2_2542 Output nets */
wire t_7390,   t_7391,   t_7392;
/* u2_2543 Output nets */
wire t_7393,   t_7394,   t_7395;
/* u2_2544 Output nets */
wire t_7396,   t_7397,   t_7398;
/* u2_2545 Output nets */
wire t_7399,   t_7400,   t_7401;
/* u2_2546 Output nets */
wire t_7402,   t_7403,   t_7404;
/* u0_2547 Output nets */
wire t_7405,   t_7406;
/* u2_2548 Output nets */
wire t_7407,   t_7408,   t_7409;
/* u2_2549 Output nets */
wire t_7410,   t_7411,   t_7412;
/* u2_2550 Output nets */
wire t_7413,   t_7414,   t_7415;
/* u2_2551 Output nets */
wire t_7416,   t_7417,   t_7418;
/* u2_2552 Output nets */
wire t_7419,   t_7420,   t_7421;
/* u2_2553 Output nets */
wire t_7422,   t_7423,   t_7424;
/* u0_2554 Output nets */
wire t_7425,   t_7426;
/* u2_2555 Output nets */
wire t_7427,   t_7428,   t_7429;
/* u2_2556 Output nets */
wire t_7430,   t_7431,   t_7432;
/* u2_2557 Output nets */
wire t_7433,   t_7434,   t_7435;
/* u2_2558 Output nets */
wire t_7436,   t_7437,   t_7438;
/* u2_2559 Output nets */
wire t_7439,   t_7440,   t_7441;
/* u2_2560 Output nets */
wire t_7442,   t_7443,   t_7444;
/* u0_2561 Output nets */
wire t_7445,   t_7446;
/* u2_2562 Output nets */
wire t_7447,   t_7448,   t_7449;
/* u2_2563 Output nets */
wire t_7450,   t_7451,   t_7452;
/* u2_2564 Output nets */
wire t_7453,   t_7454,   t_7455;
/* u2_2565 Output nets */
wire t_7456,   t_7457,   t_7458;
/* u2_2566 Output nets */
wire t_7459,   t_7460,   t_7461;
/* u2_2567 Output nets */
wire t_7462,   t_7463,   t_7464;
/* u1_2568 Output nets */
wire t_7465,   t_7466;
/* u2_2569 Output nets */
wire t_7467,   t_7468,   t_7469;
/* u2_2570 Output nets */
wire t_7470,   t_7471,   t_7472;
/* u2_2571 Output nets */
wire t_7473,   t_7474,   t_7475;
/* u2_2572 Output nets */
wire t_7476,   t_7477,   t_7478;
/* u2_2573 Output nets */
wire t_7479,   t_7480,   t_7481;
/* u2_2574 Output nets */
wire t_7482,   t_7483,   t_7484;
/* u1_2575 Output nets */
wire t_7485,   t_7486;
/* u2_2576 Output nets */
wire t_7487,   t_7488,   t_7489;
/* u2_2577 Output nets */
wire t_7490,   t_7491,   t_7492;
/* u2_2578 Output nets */
wire t_7493,   t_7494,   t_7495;
/* u2_2579 Output nets */
wire t_7496,   t_7497,   t_7498;
/* u2_2580 Output nets */
wire t_7499,   t_7500,   t_7501;
/* u2_2581 Output nets */
wire t_7502,   t_7503,   t_7504;
/* u1_2582 Output nets */
wire t_7505,   t_7506;
/* u2_2583 Output nets */
wire t_7507,   t_7508,   t_7509;
/* u2_2584 Output nets */
wire t_7510,   t_7511,   t_7512;
/* u2_2585 Output nets */
wire t_7513,   t_7514,   t_7515;
/* u2_2586 Output nets */
wire t_7516,   t_7517,   t_7518;
/* u2_2587 Output nets */
wire t_7519,   t_7520,   t_7521;
/* u2_2588 Output nets */
wire t_7522,   t_7523,   t_7524;
/* u1_2589 Output nets */
wire t_7525,   t_7526;
/* u2_2590 Output nets */
wire t_7527,   t_7528,   t_7529;
/* u2_2591 Output nets */
wire t_7530,   t_7531,   t_7532;
/* u2_2592 Output nets */
wire t_7533,   t_7534,   t_7535;
/* u2_2593 Output nets */
wire t_7536,   t_7537,   t_7538;
/* u2_2594 Output nets */
wire t_7539,   t_7540,   t_7541;
/* u2_2595 Output nets */
wire t_7542,   t_7543,   t_7544;
/* u1_2596 Output nets */
wire t_7545,   t_7546;
/* u2_2597 Output nets */
wire t_7547,   t_7548,   t_7549;
/* u2_2598 Output nets */
wire t_7550,   t_7551,   t_7552;
/* u2_2599 Output nets */
wire t_7553,   t_7554,   t_7555;
/* u2_2600 Output nets */
wire t_7556,   t_7557,   t_7558;
/* u2_2601 Output nets */
wire t_7559,   t_7560,   t_7561;
/* u2_2602 Output nets */
wire t_7562,   t_7563,   t_7564;
/* u2_2603 Output nets */
wire t_7565,   t_7566,   t_7567;
/* u2_2604 Output nets */
wire t_7568,   t_7569,   t_7570;
/* u2_2605 Output nets */
wire t_7571,   t_7572,   t_7573;
/* u2_2606 Output nets */
wire t_7574,   t_7575,   t_7576;
/* u2_2607 Output nets */
wire t_7577,   t_7578,   t_7579;
/* u2_2608 Output nets */
wire t_7580,   t_7581,   t_7582;
/* u2_2609 Output nets */
wire t_7583,   t_7584,   t_7585;
/* u1_2610 Output nets */
wire t_7586,   t_7587;
/* u2_2611 Output nets */
wire t_7588,   t_7589,   t_7590;
/* u2_2612 Output nets */
wire t_7591,   t_7592,   t_7593;
/* u2_2613 Output nets */
wire t_7594,   t_7595,   t_7596;
/* u2_2614 Output nets */
wire t_7597,   t_7598,   t_7599;
/* u2_2615 Output nets */
wire t_7600,   t_7601,   t_7602;
/* u2_2616 Output nets */
wire t_7603,   t_7604,   t_7605;
/* u1_2617 Output nets */
wire t_7606,   t_7607;
/* u2_2618 Output nets */
wire t_7608,   t_7609,   t_7610;
/* u2_2619 Output nets */
wire t_7611,   t_7612,   t_7613;
/* u2_2620 Output nets */
wire t_7614,   t_7615,   t_7616;
/* u2_2621 Output nets */
wire t_7617,   t_7618,   t_7619;
/* u2_2622 Output nets */
wire t_7620,   t_7621,   t_7622;
/* u2_2623 Output nets */
wire t_7623,   t_7624,   t_7625;
/* u2_2624 Output nets */
wire t_7626,   t_7627,   t_7628;
/* u2_2625 Output nets */
wire t_7629,   t_7630,   t_7631;
/* u2_2626 Output nets */
wire t_7632,   t_7633,   t_7634;
/* u2_2627 Output nets */
wire t_7635,   t_7636,   t_7637;
/* u2_2628 Output nets */
wire t_7638,   t_7639,   t_7640;
/* u2_2629 Output nets */
wire t_7641,   t_7642,   t_7643;
/* u2_2630 Output nets */
wire t_7644,   t_7645,   t_7646;
/* u2_2631 Output nets */
wire t_7647,   t_7648,   t_7649;
/* u2_2632 Output nets */
wire t_7650,   t_7651,   t_7652;
/* u2_2633 Output nets */
wire t_7653,   t_7654,   t_7655;
/* u2_2634 Output nets */
wire t_7656,   t_7657,   t_7658;
/* u2_2635 Output nets */
wire t_7659,   t_7660,   t_7661;
/* u2_2636 Output nets */
wire t_7662,   t_7663,   t_7664;
/* u2_2637 Output nets */
wire t_7665,   t_7666,   t_7667;
/* u2_2638 Output nets */
wire t_7668,   t_7669,   t_7670;
/* u2_2639 Output nets */
wire t_7671,   t_7672,   t_7673;
/* u2_2640 Output nets */
wire t_7674,   t_7675,   t_7676;
/* u2_2641 Output nets */
wire t_7677,   t_7678,   t_7679;
/* u2_2642 Output nets */
wire t_7680,   t_7681,   t_7682;
/* u2_2643 Output nets */
wire t_7683,   t_7684,   t_7685;
/* u2_2644 Output nets */
wire t_7686,   t_7687,   t_7688;
/* u2_2645 Output nets */
wire t_7689,   t_7690,   t_7691;
/* u2_2646 Output nets */
wire t_7692,   t_7693,   t_7694;
/* u2_2647 Output nets */
wire t_7695,   t_7696,   t_7697;
/* u2_2648 Output nets */
wire t_7698,   t_7699,   t_7700;
/* u2_2649 Output nets */
wire t_7701,   t_7702,   t_7703;
/* u2_2650 Output nets */
wire t_7704,   t_7705,   t_7706;
/* u2_2651 Output nets */
wire t_7707,   t_7708,   t_7709;
/* u2_2652 Output nets */
wire t_7710,   t_7711,   t_7712;
/* u2_2653 Output nets */
wire t_7713,   t_7714,   t_7715;
/* u2_2654 Output nets */
wire t_7716,   t_7717,   t_7718;
/* u2_2655 Output nets */
wire t_7719,   t_7720,   t_7721;
/* u2_2656 Output nets */
wire t_7722,   t_7723,   t_7724;
/* u2_2657 Output nets */
wire t_7725,   t_7726,   t_7727;
/* u2_2658 Output nets */
wire t_7728,   t_7729,   t_7730;
/* u2_2659 Output nets */
wire t_7731,   t_7732,   t_7733;
/* u0_2660 Output nets */
wire t_7734,   t_7735;
/* u2_2661 Output nets */
wire t_7736,   t_7737,   t_7738;
/* u2_2662 Output nets */
wire t_7739,   t_7740,   t_7741;
/* u2_2663 Output nets */
wire t_7742,   t_7743,   t_7744;
/* u2_2664 Output nets */
wire t_7745,   t_7746,   t_7747;
/* u2_2665 Output nets */
wire t_7748,   t_7749,   t_7750;
/* u2_2666 Output nets */
wire t_7751,   t_7752,   t_7753;
/* u2_2667 Output nets */
wire t_7754,   t_7755,   t_7756;
/* u0_2668 Output nets */
wire t_7757,   t_7758;
/* u2_2669 Output nets */
wire t_7759,   t_7760,   t_7761;
/* u2_2670 Output nets */
wire t_7762,   t_7763,   t_7764;
/* u2_2671 Output nets */
wire t_7765,   t_7766,   t_7767;
/* u2_2672 Output nets */
wire t_7768,   t_7769,   t_7770;
/* u2_2673 Output nets */
wire t_7771,   t_7772,   t_7773;
/* u2_2674 Output nets */
wire t_7774,   t_7775,   t_7776;
/* u2_2675 Output nets */
wire t_7777,   t_7778,   t_7779;
/* u0_2676 Output nets */
wire t_7780,   t_7781;
/* u2_2677 Output nets */
wire t_7782,   t_7783,   t_7784;
/* u2_2678 Output nets */
wire t_7785,   t_7786,   t_7787;
/* u2_2679 Output nets */
wire t_7788,   t_7789,   t_7790;
/* u2_2680 Output nets */
wire t_7791,   t_7792,   t_7793;
/* u2_2681 Output nets */
wire t_7794,   t_7795,   t_7796;
/* u2_2682 Output nets */
wire t_7797,   t_7798,   t_7799;
/* u2_2683 Output nets */
wire t_7800,   t_7801,   t_7802;
/* u1_2684 Output nets */
wire t_7803,   t_7804;
/* u2_2685 Output nets */
wire t_7805,   t_7806,   t_7807;
/* u2_2686 Output nets */
wire t_7808,   t_7809,   t_7810;
/* u2_2687 Output nets */
wire t_7811,   t_7812,   t_7813;
/* u2_2688 Output nets */
wire t_7814,   t_7815,   t_7816;
/* u2_2689 Output nets */
wire t_7817,   t_7818,   t_7819;
/* u2_2690 Output nets */
wire t_7820,   t_7821,   t_7822;
/* u2_2691 Output nets */
wire t_7823,   t_7824,   t_7825;
/* u1_2692 Output nets */
wire t_7826,   t_7827;
/* u2_2693 Output nets */
wire t_7828,   t_7829,   t_7830;
/* u2_2694 Output nets */
wire t_7831,   t_7832,   t_7833;
/* u2_2695 Output nets */
wire t_7834,   t_7835,   t_7836;
/* u2_2696 Output nets */
wire t_7837,   t_7838,   t_7839;
/* u2_2697 Output nets */
wire t_7840,   t_7841,   t_7842;
/* u2_2698 Output nets */
wire t_7843,   t_7844,   t_7845;
/* u2_2699 Output nets */
wire t_7846,   t_7847,   t_7848;
/* u1_2700 Output nets */
wire t_7849,   t_7850;
/* u2_2701 Output nets */
wire t_7851,   t_7852,   t_7853;
/* u2_2702 Output nets */
wire t_7854,   t_7855,   t_7856;
/* u2_2703 Output nets */
wire t_7857,   t_7858,   t_7859;
/* u2_2704 Output nets */
wire t_7860,   t_7861,   t_7862;
/* u2_2705 Output nets */
wire t_7863,   t_7864,   t_7865;
/* u2_2706 Output nets */
wire t_7866,   t_7867,   t_7868;
/* u2_2707 Output nets */
wire t_7869,   t_7870,   t_7871;
/* u1_2708 Output nets */
wire t_7872,   t_7873;
/* u2_2709 Output nets */
wire t_7874,   t_7875,   t_7876;
/* u2_2710 Output nets */
wire t_7877,   t_7878,   t_7879;
/* u2_2711 Output nets */
wire t_7880,   t_7881,   t_7882;
/* u2_2712 Output nets */
wire t_7883,   t_7884,   t_7885;
/* u2_2713 Output nets */
wire t_7886,   t_7887,   t_7888;
/* u2_2714 Output nets */
wire t_7889,   t_7890,   t_7891;
/* u2_2715 Output nets */
wire t_7892,   t_7893,   t_7894;
/* u1_2716 Output nets */
wire t_7895,   t_7896;
/* u2_2717 Output nets */
wire t_7897,   t_7898,   t_7899;
/* u2_2718 Output nets */
wire t_7900,   t_7901,   t_7902;
/* u2_2719 Output nets */
wire t_7903,   t_7904,   t_7905;
/* u2_2720 Output nets */
wire t_7906,   t_7907,   t_7908;
/* u2_2721 Output nets */
wire t_7909,   t_7910,   t_7911;
/* u2_2722 Output nets */
wire t_7912,   t_7913,   t_7914;
/* u2_2723 Output nets */
wire t_7915,   t_7916,   t_7917;
/* u2_2724 Output nets */
wire t_7918,   t_7919,   t_7920;
/* u2_2725 Output nets */
wire t_7921,   t_7922,   t_7923;
/* u2_2726 Output nets */
wire t_7924,   t_7925,   t_7926;
/* u2_2727 Output nets */
wire t_7927,   t_7928,   t_7929;
/* u2_2728 Output nets */
wire t_7930,   t_7931,   t_7932;
/* u2_2729 Output nets */
wire t_7933,   t_7934,   t_7935;
/* u2_2730 Output nets */
wire t_7936,   t_7937,   t_7938;
/* u2_2731 Output nets */
wire t_7939,   t_7940,   t_7941;
/* u1_2732 Output nets */
wire t_7942,   t_7943;
/* u2_2733 Output nets */
wire t_7944,   t_7945,   t_7946;
/* u2_2734 Output nets */
wire t_7947,   t_7948,   t_7949;
/* u2_2735 Output nets */
wire t_7950,   t_7951,   t_7952;
/* u2_2736 Output nets */
wire t_7953,   t_7954,   t_7955;
/* u2_2737 Output nets */
wire t_7956,   t_7957,   t_7958;
/* u2_2738 Output nets */
wire t_7959,   t_7960,   t_7961;
/* u2_2739 Output nets */
wire t_7962,   t_7963,   t_7964;
/* u1_2740 Output nets */
wire t_7965,   t_7966;
/* u2_2741 Output nets */
wire t_7967,   t_7968,   t_7969;
/* u2_2742 Output nets */
wire t_7970,   t_7971,   t_7972;
/* u2_2743 Output nets */
wire t_7973,   t_7974,   t_7975;
/* u2_2744 Output nets */
wire t_7976,   t_7977,   t_7978;
/* u2_2745 Output nets */
wire t_7979,   t_7980,   t_7981;
/* u2_2746 Output nets */
wire t_7982,   t_7983,   t_7984;
/* u2_2747 Output nets */
wire t_7985,   t_7986,   t_7987;
/* u2_2748 Output nets */
wire t_7988,   t_7989,   t_7990;
/* u2_2749 Output nets */
wire t_7991,   t_7992,   t_7993;
/* u2_2750 Output nets */
wire t_7994,   t_7995,   t_7996;
/* u2_2751 Output nets */
wire t_7997,   t_7998,   t_7999;
/* u2_2752 Output nets */
wire t_8000,   t_8001,   t_8002;
/* u2_2753 Output nets */
wire t_8003,   t_8004,   t_8005;
/* u2_2754 Output nets */
wire t_8006,   t_8007,   t_8008;
/* u2_2755 Output nets */
wire t_8009,   t_8010,   t_8011;
/* u2_2756 Output nets */
wire t_8012,   t_8013,   t_8014;
/* u2_2757 Output nets */
wire t_8015,   t_8016,   t_8017;
/* u2_2758 Output nets */
wire t_8018,   t_8019,   t_8020;
/* u2_2759 Output nets */
wire t_8021,   t_8022,   t_8023;
/* u2_2760 Output nets */
wire t_8024,   t_8025,   t_8026;
/* u2_2761 Output nets */
wire t_8027,   t_8028,   t_8029;
/* u2_2762 Output nets */
wire t_8030,   t_8031,   t_8032;
/* u2_2763 Output nets */
wire t_8033,   t_8034,   t_8035;
/* u2_2764 Output nets */
wire t_8036,   t_8037,   t_8038;
/* u2_2765 Output nets */
wire t_8039,   t_8040,   t_8041;
/* u2_2766 Output nets */
wire t_8042,   t_8043,   t_8044;
/* u2_2767 Output nets */
wire t_8045,   t_8046,   t_8047;
/* u2_2768 Output nets */
wire t_8048,   t_8049,   t_8050;
/* u2_2769 Output nets */
wire t_8051,   t_8052,   t_8053;
/* u2_2770 Output nets */
wire t_8054,   t_8055,   t_8056;
/* u2_2771 Output nets */
wire t_8057,   t_8058,   t_8059;
/* u2_2772 Output nets */
wire t_8060,   t_8061,   t_8062;
/* u2_2773 Output nets */
wire t_8063,   t_8064,   t_8065;
/* u2_2774 Output nets */
wire t_8066,   t_8067,   t_8068;
/* u2_2775 Output nets */
wire t_8069,   t_8070,   t_8071;
/* u2_2776 Output nets */
wire t_8072,   t_8073,   t_8074;
/* u2_2777 Output nets */
wire t_8075,   t_8076,   t_8077;
/* u2_2778 Output nets */
wire t_8078,   t_8079,   t_8080;
/* u2_2779 Output nets */
wire t_8081,   t_8082,   t_8083;
/* u2_2780 Output nets */
wire t_8084,   t_8085,   t_8086;
/* u2_2781 Output nets */
wire t_8087,   t_8088,   t_8089;
/* u2_2782 Output nets */
wire t_8090,   t_8091,   t_8092;
/* u2_2783 Output nets */
wire t_8093,   t_8094,   t_8095;
/* u2_2784 Output nets */
wire t_8096,   t_8097,   t_8098;
/* u2_2785 Output nets */
wire t_8099,   t_8100,   t_8101;
/* u2_2786 Output nets */
wire t_8102,   t_8103,   t_8104;
/* u2_2787 Output nets */
wire t_8105,   t_8106,   t_8107;
/* u2_2788 Output nets */
wire t_8108,   t_8109,   t_8110;
/* u2_2789 Output nets */
wire t_8111,   t_8112,   t_8113;
/* u2_2790 Output nets */
wire t_8114,   t_8115,   t_8116;
/* u2_2791 Output nets */
wire t_8117,   t_8118,   t_8119;
/* u2_2792 Output nets */
wire t_8120,   t_8121,   t_8122;
/* u2_2793 Output nets */
wire t_8123,   t_8124,   t_8125;
/* u2_2794 Output nets */
wire t_8126,   t_8127,   t_8128;
/* u2_2795 Output nets */
wire t_8129,   t_8130,   t_8131;
/* u2_2796 Output nets */
wire t_8132,   t_8133,   t_8134;
/* u2_2797 Output nets */
wire t_8135,   t_8136,   t_8137;
/* u2_2798 Output nets */
wire t_8138,   t_8139,   t_8140;
/* u2_2799 Output nets */
wire t_8141,   t_8142,   t_8143;
/* u2_2800 Output nets */
wire t_8144,   t_8145,   t_8146;
/* u2_2801 Output nets */
wire t_8147,   t_8148,   t_8149;
/* u2_2802 Output nets */
wire t_8150,   t_8151,   t_8152;
/* u2_2803 Output nets */
wire t_8153,   t_8154,   t_8155;
/* u2_2804 Output nets */
wire t_8156,   t_8157,   t_8158;
/* u2_2805 Output nets */
wire t_8159,   t_8160,   t_8161;
/* u2_2806 Output nets */
wire t_8162,   t_8163,   t_8164;
/* u2_2807 Output nets */
wire t_8165,   t_8166,   t_8167;
/* u2_2808 Output nets */
wire t_8168,   t_8169,   t_8170;
/* u2_2809 Output nets */
wire t_8171,   t_8172,   t_8173;
/* u2_2810 Output nets */
wire t_8174,   t_8175,   t_8176;
/* u2_2811 Output nets */
wire t_8177,   t_8178,   t_8179;
/* u2_2812 Output nets */
wire t_8180,   t_8181,   t_8182;
/* u2_2813 Output nets */
wire t_8183,   t_8184,   t_8185;
/* u2_2814 Output nets */
wire t_8186,   t_8187,   t_8188;
/* u2_2815 Output nets */
wire t_8189,   t_8190,   t_8191;
/* u2_2816 Output nets */
wire t_8192,   t_8193,   t_8194;
/* u2_2817 Output nets */
wire t_8195,   t_8196,   t_8197;
/* u2_2818 Output nets */
wire t_8198,   t_8199,   t_8200;
/* u2_2819 Output nets */
wire t_8201,   t_8202,   t_8203;
/* u1_2820 Output nets */
wire t_8204,   t_8205;
/* u2_2821 Output nets */
wire t_8206,   t_8207,   t_8208;
/* u2_2822 Output nets */
wire t_8209,   t_8210,   t_8211;
/* u2_2823 Output nets */
wire t_8212,   t_8213,   t_8214;
/* u2_2824 Output nets */
wire t_8215,   t_8216,   t_8217;
/* u2_2825 Output nets */
wire t_8218,   t_8219,   t_8220;
/* u2_2826 Output nets */
wire t_8221,   t_8222,   t_8223;
/* u2_2827 Output nets */
wire t_8224,   t_8225,   t_8226;
/* u1_2828 Output nets */
wire t_8227,   t_8228;
/* u2_2829 Output nets */
wire t_8229,   t_8230,   t_8231;
/* u2_2830 Output nets */
wire t_8232,   t_8233,   t_8234;
/* u2_2831 Output nets */
wire t_8235,   t_8236,   t_8237;
/* u2_2832 Output nets */
wire t_8238,   t_8239,   t_8240;
/* u2_2833 Output nets */
wire t_8241,   t_8242,   t_8243;
/* u2_2834 Output nets */
wire t_8244,   t_8245,   t_8246;
/* u2_2835 Output nets */
wire t_8247,   t_8248,   t_8249;
/* u1_2836 Output nets */
wire t_8250,   t_8251;
/* u2_2837 Output nets */
wire t_8252,   t_8253,   t_8254;
/* u2_2838 Output nets */
wire t_8255,   t_8256,   t_8257;
/* u2_2839 Output nets */
wire t_8258,   t_8259,   t_8260;
/* u2_2840 Output nets */
wire t_8261,   t_8262,   t_8263;
/* u2_2841 Output nets */
wire t_8264,   t_8265,   t_8266;
/* u2_2842 Output nets */
wire t_8267,   t_8268,   t_8269;
/* u2_2843 Output nets */
wire t_8270,   t_8271,   t_8272;
/* u1_2844 Output nets */
wire t_8273,   t_8274;
/* u2_2845 Output nets */
wire t_8275,   t_8276,   t_8277;
/* u2_2846 Output nets */
wire t_8278,   t_8279,   t_8280;
/* u2_2847 Output nets */
wire t_8281,   t_8282,   t_8283;
/* u2_2848 Output nets */
wire t_8284,   t_8285,   t_8286;
/* u2_2849 Output nets */
wire t_8287,   t_8288,   t_8289;
/* u2_2850 Output nets */
wire t_8290,   t_8291,   t_8292;
/* u2_2851 Output nets */
wire t_8293,   t_8294,   t_8295;
/* u1_2852 Output nets */
wire t_8296,   t_8297;
/* u2_2853 Output nets */
wire t_8298,   t_8299,   t_8300;
/* u2_2854 Output nets */
wire t_8301,   t_8302,   t_8303;
/* u2_2855 Output nets */
wire t_8304,   t_8305,   t_8306;
/* u2_2856 Output nets */
wire t_8307,   t_8308,   t_8309;
/* u2_2857 Output nets */
wire t_8310,   t_8311,   t_8312;
/* u2_2858 Output nets */
wire t_8313,   t_8314,   t_8315;
/* u2_2859 Output nets */
wire t_8316,   t_8317,   t_8318;
/* u1_2860 Output nets */
wire t_8319,   t_8320;
/* u2_2861 Output nets */
wire t_8321,   t_8322,   t_8323;
/* u2_2862 Output nets */
wire t_8324,   t_8325,   t_8326;
/* u2_2863 Output nets */
wire t_8327,   t_8328,   t_8329;
/* u2_2864 Output nets */
wire t_8330,   t_8331,   t_8332;
/* u2_2865 Output nets */
wire t_8333,   t_8334,   t_8335;
/* u2_2866 Output nets */
wire t_8336,   t_8337,   t_8338;
/* u2_2867 Output nets */
wire t_8339,   t_8340,   t_8341;
/* u1_2868 Output nets */
wire t_8342,   t_8343;
/* u2_2869 Output nets */
wire t_8344,   t_8345,   t_8346;
/* u2_2870 Output nets */
wire t_8347,   t_8348,   t_8349;
/* u2_2871 Output nets */
wire t_8350,   t_8351,   t_8352;
/* u2_2872 Output nets */
wire t_8353,   t_8354,   t_8355;
/* u2_2873 Output nets */
wire t_8356,   t_8357,   t_8358;
/* u2_2874 Output nets */
wire t_8359,   t_8360,   t_8361;
/* u2_2875 Output nets */
wire t_8362,   t_8363,   t_8364;
/* u1_2876 Output nets */
wire t_8365,   t_8366;
/* u2_2877 Output nets */
wire t_8367,   t_8368,   t_8369;
/* u2_2878 Output nets */
wire t_8370,   t_8371,   t_8372;
/* u2_2879 Output nets */
wire t_8373,   t_8374,   t_8375;
/* u2_2880 Output nets */
wire t_8376,   t_8377,   t_8378;
/* u2_2881 Output nets */
wire t_8379,   t_8380,   t_8381;
/* u2_2882 Output nets */
wire t_8382,   t_8383,   t_8384;
/* u2_2883 Output nets */
wire t_8385,   t_8386,   t_8387;
/* u0_2884 Output nets */
wire t_8388,   t_8389;
/* u2_2885 Output nets */
wire t_8390,   t_8391,   t_8392;
/* u2_2886 Output nets */
wire t_8393,   t_8394,   t_8395;
/* u2_2887 Output nets */
wire t_8396,   t_8397,   t_8398;
/* u2_2888 Output nets */
wire t_8399,   t_8400,   t_8401;
/* u2_2889 Output nets */
wire t_8402,   t_8403,   t_8404;
/* u2_2890 Output nets */
wire t_8405,   t_8406,   t_8407;
/* u2_2891 Output nets */
wire t_8408,   t_8409,   t_8410;
/* u0_2892 Output nets */
wire t_8411,   t_8412;
/* u2_2893 Output nets */
wire t_8413,   t_8414,   t_8415;
/* u2_2894 Output nets */
wire t_8416,   t_8417,   t_8418;
/* u2_2895 Output nets */
wire t_8419,   t_8420,   t_8421;
/* u2_2896 Output nets */
wire t_8422,   t_8423,   t_8424;
/* u2_2897 Output nets */
wire t_8425,   t_8426,   t_8427;
/* u2_2898 Output nets */
wire t_8428,   t_8429,   t_8430;
/* u2_2899 Output nets */
wire t_8431,   t_8432,   t_8433;
/* u0_2900 Output nets */
wire t_8434,   t_8435;
/* u2_2901 Output nets */
wire t_8436,   t_8437,   t_8438;
/* u2_2902 Output nets */
wire t_8439,   t_8440,   t_8441;
/* u2_2903 Output nets */
wire t_8442,   t_8443,   t_8444;
/* u2_2904 Output nets */
wire t_8445,   t_8446,   t_8447;
/* u2_2905 Output nets */
wire t_8448,   t_8449,   t_8450;
/* u2_2906 Output nets */
wire t_8451,   t_8452,   t_8453;
/* u2_2907 Output nets */
wire t_8454,   t_8455,   t_8456;
/* u0_2908 Output nets */
wire t_8457,   t_8458;
/* u2_2909 Output nets */
wire t_8459,   t_8460,   t_8461;
/* u2_2910 Output nets */
wire t_8462,   t_8463,   t_8464;
/* u2_2911 Output nets */
wire t_8465,   t_8466,   t_8467;
/* u2_2912 Output nets */
wire t_8468,   t_8469,   t_8470;
/* u2_2913 Output nets */
wire t_8471,   t_8472,   t_8473;
/* u2_2914 Output nets */
wire t_8474,   t_8475,   t_8476;
/* u2_2915 Output nets */
wire t_8477,   t_8478,   t_8479;
/* u0_2916 Output nets */
wire t_8480,   t_8481;
/* u2_2917 Output nets */
wire t_8482,   t_8483,   t_8484;
/* u2_2918 Output nets */
wire t_8485,   t_8486,   t_8487;
/* u2_2919 Output nets */
wire t_8488,   t_8489,   t_8490;
/* u2_2920 Output nets */
wire t_8491,   t_8492,   t_8493;
/* u2_2921 Output nets */
wire t_8494,   t_8495,   t_8496;
/* u2_2922 Output nets */
wire t_8497,   t_8498,   t_8499;
/* u2_2923 Output nets */
wire t_8500,   t_8501,   t_8502;
/* u2_2924 Output nets */
wire t_8503,   t_8504,   t_8505;
/* u2_2925 Output nets */
wire t_8506,   t_8507,   t_8508;
/* u2_2926 Output nets */
wire t_8509,   t_8510,   t_8511;
/* u2_2927 Output nets */
wire t_8512,   t_8513,   t_8514;
/* u2_2928 Output nets */
wire t_8515,   t_8516,   t_8517;
/* u2_2929 Output nets */
wire t_8518,   t_8519,   t_8520;
/* u2_2930 Output nets */
wire t_8521,   t_8522,   t_8523;
/* u2_2931 Output nets */
wire t_8524,   t_8525,   t_8526;
/* u2_2932 Output nets */
wire t_8527,   t_8528,   t_8529;
/* u2_2933 Output nets */
wire t_8530,   t_8531,   t_8532;
/* u2_2934 Output nets */
wire t_8533,   t_8534,   t_8535;
/* u2_2935 Output nets */
wire t_8536,   t_8537,   t_8538;
/* u2_2936 Output nets */
wire t_8539,   t_8540,   t_8541;
/* u2_2937 Output nets */
wire t_8542,   t_8543,   t_8544;
/* u2_2938 Output nets */
wire t_8545,   t_8546,   t_8547;
/* u2_2939 Output nets */
wire t_8548,   t_8549,   t_8550;
/* u2_2940 Output nets */
wire t_8551,   t_8552,   t_8553;
/* u2_2941 Output nets */
wire t_8554,   t_8555,   t_8556;
/* u2_2942 Output nets */
wire t_8557,   t_8558,   t_8559;
/* u2_2943 Output nets */
wire t_8560,   t_8561,   t_8562;
/* u1_2944 Output nets */
wire t_8563,   t_8564;
/* u2_2945 Output nets */
wire t_8565,   t_8566,   t_8567;
/* u2_2946 Output nets */
wire t_8568,   t_8569,   t_8570;
/* u2_2947 Output nets */
wire t_8571,   t_8572,   t_8573;
/* u2_2948 Output nets */
wire t_8574,   t_8575,   t_8576;
/* u2_2949 Output nets */
wire t_8577,   t_8578,   t_8579;
/* u2_2950 Output nets */
wire t_8580,   t_8581,   t_8582;
/* u1_2951 Output nets */
wire t_8583,   t_8584;
/* u2_2952 Output nets */
wire t_8585,   t_8586,   t_8587;
/* u2_2953 Output nets */
wire t_8588,   t_8589,   t_8590;
/* u2_2954 Output nets */
wire t_8591,   t_8592,   t_8593;
/* u2_2955 Output nets */
wire t_8594,   t_8595,   t_8596;
/* u2_2956 Output nets */
wire t_8597,   t_8598,   t_8599;
/* u2_2957 Output nets */
wire t_8600,   t_8601,   t_8602;
/* u1_2958 Output nets */
wire t_8603,   t_8604;
/* u2_2959 Output nets */
wire t_8605,   t_8606,   t_8607;
/* u2_2960 Output nets */
wire t_8608,   t_8609,   t_8610;
/* u2_2961 Output nets */
wire t_8611,   t_8612,   t_8613;
/* u2_2962 Output nets */
wire t_8614,   t_8615,   t_8616;
/* u2_2963 Output nets */
wire t_8617,   t_8618,   t_8619;
/* u2_2964 Output nets */
wire t_8620,   t_8621,   t_8622;
/* u1_2965 Output nets */
wire t_8623,   t_8624;
/* u2_2966 Output nets */
wire t_8625,   t_8626,   t_8627;
/* u2_2967 Output nets */
wire t_8628,   t_8629,   t_8630;
/* u2_2968 Output nets */
wire t_8631,   t_8632,   t_8633;
/* u2_2969 Output nets */
wire t_8634,   t_8635,   t_8636;
/* u2_2970 Output nets */
wire t_8637,   t_8638,   t_8639;
/* u2_2971 Output nets */
wire t_8640,   t_8641,   t_8642;
/* u1_2972 Output nets */
wire t_8643,   t_8644;
/* u2_2973 Output nets */
wire t_8645,   t_8646,   t_8647;
/* u2_2974 Output nets */
wire t_8648,   t_8649,   t_8650;
/* u2_2975 Output nets */
wire t_8651,   t_8652,   t_8653;
/* u2_2976 Output nets */
wire t_8654,   t_8655,   t_8656;
/* u2_2977 Output nets */
wire t_8657,   t_8658,   t_8659;
/* u2_2978 Output nets */
wire t_8660,   t_8661,   t_8662;
/* u1_2979 Output nets */
wire t_8663,   t_8664;
/* u2_2980 Output nets */
wire t_8665,   t_8666,   t_8667;
/* u2_2981 Output nets */
wire t_8668,   t_8669,   t_8670;
/* u2_2982 Output nets */
wire t_8671,   t_8672,   t_8673;
/* u2_2983 Output nets */
wire t_8674,   t_8675,   t_8676;
/* u2_2984 Output nets */
wire t_8677,   t_8678,   t_8679;
/* u2_2985 Output nets */
wire t_8680,   t_8681,   t_8682;
/* u1_2986 Output nets */
wire t_8683,   t_8684;
/* u2_2987 Output nets */
wire t_8685,   t_8686,   t_8687;
/* u2_2988 Output nets */
wire t_8688,   t_8689,   t_8690;
/* u2_2989 Output nets */
wire t_8691,   t_8692,   t_8693;
/* u2_2990 Output nets */
wire t_8694,   t_8695,   t_8696;
/* u2_2991 Output nets */
wire t_8697,   t_8698,   t_8699;
/* u2_2992 Output nets */
wire t_8700,   t_8701,   t_8702;
/* u1_2993 Output nets */
wire t_8703,   t_8704;
/* u2_2994 Output nets */
wire t_8705,   t_8706,   t_8707;
/* u2_2995 Output nets */
wire t_8708,   t_8709,   t_8710;
/* u2_2996 Output nets */
wire t_8711,   t_8712,   t_8713;
/* u2_2997 Output nets */
wire t_8714,   t_8715,   t_8716;
/* u2_2998 Output nets */
wire t_8717,   t_8718,   t_8719;
/* u2_2999 Output nets */
wire t_8720,   t_8721,   t_8722;
/* u0_3000 Output nets */
wire t_8723,   t_8724;
/* u2_3001 Output nets */
wire t_8725,   t_8726,   t_8727;
/* u2_3002 Output nets */
wire t_8728,   t_8729,   t_8730;
/* u2_3003 Output nets */
wire t_8731,   t_8732,   t_8733;
/* u2_3004 Output nets */
wire t_8734,   t_8735,   t_8736;
/* u2_3005 Output nets */
wire t_8737,   t_8738,   t_8739;
/* u2_3006 Output nets */
wire t_8740,   t_8741,   t_8742;
/* u0_3007 Output nets */
wire t_8743,   t_8744;
/* u2_3008 Output nets */
wire t_8745,   t_8746,   t_8747;
/* u2_3009 Output nets */
wire t_8748,   t_8749,   t_8750;
/* u2_3010 Output nets */
wire t_8751,   t_8752,   t_8753;
/* u2_3011 Output nets */
wire t_8754,   t_8755,   t_8756;
/* u2_3012 Output nets */
wire t_8757,   t_8758,   t_8759;
/* u2_3013 Output nets */
wire t_8760,   t_8761,   t_8762;
/* u0_3014 Output nets */
wire t_8763,   t_8764;
/* u2_3015 Output nets */
wire t_8765,   t_8766,   t_8767;
/* u2_3016 Output nets */
wire t_8768,   t_8769,   t_8770;
/* u2_3017 Output nets */
wire t_8771,   t_8772,   t_8773;
/* u2_3018 Output nets */
wire t_8774,   t_8775,   t_8776;
/* u2_3019 Output nets */
wire t_8777,   t_8778,   t_8779;
/* u2_3020 Output nets */
wire t_8780,   t_8781,   t_8782;
/* u0_3021 Output nets */
wire t_8783,   t_8784;
/* u2_3022 Output nets */
wire t_8785,   t_8786,   t_8787;
/* u2_3023 Output nets */
wire t_8788,   t_8789,   t_8790;
/* u2_3024 Output nets */
wire t_8791,   t_8792,   t_8793;
/* u2_3025 Output nets */
wire t_8794,   t_8795,   t_8796;
/* u2_3026 Output nets */
wire t_8797,   t_8798,   t_8799;
/* u2_3027 Output nets */
wire t_8800,   t_8801,   t_8802;
/* u0_3028 Output nets */
wire t_8803,   t_8804;
/* u2_3029 Output nets */
wire t_8805,   t_8806,   t_8807;
/* u2_3030 Output nets */
wire t_8808,   t_8809,   t_8810;
/* u2_3031 Output nets */
wire t_8811,   t_8812,   t_8813;
/* u2_3032 Output nets */
wire t_8814,   t_8815,   t_8816;
/* u2_3033 Output nets */
wire t_8817,   t_8818,   t_8819;
/* u2_3034 Output nets */
wire t_8820,   t_8821,   t_8822;
/* u2_3035 Output nets */
wire t_8823,   t_8824,   t_8825;
/* u2_3036 Output nets */
wire t_8826,   t_8827,   t_8828;
/* u2_3037 Output nets */
wire t_8829,   t_8830,   t_8831;
/* u2_3038 Output nets */
wire t_8832,   t_8833,   t_8834;
/* u2_3039 Output nets */
wire t_8835,   t_8836,   t_8837;
/* u2_3040 Output nets */
wire t_8838,   t_8839,   t_8840;
/* u2_3041 Output nets */
wire t_8841,   t_8842,   t_8843;
/* u2_3042 Output nets */
wire t_8844,   t_8845,   t_8846;
/* u2_3043 Output nets */
wire t_8847,   t_8848,   t_8849;
/* u2_3044 Output nets */
wire t_8850,   t_8851,   t_8852;
/* u2_3045 Output nets */
wire t_8853,   t_8854,   t_8855;
/* u2_3046 Output nets */
wire t_8856,   t_8857,   t_8858;
/* u2_3047 Output nets */
wire t_8859,   t_8860,   t_8861;
/* u2_3048 Output nets */
wire t_8862,   t_8863,   t_8864;
/* u2_3049 Output nets */
wire t_8865,   t_8866,   t_8867;
/* u2_3050 Output nets */
wire t_8868,   t_8869,   t_8870;
/* u2_3051 Output nets */
wire t_8871,   t_8872,   t_8873;
/* u1_3052 Output nets */
wire t_8874,   t_8875;
/* u2_3053 Output nets */
wire t_8876,   t_8877,   t_8878;
/* u2_3054 Output nets */
wire t_8879,   t_8880,   t_8881;
/* u2_3055 Output nets */
wire t_8882,   t_8883,   t_8884;
/* u2_3056 Output nets */
wire t_8885,   t_8886,   t_8887;
/* u2_3057 Output nets */
wire t_8888,   t_8889,   t_8890;
/* u1_3058 Output nets */
wire t_8891,   t_8892;
/* u2_3059 Output nets */
wire t_8893,   t_8894,   t_8895;
/* u2_3060 Output nets */
wire t_8896,   t_8897,   t_8898;
/* u2_3061 Output nets */
wire t_8899,   t_8900,   t_8901;
/* u2_3062 Output nets */
wire t_8902,   t_8903,   t_8904;
/* u2_3063 Output nets */
wire t_8905,   t_8906,   t_8907;
/* u1_3064 Output nets */
wire t_8908,   t_8909;
/* u2_3065 Output nets */
wire t_8910,   t_8911,   t_8912;
/* u2_3066 Output nets */
wire t_8913,   t_8914,   t_8915;
/* u2_3067 Output nets */
wire t_8916,   t_8917,   t_8918;
/* u2_3068 Output nets */
wire t_8919,   t_8920,   t_8921;
/* u2_3069 Output nets */
wire t_8922,   t_8923,   t_8924;
/* u1_3070 Output nets */
wire t_8925,   t_8926;
/* u2_3071 Output nets */
wire t_8927,   t_8928,   t_8929;
/* u2_3072 Output nets */
wire t_8930,   t_8931,   t_8932;
/* u2_3073 Output nets */
wire t_8933,   t_8934,   t_8935;
/* u2_3074 Output nets */
wire t_8936,   t_8937,   t_8938;
/* u2_3075 Output nets */
wire t_8939,   t_8940,   t_8941;
/* u1_3076 Output nets */
wire t_8942,   t_8943;
/* u2_3077 Output nets */
wire t_8944,   t_8945,   t_8946;
/* u2_3078 Output nets */
wire t_8947,   t_8948,   t_8949;
/* u2_3079 Output nets */
wire t_8950,   t_8951,   t_8952;
/* u2_3080 Output nets */
wire t_8953,   t_8954,   t_8955;
/* u2_3081 Output nets */
wire t_8956,   t_8957,   t_8958;
/* u1_3082 Output nets */
wire t_8959,   t_8960;
/* u2_3083 Output nets */
wire t_8961,   t_8962,   t_8963;
/* u2_3084 Output nets */
wire t_8964,   t_8965,   t_8966;
/* u2_3085 Output nets */
wire t_8967,   t_8968,   t_8969;
/* u2_3086 Output nets */
wire t_8970,   t_8971,   t_8972;
/* u2_3087 Output nets */
wire t_8973,   t_8974,   t_8975;
/* u1_3088 Output nets */
wire t_8976,   t_8977;
/* u2_3089 Output nets */
wire t_8978,   t_8979,   t_8980;
/* u2_3090 Output nets */
wire t_8981,   t_8982,   t_8983;
/* u2_3091 Output nets */
wire t_8984,   t_8985,   t_8986;
/* u2_3092 Output nets */
wire t_8987,   t_8988,   t_8989;
/* u2_3093 Output nets */
wire t_8990,   t_8991,   t_8992;
/* u1_3094 Output nets */
wire t_8993,   t_8994;
/* u2_3095 Output nets */
wire t_8995,   t_8996,   t_8997;
/* u2_3096 Output nets */
wire t_8998,   t_8999,   t_9000;
/* u2_3097 Output nets */
wire t_9001,   t_9002,   t_9003;
/* u2_3098 Output nets */
wire t_9004,   t_9005,   t_9006;
/* u2_3099 Output nets */
wire t_9007,   t_9008,   t_9009;
/* u0_3100 Output nets */
wire t_9010,   t_9011;
/* u2_3101 Output nets */
wire t_9012,   t_9013,   t_9014;
/* u2_3102 Output nets */
wire t_9015,   t_9016,   t_9017;
/* u2_3103 Output nets */
wire t_9018,   t_9019,   t_9020;
/* u2_3104 Output nets */
wire t_9021,   t_9022,   t_9023;
/* u2_3105 Output nets */
wire t_9024,   t_9025,   t_9026;
/* u0_3106 Output nets */
wire t_9027,   t_9028;
/* u2_3107 Output nets */
wire t_9029,   t_9030,   t_9031;
/* u2_3108 Output nets */
wire t_9032,   t_9033,   t_9034;
/* u2_3109 Output nets */
wire t_9035,   t_9036,   t_9037;
/* u2_3110 Output nets */
wire t_9038,   t_9039,   t_9040;
/* u2_3111 Output nets */
wire t_9041,   t_9042,   t_9043;
/* u0_3112 Output nets */
wire t_9044,   t_9045;
/* u2_3113 Output nets */
wire t_9046,   t_9047,   t_9048;
/* u2_3114 Output nets */
wire t_9049,   t_9050,   t_9051;
/* u2_3115 Output nets */
wire t_9052,   t_9053,   t_9054;
/* u2_3116 Output nets */
wire t_9055,   t_9056,   t_9057;
/* u2_3117 Output nets */
wire t_9058,   t_9059,   t_9060;
/* u0_3118 Output nets */
wire t_9061,   t_9062;
/* u2_3119 Output nets */
wire t_9063,   t_9064,   t_9065;
/* u2_3120 Output nets */
wire t_9066,   t_9067,   t_9068;
/* u2_3121 Output nets */
wire t_9069,   t_9070,   t_9071;
/* u2_3122 Output nets */
wire t_9072,   t_9073,   t_9074;
/* u2_3123 Output nets */
wire t_9075,   t_9076,   t_9077;
/* u0_3124 Output nets */
wire t_9078,   t_9079;
/* u2_3125 Output nets */
wire t_9080,   t_9081,   t_9082;
/* u2_3126 Output nets */
wire t_9083,   t_9084,   t_9085;
/* u2_3127 Output nets */
wire t_9086,   t_9087,   t_9088;
/* u2_3128 Output nets */
wire t_9089,   t_9090,   t_9091;
/* u2_3129 Output nets */
wire t_9092,   t_9093,   t_9094;
/* u2_3130 Output nets */
wire t_9095,   t_9096,   t_9097;
/* u2_3131 Output nets */
wire t_9098,   t_9099,   t_9100;
/* u2_3132 Output nets */
wire t_9101,   t_9102,   t_9103;
/* u2_3133 Output nets */
wire t_9104,   t_9105,   t_9106;
/* u2_3134 Output nets */
wire t_9107,   t_9108,   t_9109;
/* u2_3135 Output nets */
wire t_9110,   t_9111,   t_9112;
/* u2_3136 Output nets */
wire t_9113,   t_9114,   t_9115;
/* u2_3137 Output nets */
wire t_9116,   t_9117,   t_9118;
/* u2_3138 Output nets */
wire t_9119,   t_9120,   t_9121;
/* u2_3139 Output nets */
wire t_9122,   t_9123,   t_9124;
/* u2_3140 Output nets */
wire t_9125,   t_9126,   t_9127;
/* u2_3141 Output nets */
wire t_9128,   t_9129,   t_9130;
/* u2_3142 Output nets */
wire t_9131,   t_9132,   t_9133;
/* u2_3143 Output nets */
wire t_9134,   t_9135,   t_9136;
/* u1_3144 Output nets */
wire t_9137,   t_9138;
/* u2_3145 Output nets */
wire t_9139,   t_9140,   t_9141;
/* u2_3146 Output nets */
wire t_9142,   t_9143,   t_9144;
/* u2_3147 Output nets */
wire t_9145,   t_9146,   t_9147;
/* u2_3148 Output nets */
wire t_9148,   t_9149,   t_9150;
/* u1_3149 Output nets */
wire t_9151,   t_9152;
/* u2_3150 Output nets */
wire t_9153,   t_9154,   t_9155;
/* u2_3151 Output nets */
wire t_9156,   t_9157,   t_9158;
/* u2_3152 Output nets */
wire t_9159,   t_9160,   t_9161;
/* u2_3153 Output nets */
wire t_9162,   t_9163,   t_9164;
/* u1_3154 Output nets */
wire t_9165,   t_9166;
/* u2_3155 Output nets */
wire t_9167,   t_9168,   t_9169;
/* u2_3156 Output nets */
wire t_9170,   t_9171,   t_9172;
/* u2_3157 Output nets */
wire t_9173,   t_9174,   t_9175;
/* u2_3158 Output nets */
wire t_9176,   t_9177,   t_9178;
/* u1_3159 Output nets */
wire t_9179,   t_9180;
/* u2_3160 Output nets */
wire t_9181,   t_9182,   t_9183;
/* u2_3161 Output nets */
wire t_9184,   t_9185,   t_9186;
/* u2_3162 Output nets */
wire t_9187,   t_9188,   t_9189;
/* u2_3163 Output nets */
wire t_9190,   t_9191,   t_9192;
/* u1_3164 Output nets */
wire t_9193,   t_9194;
/* u2_3165 Output nets */
wire t_9195,   t_9196,   t_9197;
/* u2_3166 Output nets */
wire t_9198,   t_9199,   t_9200;
/* u2_3167 Output nets */
wire t_9201,   t_9202,   t_9203;
/* u2_3168 Output nets */
wire t_9204,   t_9205,   t_9206;
/* u1_3169 Output nets */
wire t_9207,   t_9208;
/* u2_3170 Output nets */
wire t_9209,   t_9210,   t_9211;
/* u2_3171 Output nets */
wire t_9212,   t_9213,   t_9214;
/* u2_3172 Output nets */
wire t_9215,   t_9216,   t_9217;
/* u2_3173 Output nets */
wire t_9218,   t_9219,   t_9220;
/* u1_3174 Output nets */
wire t_9221,   t_9222;
/* u2_3175 Output nets */
wire t_9223,   t_9224,   t_9225;
/* u2_3176 Output nets */
wire t_9226,   t_9227,   t_9228;
/* u2_3177 Output nets */
wire t_9229,   t_9230,   t_9231;
/* u2_3178 Output nets */
wire t_9232,   t_9233,   t_9234;
/* u1_3179 Output nets */
wire t_9235,   t_9236;
/* u2_3180 Output nets */
wire t_9237,   t_9238,   t_9239;
/* u2_3181 Output nets */
wire t_9240,   t_9241,   t_9242;
/* u2_3182 Output nets */
wire t_9243,   t_9244,   t_9245;
/* u2_3183 Output nets */
wire t_9246,   t_9247,   t_9248;
/* u0_3184 Output nets */
wire t_9249,   t_9250;
/* u2_3185 Output nets */
wire t_9251,   t_9252,   t_9253;
/* u2_3186 Output nets */
wire t_9254,   t_9255,   t_9256;
/* u2_3187 Output nets */
wire t_9257,   t_9258,   t_9259;
/* u2_3188 Output nets */
wire t_9260,   t_9261,   t_9262;
/* u0_3189 Output nets */
wire t_9263,   t_9264;
/* u2_3190 Output nets */
wire t_9265,   t_9266,   t_9267;
/* u2_3191 Output nets */
wire t_9268,   t_9269,   t_9270;
/* u2_3192 Output nets */
wire t_9271,   t_9272,   t_9273;
/* u2_3193 Output nets */
wire t_9274,   t_9275,   t_9276;
/* u0_3194 Output nets */
wire t_9277,   t_9278;
/* u2_3195 Output nets */
wire t_9279,   t_9280,   t_9281;
/* u2_3196 Output nets */
wire t_9282,   t_9283,   t_9284;
/* u2_3197 Output nets */
wire t_9285,   t_9286,   t_9287;
/* u2_3198 Output nets */
wire t_9288,   t_9289,   t_9290;
/* u0_3199 Output nets */
wire t_9291,   t_9292;
/* u2_3200 Output nets */
wire t_9293,   t_9294,   t_9295;
/* u2_3201 Output nets */
wire t_9296,   t_9297,   t_9298;
/* u2_3202 Output nets */
wire t_9299,   t_9300,   t_9301;
/* u2_3203 Output nets */
wire t_9302,   t_9303,   t_9304;
/* u0_3204 Output nets */
wire t_9305,   t_9306;
/* u2_3205 Output nets */
wire t_9307,   t_9308,   t_9309;
/* u2_3206 Output nets */
wire t_9310,   t_9311,   t_9312;
/* u2_3207 Output nets */
wire t_9313,   t_9314,   t_9315;
/* u2_3208 Output nets */
wire t_9316,   t_9317,   t_9318;
/* u2_3209 Output nets */
wire t_9319,   t_9320,   t_9321;
/* u2_3210 Output nets */
wire t_9322,   t_9323,   t_9324;
/* u2_3211 Output nets */
wire t_9325,   t_9326,   t_9327;
/* u2_3212 Output nets */
wire t_9328,   t_9329,   t_9330;
/* u2_3213 Output nets */
wire t_9331,   t_9332,   t_9333;
/* u2_3214 Output nets */
wire t_9334,   t_9335,   t_9336;
/* u2_3215 Output nets */
wire t_9337,   t_9338,   t_9339;
/* u2_3216 Output nets */
wire t_9340,   t_9341,   t_9342;
/* u2_3217 Output nets */
wire t_9343,   t_9344,   t_9345;
/* u2_3218 Output nets */
wire t_9346,   t_9347,   t_9348;
/* u2_3219 Output nets */
wire t_9349,   t_9350,   t_9351;
/* u1_3220 Output nets */
wire t_9352,   t_9353;
/* u2_3221 Output nets */
wire t_9354,   t_9355,   t_9356;
/* u2_3222 Output nets */
wire t_9357,   t_9358,   t_9359;
/* u2_3223 Output nets */
wire t_9360,   t_9361,   t_9362;
/* u1_3224 Output nets */
wire t_9363,   t_9364;
/* u2_3225 Output nets */
wire t_9365,   t_9366,   t_9367;
/* u2_3226 Output nets */
wire t_9368,   t_9369,   t_9370;
/* u2_3227 Output nets */
wire t_9371,   t_9372,   t_9373;
/* u1_3228 Output nets */
wire t_9374,   t_9375;
/* u2_3229 Output nets */
wire t_9376,   t_9377,   t_9378;
/* u2_3230 Output nets */
wire t_9379,   t_9380,   t_9381;
/* u2_3231 Output nets */
wire t_9382,   t_9383,   t_9384;
/* u1_3232 Output nets */
wire t_9385,   t_9386;
/* u2_3233 Output nets */
wire t_9387,   t_9388,   t_9389;
/* u2_3234 Output nets */
wire t_9390,   t_9391,   t_9392;
/* u2_3235 Output nets */
wire t_9393,   t_9394,   t_9395;
/* u1_3236 Output nets */
wire t_9396,   t_9397;
/* u2_3237 Output nets */
wire t_9398,   t_9399,   t_9400;
/* u2_3238 Output nets */
wire t_9401,   t_9402,   t_9403;
/* u2_3239 Output nets */
wire t_9404,   t_9405,   t_9406;
/* u1_3240 Output nets */
wire t_9407,   t_9408;
/* u2_3241 Output nets */
wire t_9409,   t_9410,   t_9411;
/* u2_3242 Output nets */
wire t_9412,   t_9413,   t_9414;
/* u2_3243 Output nets */
wire t_9415,   t_9416,   t_9417;
/* u1_3244 Output nets */
wire t_9418,   t_9419;
/* u2_3245 Output nets */
wire t_9420,   t_9421,   t_9422;
/* u2_3246 Output nets */
wire t_9423,   t_9424,   t_9425;
/* u2_3247 Output nets */
wire t_9426,   t_9427,   t_9428;
/* u1_3248 Output nets */
wire t_9429,   t_9430;
/* u2_3249 Output nets */
wire t_9431,   t_9432,   t_9433;
/* u2_3250 Output nets */
wire t_9434,   t_9435,   t_9436;
/* u2_3251 Output nets */
wire t_9437,   t_9438,   t_9439;
/* u0_3252 Output nets */
wire t_9440,   t_9441;
/* u2_3253 Output nets */
wire t_9442,   t_9443,   t_9444;
/* u2_3254 Output nets */
wire t_9445,   t_9446,   t_9447;
/* u2_3255 Output nets */
wire t_9448,   t_9449,   t_9450;
/* u0_3256 Output nets */
wire t_9451,   t_9452;
/* u2_3257 Output nets */
wire t_9453,   t_9454,   t_9455;
/* u2_3258 Output nets */
wire t_9456,   t_9457,   t_9458;
/* u2_3259 Output nets */
wire t_9459,   t_9460,   t_9461;
/* u0_3260 Output nets */
wire t_9462,   t_9463;
/* u2_3261 Output nets */
wire t_9464,   t_9465,   t_9466;
/* u2_3262 Output nets */
wire t_9467,   t_9468,   t_9469;
/* u2_3263 Output nets */
wire t_9470,   t_9471,   t_9472;
/* u0_3264 Output nets */
wire t_9473,   t_9474;
/* u2_3265 Output nets */
wire t_9475,   t_9476,   t_9477;
/* u2_3266 Output nets */
wire t_9478,   t_9479,   t_9480;
/* u2_3267 Output nets */
wire t_9481,   t_9482,   t_9483;
/* u0_3268 Output nets */
wire t_9484,   t_9485;
/* u2_3269 Output nets */
wire t_9486,   t_9487,   t_9488;
/* u2_3270 Output nets */
wire t_9489,   t_9490,   t_9491;
/* u2_3271 Output nets */
wire t_9492,   t_9493,   t_9494;
/* u2_3272 Output nets */
wire t_9495,   t_9496,   t_9497;
/* u2_3273 Output nets */
wire t_9498,   t_9499,   t_9500;
/* u2_3274 Output nets */
wire t_9501,   t_9502,   t_9503;
/* u2_3275 Output nets */
wire t_9504,   t_9505,   t_9506;
/* u2_3276 Output nets */
wire t_9507,   t_9508,   t_9509;
/* u2_3277 Output nets */
wire t_9510,   t_9511,   t_9512;
/* u2_3278 Output nets */
wire t_9513,   t_9514,   t_9515;
/* u2_3279 Output nets */
wire t_9516,   t_9517,   t_9518;
/* u1_3280 Output nets */
wire t_9519,   t_9520;
/* u2_3281 Output nets */
wire t_9521,   t_9522,   t_9523;
/* u2_3282 Output nets */
wire t_9524,   t_9525,   t_9526;
/* u1_3283 Output nets */
wire t_9527,   t_9528;
/* u2_3284 Output nets */
wire t_9529,   t_9530,   t_9531;
/* u2_3285 Output nets */
wire t_9532,   t_9533,   t_9534;
/* u1_3286 Output nets */
wire t_9535,   t_9536;
/* u2_3287 Output nets */
wire t_9537,   t_9538,   t_9539;
/* u2_3288 Output nets */
wire t_9540,   t_9541,   t_9542;
/* u1_3289 Output nets */
wire t_9543,   t_9544;
/* u2_3290 Output nets */
wire t_9545,   t_9546,   t_9547;
/* u2_3291 Output nets */
wire t_9548,   t_9549,   t_9550;
/* u1_3292 Output nets */
wire t_9551,   t_9552;
/* u2_3293 Output nets */
wire t_9553,   t_9554,   t_9555;
/* u2_3294 Output nets */
wire t_9556,   t_9557,   t_9558;
/* u1_3295 Output nets */
wire t_9559,   t_9560;
/* u2_3296 Output nets */
wire t_9561,   t_9562,   t_9563;
/* u2_3297 Output nets */
wire t_9564,   t_9565,   t_9566;
/* u1_3298 Output nets */
wire t_9567,   t_9568;
/* u2_3299 Output nets */
wire t_9569,   t_9570,   t_9571;
/* u2_3300 Output nets */
wire t_9572,   t_9573,   t_9574;
/* u1_3301 Output nets */
wire t_9575,   t_9576;
/* u2_3302 Output nets */
wire t_9577,   t_9578,   t_9579;
/* u2_3303 Output nets */
wire t_9580,   t_9581,   t_9582;
/* u0_3304 Output nets */
wire t_9583,   t_9584;
/* u2_3305 Output nets */
wire t_9585,   t_9586,   t_9587;
/* u2_3306 Output nets */
wire t_9588,   t_9589,   t_9590;
/* u0_3307 Output nets */
wire t_9591,   t_9592;
/* u2_3308 Output nets */
wire t_9593,   t_9594,   t_9595;
/* u2_3309 Output nets */
wire t_9596,   t_9597,   t_9598;
/* u0_3310 Output nets */
wire t_9599,   t_9600;
/* u2_3311 Output nets */
wire t_9601,   t_9602,   t_9603;
/* u2_3312 Output nets */
wire t_9604,   t_9605,   t_9606;
/* u0_3313 Output nets */
wire t_9607,   t_9608;
/* u2_3314 Output nets */
wire t_9609,   t_9610,   t_9611;
/* u2_3315 Output nets */
wire t_9612,   t_9613,   t_9614;
/* u0_3316 Output nets */
wire t_9615,   t_9616;
/* u2_3317 Output nets */
wire t_9617,   t_9618,   t_9619;
/* u2_3318 Output nets */
wire t_9620,   t_9621,   t_9622;
/* u2_3319 Output nets */
wire t_9623,   t_9624,   t_9625;
/* u2_3320 Output nets */
wire t_9626,   t_9627,   t_9628;
/* u2_3321 Output nets */
wire t_9629,   t_9630,   t_9631;
/* u2_3322 Output nets */
wire t_9632,   t_9633,   t_9634;
/* u2_3323 Output nets */
wire t_9635,   t_9636,   t_9637;
/* u1_3324 Output nets */
wire t_9638,   t_9639;
/* u2_3325 Output nets */
wire t_9640,   t_9641,   t_9642;
/* u1_3326 Output nets */
wire t_9643,   t_9644;
/* u2_3327 Output nets */
wire t_9645,   t_9646,   t_9647;
/* u1_3328 Output nets */
wire t_9648,   t_9649;
/* u2_3329 Output nets */
wire t_9650,   t_9651,   t_9652;
/* u1_3330 Output nets */
wire t_9653,   t_9654;
/* u2_3331 Output nets */
wire t_9655,   t_9656,   t_9657;
/* u1_3332 Output nets */
wire t_9658,   t_9659;
/* u2_3333 Output nets */
wire t_9660,   t_9661,   t_9662;
/* u1_3334 Output nets */
wire t_9663,   t_9664;
/* u2_3335 Output nets */
wire t_9665,   t_9666,   t_9667;
/* u1_3336 Output nets */
wire t_9668,   t_9669;
/* u2_3337 Output nets */
wire t_9670,   t_9671,   t_9672;
/* u1_3338 Output nets */
wire t_9673,   t_9674;
/* u2_3339 Output nets */
wire t_9675,   t_9676,   t_9677;
/* u0_3340 Output nets */
wire t_9678,   t_9679;
/* u2_3341 Output nets */
wire t_9680,   t_9681,   t_9682;
/* u0_3342 Output nets */
wire t_9683,   t_9684;
/* u2_3343 Output nets */
wire t_9685,   t_9686,   t_9687;
/* u0_3344 Output nets */
wire t_9688,   t_9689;
/* u2_3345 Output nets */
wire t_9690,   t_9691,   t_9692;
/* u0_3346 Output nets */
wire t_9693,   t_9694;
/* u2_3347 Output nets */
wire t_9695,   t_9696,   t_9697;
/* u0_3348 Output nets */
wire t_9698,   t_9699;
/* u2_3349 Output nets */
wire t_9700,   t_9701,   t_9702;
/* u2_3350 Output nets */
wire t_9703,   t_9704,   t_9705;
/* u2_3351 Output nets */
wire t_9706,   t_9707,   t_9708;
/* u1_3352 Output nets */
wire t_9709,   t_9710;
/* u1_3353 Output nets */
wire t_9711,   t_9712;
/* u1_3354 Output nets */
wire t_9713,   t_9714;
/* u1_3355 Output nets */
wire t_9715,   t_9716;
/* u1_3356 Output nets */
wire t_9717,   t_9718;
/* u0_3357 Output nets */
wire t_9719,   t_9720;
/* u1_3358 Output nets */
wire t_9721,   t_9722;
/* u0_3359 Output nets */
wire t_9723,   t_9724;
/* u0_3360 Output nets */
wire t_9725,   t_9726;
/* u0_3361 Output nets */
wire t_9727;

/* compress stage 2 */
half_adder u0_2206(.a(t_1), .b(s_1_0), .o(t_6441), .cout(t_6442));
half_adder u0_2207(.a(t_3), .b(t_4), .o(t_6443), .cout(t_6444));
compressor_3_2 u1_2208(.a(t_7), .b(t_9), .cin(s_5_2), .o(t_6445), .cout(t_6446));
half_adder u0_2209(.a(t_10), .b(t_11), .o(t_6447), .cout(t_6448));
half_adder u0_2210(.a(t_12), .b(t_14), .o(t_6449), .cout(t_6450));
compressor_3_2 u1_2211(.a(t_15), .b(t_20), .cin(t_17), .o(t_6451), .cout(t_6452));
compressor_3_2 u1_2212(.a(t_18), .b(t_25), .cin(t_22), .o(t_6453), .cout(t_6454));
compressor_4_2 u2_2213(.a(t_23), .b(t_30), .c(t_27), .d(s_10_6), .cin(t_6454), .o(t_6455), .co(t_6456), .cout(t_6457));
compressor_3_2 u1_2214(.a(t_35), .b(t_32), .cin(t_6457), .o(t_6458), .cout(t_6459));
compressor_3_2 u1_2215(.a(t_33), .b(t_40), .cin(t_37), .o(t_6460), .cout(t_6461));
compressor_4_2 u2_2216(.a(t_38), .b(t_46), .c(t_43), .d(s_13_6), .cin(t_6461), .o(t_6462), .co(t_6463), .cout(t_6464));
compressor_4_2 u2_2217(.a(t_44), .b(t_51), .c(t_48), .d(s_14_8), .cin(t_6464), .o(t_6465), .co(t_6466), .cout(t_6467));
compressor_4_2 u2_2218(.a(t_52), .b(t_49), .c(t_57), .d(t_54), .cin(t_6467), .o(t_6468), .co(t_6469), .cout(t_6470));
compressor_4_2 u2_2219(.a(t_55), .b(t_66), .c(t_63), .d(t_60), .cin(t_6470), .o(t_6471), .co(t_6472), .cout(t_6473));
compressor_4_2 u2_2220(.a(t_61), .b(t_74), .c(t_71), .d(t_68), .cin(t_6473), .o(t_6474), .co(t_6475), .cout(t_6476));
compressor_4_2 u2_2221(.a(t_82), .b(t_79), .c(t_76), .d(s_18_10), .cin(t_6476), .o(t_6477), .co(t_6478), .cout(t_6479));
half_adder u0_2222(.a(t_72), .b(t_69), .o(t_6480), .cout(t_6481));
compressor_4_2 u2_2223(.a(t_90), .b(t_87), .c(t_84), .d(t_6479), .cin(t_6481), .o(t_6482), .co(t_6483), .cout(t_6484));
half_adder u0_2224(.a(t_80), .b(t_77), .o(t_6485), .cout(t_6486));
compressor_4_2 u2_2225(.a(t_98), .b(t_95), .c(t_92), .d(t_6484), .cin(t_6486), .o(t_6487), .co(t_6488), .cout(t_6489));
half_adder u0_2226(.a(t_88), .b(t_85), .o(t_6490), .cout(t_6491));
compressor_4_2 u2_2227(.a(t_104), .b(t_101), .c(s_21_10), .d(t_6489), .cin(t_6491), .o(t_6492), .co(t_6493), .cout(t_6494));
compressor_3_2 u1_2228(.a(t_96), .b(t_93), .cin(t_107), .o(t_6495), .cout(t_6496));
compressor_4_2 u2_2229(.a(t_112), .b(t_109), .c(s_22_12), .d(t_6494), .cin(t_6496), .o(t_6497), .co(t_6498), .cout(t_6499));
compressor_3_2 u1_2230(.a(t_105), .b(t_102), .cin(t_115), .o(t_6500), .cout(t_6501));
compressor_4_2 u2_2231(.a(t_124), .b(t_121), .c(t_118), .d(t_6499), .cin(t_6501), .o(t_6502), .co(t_6503), .cout(t_6504));
compressor_3_2 u1_2232(.a(t_116), .b(t_113), .cin(t_110), .o(t_6505), .cout(t_6506));
compressor_4_2 u2_2233(.a(t_133), .b(t_130), .c(t_127), .d(t_6504), .cin(t_6506), .o(t_6507), .co(t_6508), .cout(t_6509));
compressor_3_2 u1_2234(.a(t_122), .b(t_119), .cin(t_136), .o(t_6510), .cout(t_6511));
compressor_4_2 u2_2235(.a(t_144), .b(t_141), .c(t_138), .d(t_6509), .cin(t_6511), .o(t_6512), .co(t_6513), .cout(t_6514));
compressor_3_2 u1_2236(.a(t_131), .b(t_128), .cin(t_147), .o(t_6515), .cout(t_6516));
compressor_4_2 u2_2237(.a(t_152), .b(t_149), .c(s_26_14), .d(t_6514), .cin(t_6516), .o(t_6517), .co(t_6518), .cout(t_6519));
compressor_4_2 u2_2238(.a(t_145), .b(t_142), .c(t_139), .d(t_158), .cin(t_155), .o(t_6520), .co(t_6521), .cout(t_6522));
compressor_4_2 u2_2239(.a(t_166), .b(t_163), .c(t_160), .d(t_6519), .cin(t_6522), .o(t_6523), .co(t_6524), .cout(t_6525));
compressor_3_2 u1_2240(.a(t_153), .b(t_150), .cin(t_169), .o(t_6526), .cout(t_6527));
compressor_4_2 u2_2241(.a(t_177), .b(t_174), .c(t_171), .d(t_6525), .cin(t_6527), .o(t_6528), .co(t_6529), .cout(t_6530));
compressor_3_2 u1_2242(.a(t_164), .b(t_161), .cin(t_180), .o(t_6531), .cout(t_6532));
compressor_4_2 u2_2243(.a(t_186), .b(t_183), .c(s_29_14), .d(t_6530), .cin(t_6532), .o(t_6533), .co(t_6534), .cout(t_6535));
compressor_4_2 u2_2244(.a(t_178), .b(t_175), .c(t_172), .d(t_192), .cin(t_189), .o(t_6536), .co(t_6537), .cout(t_6538));
compressor_4_2 u2_2245(.a(t_197), .b(t_194), .c(s_30_16), .d(t_6535), .cin(t_6538), .o(t_6539), .co(t_6540), .cout(t_6541));
compressor_4_2 u2_2246(.a(t_190), .b(t_187), .c(t_184), .d(t_203), .cin(t_200), .o(t_6542), .co(t_6543), .cout(t_6544));
compressor_4_2 u2_2247(.a(t_212), .b(t_209), .c(t_206), .d(t_6541), .cin(t_6544), .o(t_6545), .co(t_6546), .cout(t_6547));
compressor_4_2 u2_2248(.a(t_204), .b(t_201), .c(t_198), .d(t_195), .cin(t_215), .o(t_6548), .co(t_6549), .cout(t_6550));
compressor_4_2 u2_2249(.a(t_224), .b(t_221), .c(t_218), .d(t_6547), .cin(t_6550), .o(t_6551), .co(t_6552), .cout(t_6553));
compressor_4_2 u2_2250(.a(t_213), .b(t_210), .c(t_207), .d(t_230), .cin(t_227), .o(t_6554), .co(t_6555), .cout(t_6556));
compressor_4_2 u2_2251(.a(t_238), .b(t_235), .c(t_232), .d(t_6553), .cin(t_6556), .o(t_6557), .co(t_6558), .cout(t_6559));
compressor_4_2 u2_2252(.a(t_225), .b(t_222), .c(t_219), .d(t_244), .cin(t_241), .o(t_6560), .co(t_6561), .cout(t_6562));
compressor_4_2 u2_2253(.a(t_249), .b(t_246), .c(s_34_18), .d(t_6559), .cin(t_6562), .o(t_6563), .co(t_6564), .cout(t_6565));
compressor_4_2 u2_2254(.a(t_236), .b(t_233), .c(t_258), .d(t_255), .cin(t_252), .o(t_6566), .co(t_6567), .cout(t_6568));
half_adder u0_2255(.a(t_242), .b(t_239), .o(t_6569), .cout(t_6570));
compressor_4_2 u2_2256(.a(t_266), .b(t_263), .c(t_260), .d(t_6565), .cin(t_6568), .o(t_6571), .co(t_6572), .cout(t_6573));
compressor_4_2 u2_2257(.a(t_250), .b(t_247), .c(t_272), .d(t_269), .cin(t_6570), .o(t_6574), .co(t_6575), .cout(t_6576));
half_adder u0_2258(.a(t_256), .b(t_253), .o(t_6577), .cout(t_6578));
compressor_4_2 u2_2259(.a(t_280), .b(t_277), .c(t_274), .d(t_6573), .cin(t_6576), .o(t_6579), .co(t_6580), .cout(t_6581));
compressor_4_2 u2_2260(.a(t_264), .b(t_261), .c(t_286), .d(t_283), .cin(t_6578), .o(t_6582), .co(t_6583), .cout(t_6584));
half_adder u0_2261(.a(t_270), .b(t_267), .o(t_6585), .cout(t_6586));
compressor_4_2 u2_2262(.a(t_292), .b(t_289), .c(s_37_18), .d(t_6581), .cin(t_6584), .o(t_6587), .co(t_6588), .cout(t_6589));
compressor_4_2 u2_2263(.a(t_275), .b(t_301), .c(t_298), .d(t_295), .cin(t_6586), .o(t_6590), .co(t_6591), .cout(t_6592));
compressor_3_2 u1_2264(.a(t_284), .b(t_281), .cin(t_278), .o(t_6593), .cout(t_6594));
compressor_4_2 u2_2265(.a(t_306), .b(t_303), .c(s_38_20), .d(t_6589), .cin(t_6592), .o(t_6595), .co(t_6596), .cout(t_6597));
compressor_4_2 u2_2266(.a(t_290), .b(t_315), .c(t_312), .d(t_309), .cin(t_6594), .o(t_6598), .co(t_6599), .cout(t_6600));
compressor_3_2 u1_2267(.a(t_299), .b(t_296), .cin(t_293), .o(t_6601), .cout(t_6602));
compressor_4_2 u2_2268(.a(t_324), .b(t_321), .c(t_318), .d(t_6597), .cin(t_6600), .o(t_6603), .co(t_6604), .cout(t_6605));
compressor_4_2 u2_2269(.a(t_307), .b(t_304), .c(t_330), .d(t_327), .cin(t_6602), .o(t_6606), .co(t_6607), .cout(t_6608));
compressor_3_2 u1_2270(.a(t_316), .b(t_313), .cin(t_310), .o(t_6609), .cout(t_6610));
compressor_4_2 u2_2271(.a(t_339), .b(t_336), .c(t_333), .d(t_6605), .cin(t_6608), .o(t_6611), .co(t_6612), .cout(t_6613));
compressor_4_2 u2_2272(.a(t_319), .b(t_348), .c(t_345), .d(t_342), .cin(t_6610), .o(t_6614), .co(t_6615), .cout(t_6616));
compressor_3_2 u1_2273(.a(t_328), .b(t_325), .cin(t_322), .o(t_6617), .cout(t_6618));
compressor_4_2 u2_2274(.a(t_356), .b(t_353), .c(t_350), .d(t_6613), .cin(t_6616), .o(t_6619), .co(t_6620), .cout(t_6621));
compressor_4_2 u2_2275(.a(t_334), .b(t_365), .c(t_362), .d(t_359), .cin(t_6618), .o(t_6622), .co(t_6623), .cout(t_6624));
compressor_3_2 u1_2276(.a(t_343), .b(t_340), .cin(t_337), .o(t_6625), .cout(t_6626));
compressor_4_2 u2_2277(.a(t_370), .b(t_367), .c(s_42_22), .d(t_6621), .cin(t_6624), .o(t_6627), .co(t_6628), .cout(t_6629));
compressor_4_2 u2_2278(.a(t_382), .b(t_379), .c(t_376), .d(t_373), .cin(t_6626), .o(t_6630), .co(t_6631), .cout(t_6632));
compressor_4_2 u2_2279(.a(t_363), .b(t_360), .c(t_357), .d(t_354), .cin(t_351), .o(t_6633), .co(t_6634), .cout(t_6635));
compressor_4_2 u2_2280(.a(t_390), .b(t_387), .c(t_384), .d(t_6629), .cin(t_6632), .o(t_6636), .co(t_6637), .cout(t_6638));
compressor_4_2 u2_2281(.a(t_368), .b(t_399), .c(t_396), .d(t_393), .cin(t_6635), .o(t_6639), .co(t_6640), .cout(t_6641));
compressor_3_2 u1_2282(.a(t_377), .b(t_374), .cin(t_371), .o(t_6642), .cout(t_6643));
compressor_4_2 u2_2283(.a(t_407), .b(t_404), .c(t_401), .d(t_6638), .cin(t_6641), .o(t_6644), .co(t_6645), .cout(t_6646));
compressor_4_2 u2_2284(.a(t_385), .b(t_416), .c(t_413), .d(t_410), .cin(t_6643), .o(t_6647), .co(t_6648), .cout(t_6649));
compressor_3_2 u1_2285(.a(t_394), .b(t_391), .cin(t_388), .o(t_6650), .cout(t_6651));
compressor_4_2 u2_2286(.a(t_422), .b(t_419), .c(s_45_22), .d(t_6646), .cin(t_6649), .o(t_6652), .co(t_6653), .cout(t_6654));
compressor_4_2 u2_2287(.a(t_434), .b(t_431), .c(t_428), .d(t_425), .cin(t_6651), .o(t_6655), .co(t_6656), .cout(t_6657));
compressor_4_2 u2_2288(.a(t_414), .b(t_411), .c(t_408), .d(t_405), .cin(t_402), .o(t_6658), .co(t_6659), .cout(t_6660));
compressor_4_2 u2_2289(.a(t_439), .b(t_436), .c(s_46_24), .d(t_6654), .cin(t_6657), .o(t_6661), .co(t_6662), .cout(t_6663));
compressor_4_2 u2_2290(.a(t_451), .b(t_448), .c(t_445), .d(t_442), .cin(t_6660), .o(t_6664), .co(t_6665), .cout(t_6666));
compressor_4_2 u2_2291(.a(t_432), .b(t_429), .c(t_426), .d(t_423), .cin(t_420), .o(t_6667), .co(t_6668), .cout(t_6669));
compressor_4_2 u2_2292(.a(t_460), .b(t_457), .c(t_454), .d(t_6663), .cin(t_6666), .o(t_6670), .co(t_6671), .cout(t_6672));
compressor_4_2 u2_2293(.a(t_437), .b(t_469), .c(t_466), .d(t_463), .cin(t_6669), .o(t_6673), .co(t_6674), .cout(t_6675));
compressor_4_2 u2_2294(.a(t_452), .b(t_449), .c(t_446), .d(t_443), .cin(t_440), .o(t_6676), .co(t_6677), .cout(t_6678));
compressor_4_2 u2_2295(.a(t_478), .b(t_475), .c(t_472), .d(t_6672), .cin(t_6675), .o(t_6679), .co(t_6680), .cout(t_6681));
compressor_4_2 u2_2296(.a(t_490), .b(t_487), .c(t_484), .d(t_481), .cin(t_6678), .o(t_6682), .co(t_6683), .cout(t_6684));
compressor_4_2 u2_2297(.a(t_467), .b(t_464), .c(t_461), .d(t_458), .cin(t_455), .o(t_6685), .co(t_6686), .cout(t_6687));
compressor_4_2 u2_2298(.a(t_498), .b(t_495), .c(t_492), .d(t_6681), .cin(t_6684), .o(t_6688), .co(t_6689), .cout(t_6690));
compressor_4_2 u2_2299(.a(t_510), .b(t_507), .c(t_504), .d(t_501), .cin(t_6687), .o(t_6691), .co(t_6692), .cout(t_6693));
compressor_4_2 u2_2300(.a(t_485), .b(t_482), .c(t_479), .d(t_476), .cin(t_473), .o(t_6694), .co(t_6695), .cout(t_6696));
compressor_4_2 u2_2301(.a(t_515), .b(t_512), .c(s_50_26), .d(t_6690), .cin(t_6693), .o(t_6697), .co(t_6698), .cout(t_6699));
compressor_4_2 u2_2302(.a(t_527), .b(t_524), .c(t_521), .d(t_518), .cin(t_6696), .o(t_6700), .co(t_6701), .cout(t_6702));
compressor_4_2 u2_2303(.a(t_502), .b(t_499), .c(t_496), .d(t_493), .cin(t_530), .o(t_6703), .co(t_6704), .cout(t_6705));
half_adder u0_2304(.a(t_508), .b(t_505), .o(t_6706), .cout(t_6707));
compressor_4_2 u2_2305(.a(t_538), .b(t_535), .c(t_532), .d(t_6699), .cin(t_6702), .o(t_6708), .co(t_6709), .cout(t_6710));
compressor_4_2 u2_2306(.a(t_547), .b(t_544), .c(t_541), .d(t_6705), .cin(t_6707), .o(t_6711), .co(t_6712), .cout(t_6713));
compressor_4_2 u2_2307(.a(t_522), .b(t_519), .c(t_516), .d(t_513), .cin(t_550), .o(t_6714), .co(t_6715), .cout(t_6716));
half_adder u0_2308(.a(t_528), .b(t_525), .o(t_6717), .cout(t_6718));
compressor_4_2 u2_2309(.a(t_558), .b(t_555), .c(t_552), .d(t_6710), .cin(t_6713), .o(t_6719), .co(t_6720), .cout(t_6721));
compressor_4_2 u2_2310(.a(t_567), .b(t_564), .c(t_561), .d(t_6716), .cin(t_6718), .o(t_6722), .co(t_6723), .cout(t_6724));
compressor_4_2 u2_2311(.a(t_542), .b(t_539), .c(t_536), .d(t_533), .cin(t_570), .o(t_6725), .co(t_6726), .cout(t_6727));
half_adder u0_2312(.a(t_548), .b(t_545), .o(t_6728), .cout(t_6729));
compressor_4_2 u2_2313(.a(t_576), .b(t_573), .c(s_53_26), .d(t_6721), .cin(t_6724), .o(t_6730), .co(t_6731), .cout(t_6732));
compressor_4_2 u2_2314(.a(t_585), .b(t_582), .c(t_579), .d(t_6727), .cin(t_6729), .o(t_6733), .co(t_6734), .cout(t_6735));
compressor_4_2 u2_2315(.a(t_559), .b(t_556), .c(t_553), .d(t_591), .cin(t_588), .o(t_6736), .co(t_6737), .cout(t_6738));
compressor_3_2 u1_2316(.a(t_568), .b(t_565), .cin(t_562), .o(t_6739), .cout(t_6740));
compressor_4_2 u2_2317(.a(t_596), .b(t_593), .c(s_54_28), .d(t_6732), .cin(t_6735), .o(t_6741), .co(t_6742), .cout(t_6743));
compressor_4_2 u2_2318(.a(t_605), .b(t_602), .c(t_599), .d(t_6738), .cin(t_6740), .o(t_6744), .co(t_6745), .cout(t_6746));
compressor_4_2 u2_2319(.a(t_580), .b(t_577), .c(t_574), .d(t_611), .cin(t_608), .o(t_6747), .co(t_6748), .cout(t_6749));
compressor_3_2 u1_2320(.a(t_589), .b(t_586), .cin(t_583), .o(t_6750), .cout(t_6751));
compressor_4_2 u2_2321(.a(t_620), .b(t_617), .c(t_614), .d(t_6743), .cin(t_6746), .o(t_6752), .co(t_6753), .cout(t_6754));
compressor_4_2 u2_2322(.a(t_629), .b(t_626), .c(t_623), .d(t_6749), .cin(t_6751), .o(t_6755), .co(t_6756), .cout(t_6757));
compressor_4_2 u2_2323(.a(t_603), .b(t_600), .c(t_597), .d(t_594), .cin(t_632), .o(t_6758), .co(t_6759), .cout(t_6760));
compressor_3_2 u1_2324(.a(t_612), .b(t_609), .cin(t_606), .o(t_6761), .cout(t_6762));
compressor_4_2 u2_2325(.a(t_641), .b(t_638), .c(t_635), .d(t_6754), .cin(t_6757), .o(t_6763), .co(t_6764), .cout(t_6765));
compressor_4_2 u2_2326(.a(t_650), .b(t_647), .c(t_644), .d(t_6760), .cin(t_6762), .o(t_6766), .co(t_6767), .cout(t_6768));
compressor_4_2 u2_2327(.a(t_621), .b(t_618), .c(t_615), .d(t_656), .cin(t_653), .o(t_6769), .co(t_6770), .cout(t_6771));
compressor_3_2 u1_2328(.a(t_630), .b(t_627), .cin(t_624), .o(t_6772), .cout(t_6773));
compressor_4_2 u2_2329(.a(t_664), .b(t_661), .c(t_658), .d(t_6765), .cin(t_6768), .o(t_6774), .co(t_6775), .cout(t_6776));
compressor_4_2 u2_2330(.a(t_673), .b(t_670), .c(t_667), .d(t_6771), .cin(t_6773), .o(t_6777), .co(t_6778), .cout(t_6779));
compressor_4_2 u2_2331(.a(t_642), .b(t_639), .c(t_636), .d(t_679), .cin(t_676), .o(t_6780), .co(t_6781), .cout(t_6782));
compressor_3_2 u1_2332(.a(t_651), .b(t_648), .cin(t_645), .o(t_6783), .cout(t_6784));
compressor_4_2 u2_2333(.a(t_684), .b(t_681), .c(s_58_30), .d(t_6776), .cin(t_6779), .o(t_6785), .co(t_6786), .cout(t_6787));
compressor_4_2 u2_2334(.a(t_693), .b(t_690), .c(t_687), .d(t_6782), .cin(t_6784), .o(t_6788), .co(t_6789), .cout(t_6790));
compressor_4_2 u2_2335(.a(t_662), .b(t_659), .c(t_702), .d(t_699), .cin(t_696), .o(t_6791), .co(t_6792), .cout(t_6793));
compressor_4_2 u2_2336(.a(t_677), .b(t_674), .c(t_671), .d(t_668), .cin(t_665), .o(t_6794), .co(t_6795), .cout(t_6796));
compressor_4_2 u2_2337(.a(t_710), .b(t_707), .c(t_704), .d(t_6787), .cin(t_6790), .o(t_6797), .co(t_6798), .cout(t_6799));
compressor_4_2 u2_2338(.a(t_719), .b(t_716), .c(t_713), .d(t_6793), .cin(t_6796), .o(t_6800), .co(t_6801), .cout(t_6802));
compressor_4_2 u2_2339(.a(t_688), .b(t_685), .c(t_682), .d(t_725), .cin(t_722), .o(t_6803), .co(t_6804), .cout(t_6805));
compressor_3_2 u1_2340(.a(t_697), .b(t_694), .cin(t_691), .o(t_6806), .cout(t_6807));
compressor_4_2 u2_2341(.a(t_733), .b(t_730), .c(t_727), .d(t_6799), .cin(t_6802), .o(t_6808), .co(t_6809), .cout(t_6810));
compressor_4_2 u2_2342(.a(t_742), .b(t_739), .c(t_736), .d(t_6805), .cin(t_6807), .o(t_6811), .co(t_6812), .cout(t_6813));
compressor_4_2 u2_2343(.a(t_711), .b(t_708), .c(t_705), .d(t_748), .cin(t_745), .o(t_6814), .co(t_6815), .cout(t_6816));
compressor_3_2 u1_2344(.a(t_720), .b(t_717), .cin(t_714), .o(t_6817), .cout(t_6818));
compressor_4_2 u2_2345(.a(t_754), .b(t_751), .c(s_61_30), .d(t_6810), .cin(t_6813), .o(t_6819), .co(t_6820), .cout(t_6821));
compressor_4_2 u2_2346(.a(t_763), .b(t_760), .c(t_757), .d(t_6816), .cin(t_6818), .o(t_6822), .co(t_6823), .cout(t_6824));
compressor_4_2 u2_2347(.a(t_731), .b(t_728), .c(t_772), .d(t_769), .cin(t_766), .o(t_6825), .co(t_6826), .cout(t_6827));
compressor_4_2 u2_2348(.a(t_746), .b(t_743), .c(t_740), .d(t_737), .cin(t_734), .o(t_6828), .co(t_6829), .cout(t_6830));
compressor_4_2 u2_2349(.a(t_777), .b(t_774), .c(s_62_32), .d(t_6821), .cin(t_6824), .o(t_6831), .co(t_6832), .cout(t_6833));
compressor_4_2 u2_2350(.a(t_786), .b(t_783), .c(t_780), .d(t_6827), .cin(t_6830), .o(t_6834), .co(t_6835), .cout(t_6836));
compressor_4_2 u2_2351(.a(t_755), .b(t_752), .c(t_795), .d(t_792), .cin(t_789), .o(t_6837), .co(t_6838), .cout(t_6839));
compressor_4_2 u2_2352(.a(t_770), .b(t_767), .c(t_764), .d(t_761), .cin(t_758), .o(t_6840), .co(t_6841), .cout(t_6842));
compressor_4_2 u2_2353(.a(t_804), .b(t_801), .c(t_798), .d(t_6833), .cin(t_6836), .o(t_6843), .co(t_6844), .cout(t_6845));
compressor_4_2 u2_2354(.a(t_813), .b(t_810), .c(t_807), .d(t_6839), .cin(t_6842), .o(t_6846), .co(t_6847), .cout(t_6848));
compressor_4_2 u2_2355(.a(t_781), .b(t_778), .c(t_775), .d(t_819), .cin(t_816), .o(t_6849), .co(t_6850), .cout(t_6851));
compressor_4_2 u2_2356(.a(t_796), .b(t_793), .c(t_790), .d(t_787), .cin(t_784), .o(t_6852), .co(t_6853), .cout(t_6854));
compressor_4_2 u2_2357(.a(t_828), .b(t_825), .c(t_822), .d(t_6845), .cin(t_6848), .o(t_6855), .co(t_6856), .cout(t_6857));
compressor_4_2 u2_2358(.a(t_837), .b(t_834), .c(t_831), .d(t_6851), .cin(t_6854), .o(t_6858), .co(t_6859), .cout(t_6860));
compressor_4_2 u2_2359(.a(t_802), .b(t_799), .c(t_846), .d(t_843), .cin(t_840), .o(t_6861), .co(t_6862), .cout(t_6863));
compressor_4_2 u2_2360(.a(t_817), .b(t_814), .c(t_811), .d(t_808), .cin(t_805), .o(t_6864), .co(t_6865), .cout(t_6866));
compressor_4_2 u2_2361(.a(t_854), .b(t_851), .c(t_848), .d(t_6857), .cin(t_6860), .o(t_6867), .co(t_6868), .cout(t_6869));
compressor_4_2 u2_2362(.a(t_863), .b(t_860), .c(t_857), .d(t_6863), .cin(t_6866), .o(t_6870), .co(t_6871), .cout(t_6872));
compressor_4_2 u2_2363(.a(t_826), .b(t_823), .c(t_872), .d(t_869), .cin(t_866), .o(t_6873), .co(t_6874), .cout(t_6875));
compressor_4_2 u2_2364(.a(t_841), .b(t_838), .c(t_835), .d(t_832), .cin(t_829), .o(t_6876), .co(t_6877), .cout(t_6878));
compressor_4_2 u2_2365(.a(t_877), .b(t_874), .c(s_66_34), .d(t_6869), .cin(t_6872), .o(t_6879), .co(t_6880), .cout(t_6881));
compressor_4_2 u2_2366(.a(t_886), .b(t_883), .c(t_880), .d(t_6875), .cin(t_6878), .o(t_6882), .co(t_6883), .cout(t_6884));
compressor_4_2 u2_2367(.a(t_849), .b(t_898), .c(t_895), .d(t_892), .cin(t_889), .o(t_6885), .co(t_6886), .cout(t_6887));
compressor_4_2 u2_2368(.a(t_864), .b(t_861), .c(t_858), .d(t_855), .cin(t_852), .o(t_6888), .co(t_6889), .cout(t_6890));
half_adder u0_2369(.a(t_870), .b(t_867), .o(t_6891), .cout(t_6892));
compressor_4_2 u2_2370(.a(t_906), .b(t_903), .c(t_900), .d(t_6881), .cin(t_6884), .o(t_6893), .co(t_6894), .cout(t_6895));
compressor_4_2 u2_2371(.a(t_915), .b(t_912), .c(t_909), .d(t_6887), .cin(t_6890), .o(t_6896), .co(t_6897), .cout(t_6898));
compressor_4_2 u2_2372(.a(t_875), .b(t_924), .c(t_921), .d(t_918), .cin(t_6892), .o(t_6899), .co(t_6900), .cout(t_6901));
compressor_4_2 u2_2373(.a(t_890), .b(t_887), .c(t_884), .d(t_881), .cin(t_878), .o(t_6902), .co(t_6903), .cout(t_6904));
half_adder u0_2374(.a(t_896), .b(t_893), .o(t_6905), .cout(t_6906));
compressor_4_2 u2_2375(.a(t_932), .b(t_929), .c(t_926), .d(t_6895), .cin(t_6898), .o(t_6907), .co(t_6908), .cout(t_6909));
compressor_4_2 u2_2376(.a(t_941), .b(t_938), .c(t_935), .d(t_6901), .cin(t_6904), .o(t_6910), .co(t_6911), .cout(t_6912));
compressor_4_2 u2_2377(.a(t_901), .b(t_950), .c(t_947), .d(t_944), .cin(t_6906), .o(t_6913), .co(t_6914), .cout(t_6915));
compressor_4_2 u2_2378(.a(t_916), .b(t_913), .c(t_910), .d(t_907), .cin(t_904), .o(t_6916), .co(t_6917), .cout(t_6918));
half_adder u0_2379(.a(t_922), .b(t_919), .o(t_6919), .cout(t_6920));
compressor_4_2 u2_2380(.a(t_956), .b(t_953), .c(s_69_34), .d(t_6909), .cin(t_6912), .o(t_6921), .co(t_6922), .cout(t_6923));
compressor_4_2 u2_2381(.a(t_965), .b(t_962), .c(t_959), .d(t_6915), .cin(t_6918), .o(t_6924), .co(t_6925), .cout(t_6926));
compressor_4_2 u2_2382(.a(t_977), .b(t_974), .c(t_971), .d(t_968), .cin(t_6920), .o(t_6927), .co(t_6928), .cout(t_6929));
compressor_4_2 u2_2383(.a(t_939), .b(t_936), .c(t_933), .d(t_930), .cin(t_927), .o(t_6930), .co(t_6931), .cout(t_6932));
compressor_3_2 u1_2384(.a(t_948), .b(t_945), .cin(t_942), .o(t_6933), .cout(t_6934));
compressor_4_2 u2_2385(.a(t_982), .b(t_979), .c(s_70_36), .d(t_6923), .cin(t_6926), .o(t_6935), .co(t_6936), .cout(t_6937));
compressor_4_2 u2_2386(.a(t_991), .b(t_988), .c(t_985), .d(t_6929), .cin(t_6932), .o(t_6938), .co(t_6939), .cout(t_6940));
compressor_4_2 u2_2387(.a(t_1003), .b(t_1000), .c(t_997), .d(t_994), .cin(t_6934), .o(t_6941), .co(t_6942), .cout(t_6943));
compressor_4_2 u2_2388(.a(t_966), .b(t_963), .c(t_960), .d(t_957), .cin(t_954), .o(t_6944), .co(t_6945), .cout(t_6946));
compressor_3_2 u1_2389(.a(t_975), .b(t_972), .cin(t_969), .o(t_6947), .cout(t_6948));
compressor_4_2 u2_2390(.a(t_1012), .b(t_1009), .c(t_1006), .d(t_6937), .cin(t_6940), .o(t_6949), .co(t_6950), .cout(t_6951));
compressor_4_2 u2_2391(.a(t_1021), .b(t_1018), .c(t_1015), .d(t_6943), .cin(t_6946), .o(t_6952), .co(t_6953), .cout(t_6954));
compressor_4_2 u2_2392(.a(t_980), .b(t_1030), .c(t_1027), .d(t_1024), .cin(t_6948), .o(t_6955), .co(t_6956), .cout(t_6957));
compressor_4_2 u2_2393(.a(t_995), .b(t_992), .c(t_989), .d(t_986), .cin(t_983), .o(t_6958), .co(t_6959), .cout(t_6960));
compressor_3_2 u1_2394(.a(t_1004), .b(t_1001), .cin(t_998), .o(t_6961), .cout(t_6962));
compressor_4_2 u2_2395(.a(t_1039), .b(t_1036), .c(t_1033), .d(t_6951), .cin(t_6954), .o(t_6963), .co(t_6964), .cout(t_6965));
compressor_4_2 u2_2396(.a(t_1048), .b(t_1045), .c(t_1042), .d(t_6957), .cin(t_6960), .o(t_6966), .co(t_6967), .cout(t_6968));
compressor_4_2 u2_2397(.a(t_1060), .b(t_1057), .c(t_1054), .d(t_1051), .cin(t_6962), .o(t_6969), .co(t_6970), .cout(t_6971));
compressor_4_2 u2_2398(.a(t_1019), .b(t_1016), .c(t_1013), .d(t_1010), .cin(t_1007), .o(t_6972), .co(t_6973), .cout(t_6974));
compressor_3_2 u1_2399(.a(t_1028), .b(t_1025), .cin(t_1022), .o(t_6975), .cout(t_6976));
compressor_4_2 u2_2400(.a(t_1068), .b(t_1065), .c(t_1062), .d(t_6965), .cin(t_6968), .o(t_6977), .co(t_6978), .cout(t_6979));
compressor_4_2 u2_2401(.a(t_1077), .b(t_1074), .c(t_1071), .d(t_6971), .cin(t_6974), .o(t_6980), .co(t_6981), .cout(t_6982));
compressor_4_2 u2_2402(.a(t_1089), .b(t_1086), .c(t_1083), .d(t_1080), .cin(t_6976), .o(t_6983), .co(t_6984), .cout(t_6985));
compressor_4_2 u2_2403(.a(t_1046), .b(t_1043), .c(t_1040), .d(t_1037), .cin(t_1034), .o(t_6986), .co(t_6987), .cout(t_6988));
compressor_3_2 u1_2404(.a(t_1055), .b(t_1052), .cin(t_1049), .o(t_6989), .cout(t_6990));
compressor_4_2 u2_2405(.a(t_1094), .b(t_1091), .c(s_74_38), .d(t_6979), .cin(t_6982), .o(t_6991), .co(t_6992), .cout(t_6993));
compressor_4_2 u2_2406(.a(t_1103), .b(t_1100), .c(t_1097), .d(t_6985), .cin(t_6988), .o(t_6994), .co(t_6995), .cout(t_6996));
compressor_4_2 u2_2407(.a(t_1115), .b(t_1112), .c(t_1109), .d(t_1106), .cin(t_6990), .o(t_6997), .co(t_6998), .cout(t_6999));
compressor_4_2 u2_2408(.a(t_1072), .b(t_1069), .c(t_1066), .d(t_1063), .cin(t_1118), .o(t_7000), .co(t_7001), .cout(t_7002));
compressor_4_2 u2_2409(.a(t_1087), .b(t_1084), .c(t_1081), .d(t_1078), .cin(t_1075), .o(t_7003), .co(t_7004), .cout(t_7005));
compressor_4_2 u2_2410(.a(t_1126), .b(t_1123), .c(t_1120), .d(t_6993), .cin(t_6996), .o(t_7006), .co(t_7007), .cout(t_7008));
compressor_4_2 u2_2411(.a(t_1135), .b(t_1132), .c(t_1129), .d(t_6999), .cin(t_7002), .o(t_7009), .co(t_7010), .cout(t_7011));
compressor_4_2 u2_2412(.a(t_1147), .b(t_1144), .c(t_1141), .d(t_1138), .cin(t_7005), .o(t_7012), .co(t_7013), .cout(t_7014));
compressor_4_2 u2_2413(.a(t_1104), .b(t_1101), .c(t_1098), .d(t_1095), .cin(t_1092), .o(t_7015), .co(t_7016), .cout(t_7017));
compressor_3_2 u1_2414(.a(t_1113), .b(t_1110), .cin(t_1107), .o(t_7018), .cout(t_7019));
compressor_4_2 u2_2415(.a(t_1155), .b(t_1152), .c(t_1149), .d(t_7008), .cin(t_7011), .o(t_7020), .co(t_7021), .cout(t_7022));
compressor_4_2 u2_2416(.a(t_1164), .b(t_1161), .c(t_1158), .d(t_7014), .cin(t_7017), .o(t_7023), .co(t_7024), .cout(t_7025));
compressor_4_2 u2_2417(.a(t_1176), .b(t_1173), .c(t_1170), .d(t_1167), .cin(t_7019), .o(t_7026), .co(t_7027), .cout(t_7028));
compressor_4_2 u2_2418(.a(t_1133), .b(t_1130), .c(t_1127), .d(t_1124), .cin(t_1121), .o(t_7029), .co(t_7030), .cout(t_7031));
compressor_3_2 u1_2419(.a(t_1142), .b(t_1139), .cin(t_1136), .o(t_7032), .cout(t_7033));
compressor_4_2 u2_2420(.a(t_1182), .b(t_1179), .c(s_77_38), .d(t_7022), .cin(t_7025), .o(t_7034), .co(t_7035), .cout(t_7036));
compressor_4_2 u2_2421(.a(t_1191), .b(t_1188), .c(t_1185), .d(t_7028), .cin(t_7031), .o(t_7037), .co(t_7038), .cout(t_7039));
compressor_4_2 u2_2422(.a(t_1203), .b(t_1200), .c(t_1197), .d(t_1194), .cin(t_7033), .o(t_7040), .co(t_7041), .cout(t_7042));
compressor_4_2 u2_2423(.a(t_1159), .b(t_1156), .c(t_1153), .d(t_1150), .cin(t_1206), .o(t_7043), .co(t_7044), .cout(t_7045));
compressor_4_2 u2_2424(.a(t_1174), .b(t_1171), .c(t_1168), .d(t_1165), .cin(t_1162), .o(t_7046), .co(t_7047), .cout(t_7048));
compressor_4_2 u2_2425(.a(t_1211), .b(t_1208), .c(s_78_40), .d(t_7036), .cin(t_7039), .o(t_7049), .co(t_7050), .cout(t_7051));
compressor_4_2 u2_2426(.a(t_1220), .b(t_1217), .c(t_1214), .d(t_7042), .cin(t_7045), .o(t_7052), .co(t_7053), .cout(t_7054));
compressor_4_2 u2_2427(.a(t_1232), .b(t_1229), .c(t_1226), .d(t_1223), .cin(t_7048), .o(t_7055), .co(t_7056), .cout(t_7057));
compressor_4_2 u2_2428(.a(t_1189), .b(t_1186), .c(t_1183), .d(t_1180), .cin(t_1235), .o(t_7058), .co(t_7059), .cout(t_7060));
compressor_4_2 u2_2429(.a(t_1204), .b(t_1201), .c(t_1198), .d(t_1195), .cin(t_1192), .o(t_7061), .co(t_7062), .cout(t_7063));
compressor_4_2 u2_2430(.a(t_1244), .b(t_1241), .c(t_1238), .d(t_7051), .cin(t_7054), .o(t_7064), .co(t_7065), .cout(t_7066));
compressor_4_2 u2_2431(.a(t_1253), .b(t_1250), .c(t_1247), .d(t_7057), .cin(t_7060), .o(t_7067), .co(t_7068), .cout(t_7069));
compressor_4_2 u2_2432(.a(t_1265), .b(t_1262), .c(t_1259), .d(t_1256), .cin(t_7063), .o(t_7070), .co(t_7071), .cout(t_7072));
compressor_4_2 u2_2433(.a(t_1221), .b(t_1218), .c(t_1215), .d(t_1212), .cin(t_1209), .o(t_7073), .co(t_7074), .cout(t_7075));
compressor_4_2 u2_2434(.a(t_1236), .b(t_1233), .c(t_1230), .d(t_1227), .cin(t_1224), .o(t_7076), .co(t_7077), .cout(t_7078));
compressor_4_2 u2_2435(.a(t_1274), .b(t_1271), .c(t_1268), .d(t_7066), .cin(t_7069), .o(t_7079), .co(t_7080), .cout(t_7081));
compressor_4_2 u2_2436(.a(t_1283), .b(t_1280), .c(t_1277), .d(t_7072), .cin(t_7075), .o(t_7082), .co(t_7083), .cout(t_7084));
compressor_4_2 u2_2437(.a(t_1295), .b(t_1292), .c(t_1289), .d(t_1286), .cin(t_7078), .o(t_7085), .co(t_7086), .cout(t_7087));
compressor_4_2 u2_2438(.a(t_1248), .b(t_1245), .c(t_1242), .d(t_1239), .cin(t_1298), .o(t_7088), .co(t_7089), .cout(t_7090));
compressor_4_2 u2_2439(.a(t_1263), .b(t_1260), .c(t_1257), .d(t_1254), .cin(t_1251), .o(t_7091), .co(t_7092), .cout(t_7093));
compressor_4_2 u2_2440(.a(t_1306), .b(t_1303), .c(t_1300), .d(t_7081), .cin(t_7084), .o(t_7094), .co(t_7095), .cout(t_7096));
compressor_4_2 u2_2441(.a(t_1315), .b(t_1312), .c(t_1309), .d(t_7087), .cin(t_7090), .o(t_7097), .co(t_7098), .cout(t_7099));
compressor_4_2 u2_2442(.a(t_1327), .b(t_1324), .c(t_1321), .d(t_1318), .cin(t_7093), .o(t_7100), .co(t_7101), .cout(t_7102));
compressor_4_2 u2_2443(.a(t_1278), .b(t_1275), .c(t_1272), .d(t_1269), .cin(t_1330), .o(t_7103), .co(t_7104), .cout(t_7105));
compressor_4_2 u2_2444(.a(t_1293), .b(t_1290), .c(t_1287), .d(t_1284), .cin(t_1281), .o(t_7106), .co(t_7107), .cout(t_7108));
compressor_4_2 u2_2445(.a(t_1335), .b(t_1332), .c(s_82_42), .d(t_7096), .cin(t_7099), .o(t_7109), .co(t_7110), .cout(t_7111));
compressor_4_2 u2_2446(.a(t_1344), .b(t_1341), .c(t_1338), .d(t_7102), .cin(t_7105), .o(t_7112), .co(t_7113), .cout(t_7114));
compressor_4_2 u2_2447(.a(t_1356), .b(t_1353), .c(t_1350), .d(t_1347), .cin(t_7108), .o(t_7115), .co(t_7116), .cout(t_7117));
compressor_4_2 u2_2448(.a(t_1307), .b(t_1304), .c(t_1301), .d(t_1362), .cin(t_1359), .o(t_7118), .co(t_7119), .cout(t_7120));
compressor_4_2 u2_2449(.a(t_1322), .b(t_1319), .c(t_1316), .d(t_1313), .cin(t_1310), .o(t_7121), .co(t_7122), .cout(t_7123));
half_adder u0_2450(.a(t_1328), .b(t_1325), .o(t_7124), .cout(t_7125));
compressor_4_2 u2_2451(.a(t_1370), .b(t_1367), .c(t_1364), .d(t_7111), .cin(t_7114), .o(t_7126), .co(t_7127), .cout(t_7128));
compressor_4_2 u2_2452(.a(t_1379), .b(t_1376), .c(t_1373), .d(t_7117), .cin(t_7120), .o(t_7129), .co(t_7130), .cout(t_7131));
compressor_4_2 u2_2453(.a(t_1388), .b(t_1385), .c(t_1382), .d(t_7123), .cin(t_7125), .o(t_7132), .co(t_7133), .cout(t_7134));
compressor_4_2 u2_2454(.a(t_1339), .b(t_1336), .c(t_1333), .d(t_1394), .cin(t_1391), .o(t_7135), .co(t_7136), .cout(t_7137));
compressor_4_2 u2_2455(.a(t_1354), .b(t_1351), .c(t_1348), .d(t_1345), .cin(t_1342), .o(t_7138), .co(t_7139), .cout(t_7140));
half_adder u0_2456(.a(t_1360), .b(t_1357), .o(t_7141), .cout(t_7142));
compressor_4_2 u2_2457(.a(t_1402), .b(t_1399), .c(t_1396), .d(t_7128), .cin(t_7131), .o(t_7143), .co(t_7144), .cout(t_7145));
compressor_4_2 u2_2458(.a(t_1411), .b(t_1408), .c(t_1405), .d(t_7134), .cin(t_7137), .o(t_7146), .co(t_7147), .cout(t_7148));
compressor_4_2 u2_2459(.a(t_1420), .b(t_1417), .c(t_1414), .d(t_7140), .cin(t_7142), .o(t_7149), .co(t_7150), .cout(t_7151));
compressor_4_2 u2_2460(.a(t_1371), .b(t_1368), .c(t_1365), .d(t_1426), .cin(t_1423), .o(t_7152), .co(t_7153), .cout(t_7154));
compressor_4_2 u2_2461(.a(t_1386), .b(t_1383), .c(t_1380), .d(t_1377), .cin(t_1374), .o(t_7155), .co(t_7156), .cout(t_7157));
half_adder u0_2462(.a(t_1392), .b(t_1389), .o(t_7158), .cout(t_7159));
compressor_4_2 u2_2463(.a(t_1432), .b(t_1429), .c(s_85_42), .d(t_7145), .cin(t_7148), .o(t_7160), .co(t_7161), .cout(t_7162));
compressor_4_2 u2_2464(.a(t_1441), .b(t_1438), .c(t_1435), .d(t_7151), .cin(t_7154), .o(t_7163), .co(t_7164), .cout(t_7165));
compressor_4_2 u2_2465(.a(t_1450), .b(t_1447), .c(t_1444), .d(t_7157), .cin(t_7159), .o(t_7166), .co(t_7167), .cout(t_7168));
compressor_4_2 u2_2466(.a(t_1400), .b(t_1397), .c(t_1459), .d(t_1456), .cin(t_1453), .o(t_7169), .co(t_7170), .cout(t_7171));
compressor_4_2 u2_2467(.a(t_1415), .b(t_1412), .c(t_1409), .d(t_1406), .cin(t_1403), .o(t_7172), .co(t_7173), .cout(t_7174));
compressor_3_2 u1_2468(.a(t_1424), .b(t_1421), .cin(t_1418), .o(t_7175), .cout(t_7176));
compressor_4_2 u2_2469(.a(t_1464), .b(t_1461), .c(s_86_44), .d(t_7162), .cin(t_7165), .o(t_7177), .co(t_7178), .cout(t_7179));
compressor_4_2 u2_2470(.a(t_1473), .b(t_1470), .c(t_1467), .d(t_7168), .cin(t_7171), .o(t_7180), .co(t_7181), .cout(t_7182));
compressor_4_2 u2_2471(.a(t_1482), .b(t_1479), .c(t_1476), .d(t_7174), .cin(t_7176), .o(t_7183), .co(t_7184), .cout(t_7185));
compressor_4_2 u2_2472(.a(t_1433), .b(t_1430), .c(t_1491), .d(t_1488), .cin(t_1485), .o(t_7186), .co(t_7187), .cout(t_7188));
compressor_4_2 u2_2473(.a(t_1448), .b(t_1445), .c(t_1442), .d(t_1439), .cin(t_1436), .o(t_7189), .co(t_7190), .cout(t_7191));
compressor_3_2 u1_2474(.a(t_1457), .b(t_1454), .cin(t_1451), .o(t_7192), .cout(t_7193));
compressor_4_2 u2_2475(.a(t_1500), .b(t_1497), .c(t_1494), .d(t_7179), .cin(t_7182), .o(t_7194), .co(t_7195), .cout(t_7196));
compressor_4_2 u2_2476(.a(t_1509), .b(t_1506), .c(t_1503), .d(t_7185), .cin(t_7188), .o(t_7197), .co(t_7198), .cout(t_7199));
compressor_4_2 u2_2477(.a(t_1518), .b(t_1515), .c(t_1512), .d(t_7191), .cin(t_7193), .o(t_7200), .co(t_7201), .cout(t_7202));
compressor_4_2 u2_2478(.a(t_1468), .b(t_1465), .c(t_1462), .d(t_1524), .cin(t_1521), .o(t_7203), .co(t_7204), .cout(t_7205));
compressor_4_2 u2_2479(.a(t_1483), .b(t_1480), .c(t_1477), .d(t_1474), .cin(t_1471), .o(t_7206), .co(t_7207), .cout(t_7208));
compressor_3_2 u1_2480(.a(t_1492), .b(t_1489), .cin(t_1486), .o(t_7209), .cout(t_7210));
compressor_4_2 u2_2481(.a(t_1533), .b(t_1530), .c(t_1527), .d(t_7196), .cin(t_7199), .o(t_7211), .co(t_7212), .cout(t_7213));
compressor_4_2 u2_2482(.a(t_1542), .b(t_1539), .c(t_1536), .d(t_7202), .cin(t_7205), .o(t_7214), .co(t_7215), .cout(t_7216));
compressor_4_2 u2_2483(.a(t_1551), .b(t_1548), .c(t_1545), .d(t_7208), .cin(t_7210), .o(t_7217), .co(t_7218), .cout(t_7219));
compressor_4_2 u2_2484(.a(t_1498), .b(t_1495), .c(t_1560), .d(t_1557), .cin(t_1554), .o(t_7220), .co(t_7221), .cout(t_7222));
compressor_4_2 u2_2485(.a(t_1513), .b(t_1510), .c(t_1507), .d(t_1504), .cin(t_1501), .o(t_7223), .co(t_7224), .cout(t_7225));
compressor_3_2 u1_2486(.a(t_1522), .b(t_1519), .cin(t_1516), .o(t_7226), .cout(t_7227));
compressor_4_2 u2_2487(.a(t_1568), .b(t_1565), .c(t_1562), .d(t_7213), .cin(t_7216), .o(t_7228), .co(t_7229), .cout(t_7230));
compressor_4_2 u2_2488(.a(t_1577), .b(t_1574), .c(t_1571), .d(t_7219), .cin(t_7222), .o(t_7231), .co(t_7232), .cout(t_7233));
compressor_4_2 u2_2489(.a(t_1586), .b(t_1583), .c(t_1580), .d(t_7225), .cin(t_7227), .o(t_7234), .co(t_7235), .cout(t_7236));
compressor_4_2 u2_2490(.a(t_1531), .b(t_1528), .c(t_1595), .d(t_1592), .cin(t_1589), .o(t_7237), .co(t_7238), .cout(t_7239));
compressor_4_2 u2_2491(.a(t_1546), .b(t_1543), .c(t_1540), .d(t_1537), .cin(t_1534), .o(t_7240), .co(t_7241), .cout(t_7242));
compressor_3_2 u1_2492(.a(t_1555), .b(t_1552), .cin(t_1549), .o(t_7243), .cout(t_7244));
compressor_4_2 u2_2493(.a(t_1600), .b(t_1597), .c(s_90_46), .d(t_7230), .cin(t_7233), .o(t_7245), .co(t_7246), .cout(t_7247));
compressor_4_2 u2_2494(.a(t_1609), .b(t_1606), .c(t_1603), .d(t_7236), .cin(t_7239), .o(t_7248), .co(t_7249), .cout(t_7250));
compressor_4_2 u2_2495(.a(t_1618), .b(t_1615), .c(t_1612), .d(t_7242), .cin(t_7244), .o(t_7251), .co(t_7252), .cout(t_7253));
compressor_4_2 u2_2496(.a(t_1563), .b(t_1630), .c(t_1627), .d(t_1624), .cin(t_1621), .o(t_7254), .co(t_7255), .cout(t_7256));
compressor_4_2 u2_2497(.a(t_1578), .b(t_1575), .c(t_1572), .d(t_1569), .cin(t_1566), .o(t_7257), .co(t_7258), .cout(t_7259));
compressor_4_2 u2_2498(.a(t_1593), .b(t_1590), .c(t_1587), .d(t_1584), .cin(t_1581), .o(t_7260), .co(t_7261), .cout(t_7262));
compressor_4_2 u2_2499(.a(t_1638), .b(t_1635), .c(t_1632), .d(t_7247), .cin(t_7250), .o(t_7263), .co(t_7264), .cout(t_7265));
compressor_4_2 u2_2500(.a(t_1647), .b(t_1644), .c(t_1641), .d(t_7253), .cin(t_7256), .o(t_7266), .co(t_7267), .cout(t_7268));
compressor_4_2 u2_2501(.a(t_1656), .b(t_1653), .c(t_1650), .d(t_7259), .cin(t_7262), .o(t_7269), .co(t_7270), .cout(t_7271));
compressor_4_2 u2_2502(.a(t_1601), .b(t_1598), .c(t_1665), .d(t_1662), .cin(t_1659), .o(t_7272), .co(t_7273), .cout(t_7274));
compressor_4_2 u2_2503(.a(t_1616), .b(t_1613), .c(t_1610), .d(t_1607), .cin(t_1604), .o(t_7275), .co(t_7276), .cout(t_7277));
compressor_3_2 u1_2504(.a(t_1625), .b(t_1622), .cin(t_1619), .o(t_7278), .cout(t_7279));
compressor_4_2 u2_2505(.a(t_1673), .b(t_1670), .c(t_1667), .d(t_7265), .cin(t_7268), .o(t_7280), .co(t_7281), .cout(t_7282));
compressor_4_2 u2_2506(.a(t_1682), .b(t_1679), .c(t_1676), .d(t_7271), .cin(t_7274), .o(t_7283), .co(t_7284), .cout(t_7285));
compressor_4_2 u2_2507(.a(t_1691), .b(t_1688), .c(t_1685), .d(t_7277), .cin(t_7279), .o(t_7286), .co(t_7287), .cout(t_7288));
compressor_4_2 u2_2508(.a(t_1636), .b(t_1633), .c(t_1700), .d(t_1697), .cin(t_1694), .o(t_7289), .co(t_7290), .cout(t_7291));
compressor_4_2 u2_2509(.a(t_1651), .b(t_1648), .c(t_1645), .d(t_1642), .cin(t_1639), .o(t_7292), .co(t_7293), .cout(t_7294));
compressor_3_2 u1_2510(.a(t_1660), .b(t_1657), .cin(t_1654), .o(t_7295), .cout(t_7296));
compressor_4_2 u2_2511(.a(t_1706), .b(t_1703), .c(s_93_46), .d(t_7282), .cin(t_7285), .o(t_7297), .co(t_7298), .cout(t_7299));
compressor_4_2 u2_2512(.a(t_1715), .b(t_1712), .c(t_1709), .d(t_7288), .cin(t_7291), .o(t_7300), .co(t_7301), .cout(t_7302));
compressor_4_2 u2_2513(.a(t_1724), .b(t_1721), .c(t_1718), .d(t_7294), .cin(t_7296), .o(t_7303), .co(t_7304), .cout(t_7305));
compressor_4_2 u2_2514(.a(t_1668), .b(t_1736), .c(t_1733), .d(t_1730), .cin(t_1727), .o(t_7306), .co(t_7307), .cout(t_7308));
compressor_4_2 u2_2515(.a(t_1683), .b(t_1680), .c(t_1677), .d(t_1674), .cin(t_1671), .o(t_7309), .co(t_7310), .cout(t_7311));
compressor_4_2 u2_2516(.a(t_1698), .b(t_1695), .c(t_1692), .d(t_1689), .cin(t_1686), .o(t_7312), .co(t_7313), .cout(t_7314));
compressor_4_2 u2_2517(.a(t_1741), .b(t_1738), .c(s_94_48), .d(t_7299), .cin(t_7302), .o(t_7315), .co(t_7316), .cout(t_7317));
compressor_4_2 u2_2518(.a(t_1750), .b(t_1747), .c(t_1744), .d(t_7305), .cin(t_7308), .o(t_7318), .co(t_7319), .cout(t_7320));
compressor_4_2 u2_2519(.a(t_1759), .b(t_1756), .c(t_1753), .d(t_7311), .cin(t_7314), .o(t_7321), .co(t_7322), .cout(t_7323));
compressor_4_2 u2_2520(.a(t_1704), .b(t_1771), .c(t_1768), .d(t_1765), .cin(t_1762), .o(t_7324), .co(t_7325), .cout(t_7326));
compressor_4_2 u2_2521(.a(t_1719), .b(t_1716), .c(t_1713), .d(t_1710), .cin(t_1707), .o(t_7327), .co(t_7328), .cout(t_7329));
compressor_4_2 u2_2522(.a(t_1734), .b(t_1731), .c(t_1728), .d(t_1725), .cin(t_1722), .o(t_7330), .co(t_7331), .cout(t_7332));
compressor_4_2 u2_2523(.a(t_1780), .b(t_1777), .c(t_1774), .d(t_7317), .cin(t_7320), .o(t_7333), .co(t_7334), .cout(t_7335));
compressor_4_2 u2_2524(.a(t_1789), .b(t_1786), .c(t_1783), .d(t_7323), .cin(t_7326), .o(t_7336), .co(t_7337), .cout(t_7338));
compressor_4_2 u2_2525(.a(t_1798), .b(t_1795), .c(t_1792), .d(t_7329), .cin(t_7332), .o(t_7339), .co(t_7340), .cout(t_7341));
compressor_4_2 u2_2526(.a(t_1742), .b(t_1739), .c(t_1807), .d(t_1804), .cin(t_1801), .o(t_7342), .co(t_7343), .cout(t_7344));
compressor_4_2 u2_2527(.a(t_1757), .b(t_1754), .c(t_1751), .d(t_1748), .cin(t_1745), .o(t_7345), .co(t_7346), .cout(t_7347));
compressor_4_2 u2_2528(.a(t_1772), .b(t_1769), .c(t_1766), .d(t_1763), .cin(t_1760), .o(t_7348), .co(t_7349), .cout(t_7350));
compressor_4_2 u2_2529(.a(t_1816), .b(t_1813), .c(t_1810), .d(t_7335), .cin(t_7338), .o(t_7351), .co(t_7352), .cout(t_7353));
compressor_4_2 u2_2530(.a(t_1825), .b(t_1822), .c(t_1819), .d(t_7341), .cin(t_7344), .o(t_7354), .co(t_7355), .cout(t_7356));
compressor_4_2 u2_2531(.a(t_1834), .b(t_1831), .c(t_1828), .d(t_7347), .cin(t_7350), .o(t_7357), .co(t_7358), .cout(t_7359));
compressor_4_2 u2_2532(.a(t_1775), .b(t_1846), .c(t_1843), .d(t_1840), .cin(t_1837), .o(t_7360), .co(t_7361), .cout(t_7362));
compressor_4_2 u2_2533(.a(t_1790), .b(t_1787), .c(t_1784), .d(t_1781), .cin(t_1778), .o(t_7363), .co(t_7364), .cout(t_7365));
compressor_4_2 u2_2534(.a(t_1805), .b(t_1802), .c(t_1799), .d(t_1796), .cin(t_1793), .o(t_7366), .co(t_7367), .cout(t_7368));
compressor_4_2 u2_2535(.a(t_1854), .b(t_1851), .c(t_1848), .d(t_7353), .cin(t_7356), .o(t_7369), .co(t_7370), .cout(t_7371));
compressor_4_2 u2_2536(.a(t_1863), .b(t_1860), .c(t_1857), .d(t_7359), .cin(t_7362), .o(t_7372), .co(t_7373), .cout(t_7374));
compressor_4_2 u2_2537(.a(t_1872), .b(t_1869), .c(t_1866), .d(t_7365), .cin(t_7368), .o(t_7375), .co(t_7376), .cout(t_7377));
compressor_4_2 u2_2538(.a(t_1811), .b(t_1884), .c(t_1881), .d(t_1878), .cin(t_1875), .o(t_7378), .co(t_7379), .cout(t_7380));
compressor_4_2 u2_2539(.a(t_1826), .b(t_1823), .c(t_1820), .d(t_1817), .cin(t_1814), .o(t_7381), .co(t_7382), .cout(t_7383));
compressor_4_2 u2_2540(.a(t_1841), .b(t_1838), .c(t_1835), .d(t_1832), .cin(t_1829), .o(t_7384), .co(t_7385), .cout(t_7386));
compressor_4_2 u2_2541(.a(t_1889), .b(t_1886), .c(s_98_50), .d(t_7371), .cin(t_7374), .o(t_7387), .co(t_7388), .cout(t_7389));
compressor_4_2 u2_2542(.a(t_1898), .b(t_1895), .c(t_1892), .d(t_7377), .cin(t_7380), .o(t_7390), .co(t_7391), .cout(t_7392));
compressor_4_2 u2_2543(.a(t_1907), .b(t_1904), .c(t_1901), .d(t_7383), .cin(t_7386), .o(t_7393), .co(t_7394), .cout(t_7395));
compressor_4_2 u2_2544(.a(t_1922), .b(t_1919), .c(t_1916), .d(t_1913), .cin(t_1910), .o(t_7396), .co(t_7397), .cout(t_7398));
compressor_4_2 u2_2545(.a(t_1861), .b(t_1858), .c(t_1855), .d(t_1852), .cin(t_1849), .o(t_7399), .co(t_7400), .cout(t_7401));
compressor_4_2 u2_2546(.a(t_1876), .b(t_1873), .c(t_1870), .d(t_1867), .cin(t_1864), .o(t_7402), .co(t_7403), .cout(t_7404));
half_adder u0_2547(.a(t_1882), .b(t_1879), .o(t_7405), .cout(t_7406));
compressor_4_2 u2_2548(.a(t_1930), .b(t_1927), .c(t_1924), .d(t_7389), .cin(t_7392), .o(t_7407), .co(t_7408), .cout(t_7409));
compressor_4_2 u2_2549(.a(t_1939), .b(t_1936), .c(t_1933), .d(t_7395), .cin(t_7398), .o(t_7410), .co(t_7411), .cout(t_7412));
compressor_4_2 u2_2550(.a(t_1948), .b(t_1945), .c(t_1942), .d(t_7401), .cin(t_7404), .o(t_7413), .co(t_7414), .cout(t_7415));
compressor_4_2 u2_2551(.a(t_1960), .b(t_1957), .c(t_1954), .d(t_1951), .cin(t_7406), .o(t_7416), .co(t_7417), .cout(t_7418));
compressor_4_2 u2_2552(.a(t_1899), .b(t_1896), .c(t_1893), .d(t_1890), .cin(t_1887), .o(t_7419), .co(t_7420), .cout(t_7421));
compressor_4_2 u2_2553(.a(t_1914), .b(t_1911), .c(t_1908), .d(t_1905), .cin(t_1902), .o(t_7422), .co(t_7423), .cout(t_7424));
half_adder u0_2554(.a(t_1920), .b(t_1917), .o(t_7425), .cout(t_7426));
compressor_4_2 u2_2555(.a(t_1968), .b(t_1965), .c(t_1962), .d(t_7409), .cin(t_7412), .o(t_7427), .co(t_7428), .cout(t_7429));
compressor_4_2 u2_2556(.a(t_1977), .b(t_1974), .c(t_1971), .d(t_7415), .cin(t_7418), .o(t_7430), .co(t_7431), .cout(t_7432));
compressor_4_2 u2_2557(.a(t_1986), .b(t_1983), .c(t_1980), .d(t_7421), .cin(t_7424), .o(t_7433), .co(t_7434), .cout(t_7435));
compressor_4_2 u2_2558(.a(t_1998), .b(t_1995), .c(t_1992), .d(t_1989), .cin(t_7426), .o(t_7436), .co(t_7437), .cout(t_7438));
compressor_4_2 u2_2559(.a(t_1937), .b(t_1934), .c(t_1931), .d(t_1928), .cin(t_1925), .o(t_7439), .co(t_7440), .cout(t_7441));
compressor_4_2 u2_2560(.a(t_1952), .b(t_1949), .c(t_1946), .d(t_1943), .cin(t_1940), .o(t_7442), .co(t_7443), .cout(t_7444));
half_adder u0_2561(.a(t_1958), .b(t_1955), .o(t_7445), .cout(t_7446));
compressor_4_2 u2_2562(.a(t_2004), .b(t_2001), .c(s_101_50), .d(t_7429), .cin(t_7432), .o(t_7447), .co(t_7448), .cout(t_7449));
compressor_4_2 u2_2563(.a(t_2013), .b(t_2010), .c(t_2007), .d(t_7435), .cin(t_7438), .o(t_7450), .co(t_7451), .cout(t_7452));
compressor_4_2 u2_2564(.a(t_2022), .b(t_2019), .c(t_2016), .d(t_7441), .cin(t_7444), .o(t_7453), .co(t_7454), .cout(t_7455));
compressor_4_2 u2_2565(.a(t_2034), .b(t_2031), .c(t_2028), .d(t_2025), .cin(t_7446), .o(t_7456), .co(t_7457), .cout(t_7458));
compressor_4_2 u2_2566(.a(t_1972), .b(t_1969), .c(t_1966), .d(t_1963), .cin(t_2037), .o(t_7459), .co(t_7460), .cout(t_7461));
compressor_4_2 u2_2567(.a(t_1987), .b(t_1984), .c(t_1981), .d(t_1978), .cin(t_1975), .o(t_7462), .co(t_7463), .cout(t_7464));
compressor_3_2 u1_2568(.a(t_1996), .b(t_1993), .cin(t_1990), .o(t_7465), .cout(t_7466));
compressor_4_2 u2_2569(.a(t_2042), .b(t_2039), .c(s_102_52), .d(t_7449), .cin(t_7452), .o(t_7467), .co(t_7468), .cout(t_7469));
compressor_4_2 u2_2570(.a(t_2051), .b(t_2048), .c(t_2045), .d(t_7455), .cin(t_7458), .o(t_7470), .co(t_7471), .cout(t_7472));
compressor_4_2 u2_2571(.a(t_2060), .b(t_2057), .c(t_2054), .d(t_7461), .cin(t_7464), .o(t_7473), .co(t_7474), .cout(t_7475));
compressor_4_2 u2_2572(.a(t_2072), .b(t_2069), .c(t_2066), .d(t_2063), .cin(t_7466), .o(t_7476), .co(t_7477), .cout(t_7478));
compressor_4_2 u2_2573(.a(t_2011), .b(t_2008), .c(t_2005), .d(t_2002), .cin(t_2075), .o(t_7479), .co(t_7480), .cout(t_7481));
compressor_4_2 u2_2574(.a(t_2026), .b(t_2023), .c(t_2020), .d(t_2017), .cin(t_2014), .o(t_7482), .co(t_7483), .cout(t_7484));
compressor_3_2 u1_2575(.a(t_2035), .b(t_2032), .cin(t_2029), .o(t_7485), .cout(t_7486));
compressor_4_2 u2_2576(.a(t_2084), .b(t_2081), .c(t_2078), .d(t_7469), .cin(t_7472), .o(t_7487), .co(t_7488), .cout(t_7489));
compressor_4_2 u2_2577(.a(t_2093), .b(t_2090), .c(t_2087), .d(t_7475), .cin(t_7478), .o(t_7490), .co(t_7491), .cout(t_7492));
compressor_4_2 u2_2578(.a(t_2102), .b(t_2099), .c(t_2096), .d(t_7481), .cin(t_7484), .o(t_7493), .co(t_7494), .cout(t_7495));
compressor_4_2 u2_2579(.a(t_2114), .b(t_2111), .c(t_2108), .d(t_2105), .cin(t_7486), .o(t_7496), .co(t_7497), .cout(t_7498));
compressor_4_2 u2_2580(.a(t_2052), .b(t_2049), .c(t_2046), .d(t_2043), .cin(t_2040), .o(t_7499), .co(t_7500), .cout(t_7501));
compressor_4_2 u2_2581(.a(t_2067), .b(t_2064), .c(t_2061), .d(t_2058), .cin(t_2055), .o(t_7502), .co(t_7503), .cout(t_7504));
compressor_3_2 u1_2582(.a(t_2076), .b(t_2073), .cin(t_2070), .o(t_7505), .cout(t_7506));
compressor_4_2 u2_2583(.a(t_2123), .b(t_2120), .c(t_2117), .d(t_7489), .cin(t_7492), .o(t_7507), .co(t_7508), .cout(t_7509));
compressor_4_2 u2_2584(.a(t_2132), .b(t_2129), .c(t_2126), .d(t_7495), .cin(t_7498), .o(t_7510), .co(t_7511), .cout(t_7512));
compressor_4_2 u2_2585(.a(t_2141), .b(t_2138), .c(t_2135), .d(t_7501), .cin(t_7504), .o(t_7513), .co(t_7514), .cout(t_7515));
compressor_4_2 u2_2586(.a(t_2153), .b(t_2150), .c(t_2147), .d(t_2144), .cin(t_7506), .o(t_7516), .co(t_7517), .cout(t_7518));
compressor_4_2 u2_2587(.a(t_2088), .b(t_2085), .c(t_2082), .d(t_2079), .cin(t_2156), .o(t_7519), .co(t_7520), .cout(t_7521));
compressor_4_2 u2_2588(.a(t_2103), .b(t_2100), .c(t_2097), .d(t_2094), .cin(t_2091), .o(t_7522), .co(t_7523), .cout(t_7524));
compressor_3_2 u1_2589(.a(t_2112), .b(t_2109), .cin(t_2106), .o(t_7525), .cout(t_7526));
compressor_4_2 u2_2590(.a(t_2164), .b(t_2161), .c(t_2158), .d(t_7509), .cin(t_7512), .o(t_7527), .co(t_7528), .cout(t_7529));
compressor_4_2 u2_2591(.a(t_2173), .b(t_2170), .c(t_2167), .d(t_7515), .cin(t_7518), .o(t_7530), .co(t_7531), .cout(t_7532));
compressor_4_2 u2_2592(.a(t_2182), .b(t_2179), .c(t_2176), .d(t_7521), .cin(t_7524), .o(t_7533), .co(t_7534), .cout(t_7535));
compressor_4_2 u2_2593(.a(t_2194), .b(t_2191), .c(t_2188), .d(t_2185), .cin(t_7526), .o(t_7536), .co(t_7537), .cout(t_7538));
compressor_4_2 u2_2594(.a(t_2127), .b(t_2124), .c(t_2121), .d(t_2118), .cin(t_2197), .o(t_7539), .co(t_7540), .cout(t_7541));
compressor_4_2 u2_2595(.a(t_2142), .b(t_2139), .c(t_2136), .d(t_2133), .cin(t_2130), .o(t_7542), .co(t_7543), .cout(t_7544));
compressor_3_2 u1_2596(.a(t_2151), .b(t_2148), .cin(t_2145), .o(t_7545), .cout(t_7546));
compressor_4_2 u2_2597(.a(t_2202), .b(t_2199), .c(s_106_54), .d(t_7529), .cin(t_7532), .o(t_7547), .co(t_7548), .cout(t_7549));
compressor_4_2 u2_2598(.a(t_2211), .b(t_2208), .c(t_2205), .d(t_7535), .cin(t_7538), .o(t_7550), .co(t_7551), .cout(t_7552));
compressor_4_2 u2_2599(.a(t_2220), .b(t_2217), .c(t_2214), .d(t_7541), .cin(t_7544), .o(t_7553), .co(t_7554), .cout(t_7555));
compressor_4_2 u2_2600(.a(t_2232), .b(t_2229), .c(t_2226), .d(t_2223), .cin(t_7546), .o(t_7556), .co(t_7557), .cout(t_7558));
compressor_4_2 u2_2601(.a(t_2165), .b(t_2162), .c(t_2159), .d(t_2238), .cin(t_2235), .o(t_7559), .co(t_7560), .cout(t_7561));
compressor_4_2 u2_2602(.a(t_2180), .b(t_2177), .c(t_2174), .d(t_2171), .cin(t_2168), .o(t_7562), .co(t_7563), .cout(t_7564));
compressor_4_2 u2_2603(.a(t_2195), .b(t_2192), .c(t_2189), .d(t_2186), .cin(t_2183), .o(t_7565), .co(t_7566), .cout(t_7567));
compressor_4_2 u2_2604(.a(t_2246), .b(t_2243), .c(t_2240), .d(t_7549), .cin(t_7552), .o(t_7568), .co(t_7569), .cout(t_7570));
compressor_4_2 u2_2605(.a(t_2255), .b(t_2252), .c(t_2249), .d(t_7555), .cin(t_7558), .o(t_7571), .co(t_7572), .cout(t_7573));
compressor_4_2 u2_2606(.a(t_2264), .b(t_2261), .c(t_2258), .d(t_7561), .cin(t_7564), .o(t_7574), .co(t_7575), .cout(t_7576));
compressor_4_2 u2_2607(.a(t_2276), .b(t_2273), .c(t_2270), .d(t_2267), .cin(t_7567), .o(t_7577), .co(t_7578), .cout(t_7579));
compressor_4_2 u2_2608(.a(t_2209), .b(t_2206), .c(t_2203), .d(t_2200), .cin(t_2279), .o(t_7580), .co(t_7581), .cout(t_7582));
compressor_4_2 u2_2609(.a(t_2224), .b(t_2221), .c(t_2218), .d(t_2215), .cin(t_2212), .o(t_7583), .co(t_7584), .cout(t_7585));
compressor_3_2 u1_2610(.a(t_2233), .b(t_2230), .cin(t_2227), .o(t_7586), .cout(t_7587));
compressor_4_2 u2_2611(.a(t_2287), .b(t_2284), .c(t_2281), .d(t_7570), .cin(t_7573), .o(t_7588), .co(t_7589), .cout(t_7590));
compressor_4_2 u2_2612(.a(t_2296), .b(t_2293), .c(t_2290), .d(t_7576), .cin(t_7579), .o(t_7591), .co(t_7592), .cout(t_7593));
compressor_4_2 u2_2613(.a(t_2305), .b(t_2302), .c(t_2299), .d(t_7582), .cin(t_7585), .o(t_7594), .co(t_7595), .cout(t_7596));
compressor_4_2 u2_2614(.a(t_2317), .b(t_2314), .c(t_2311), .d(t_2308), .cin(t_7587), .o(t_7597), .co(t_7598), .cout(t_7599));
compressor_4_2 u2_2615(.a(t_2250), .b(t_2247), .c(t_2244), .d(t_2241), .cin(t_2320), .o(t_7600), .co(t_7601), .cout(t_7602));
compressor_4_2 u2_2616(.a(t_2265), .b(t_2262), .c(t_2259), .d(t_2256), .cin(t_2253), .o(t_7603), .co(t_7604), .cout(t_7605));
compressor_3_2 u1_2617(.a(t_2274), .b(t_2271), .cin(t_2268), .o(t_7606), .cout(t_7607));
compressor_4_2 u2_2618(.a(t_2326), .b(t_2323), .c(s_109_54), .d(t_7590), .cin(t_7593), .o(t_7608), .co(t_7609), .cout(t_7610));
compressor_4_2 u2_2619(.a(t_2335), .b(t_2332), .c(t_2329), .d(t_7596), .cin(t_7599), .o(t_7611), .co(t_7612), .cout(t_7613));
compressor_4_2 u2_2620(.a(t_2344), .b(t_2341), .c(t_2338), .d(t_7602), .cin(t_7605), .o(t_7614), .co(t_7615), .cout(t_7616));
compressor_4_2 u2_2621(.a(t_2356), .b(t_2353), .c(t_2350), .d(t_2347), .cin(t_7607), .o(t_7617), .co(t_7618), .cout(t_7619));
compressor_4_2 u2_2622(.a(t_2288), .b(t_2285), .c(t_2282), .d(t_2362), .cin(t_2359), .o(t_7620), .co(t_7621), .cout(t_7622));
compressor_4_2 u2_2623(.a(t_2303), .b(t_2300), .c(t_2297), .d(t_2294), .cin(t_2291), .o(t_7623), .co(t_7624), .cout(t_7625));
compressor_4_2 u2_2624(.a(t_2318), .b(t_2315), .c(t_2312), .d(t_2309), .cin(t_2306), .o(t_7626), .co(t_7627), .cout(t_7628));
compressor_4_2 u2_2625(.a(t_2367), .b(t_2364), .c(s_110_56), .d(t_7610), .cin(t_7613), .o(t_7629), .co(t_7630), .cout(t_7631));
compressor_4_2 u2_2626(.a(t_2376), .b(t_2373), .c(t_2370), .d(t_7616), .cin(t_7619), .o(t_7632), .co(t_7633), .cout(t_7634));
compressor_4_2 u2_2627(.a(t_2385), .b(t_2382), .c(t_2379), .d(t_7622), .cin(t_7625), .o(t_7635), .co(t_7636), .cout(t_7637));
compressor_4_2 u2_2628(.a(t_2397), .b(t_2394), .c(t_2391), .d(t_2388), .cin(t_7628), .o(t_7638), .co(t_7639), .cout(t_7640));
compressor_4_2 u2_2629(.a(t_2330), .b(t_2327), .c(t_2324), .d(t_2403), .cin(t_2400), .o(t_7641), .co(t_7642), .cout(t_7643));
compressor_4_2 u2_2630(.a(t_2345), .b(t_2342), .c(t_2339), .d(t_2336), .cin(t_2333), .o(t_7644), .co(t_7645), .cout(t_7646));
compressor_4_2 u2_2631(.a(t_2360), .b(t_2357), .c(t_2354), .d(t_2351), .cin(t_2348), .o(t_7647), .co(t_7648), .cout(t_7649));
compressor_4_2 u2_2632(.a(t_2412), .b(t_2409), .c(t_2406), .d(t_7631), .cin(t_7634), .o(t_7650), .co(t_7651), .cout(t_7652));
compressor_4_2 u2_2633(.a(t_2421), .b(t_2418), .c(t_2415), .d(t_7637), .cin(t_7640), .o(t_7653), .co(t_7654), .cout(t_7655));
compressor_4_2 u2_2634(.a(t_2430), .b(t_2427), .c(t_2424), .d(t_7643), .cin(t_7646), .o(t_7656), .co(t_7657), .cout(t_7658));
compressor_4_2 u2_2635(.a(t_2442), .b(t_2439), .c(t_2436), .d(t_2433), .cin(t_7649), .o(t_7659), .co(t_7660), .cout(t_7661));
compressor_4_2 u2_2636(.a(t_2374), .b(t_2371), .c(t_2368), .d(t_2365), .cin(t_2445), .o(t_7662), .co(t_7663), .cout(t_7664));
compressor_4_2 u2_2637(.a(t_2389), .b(t_2386), .c(t_2383), .d(t_2380), .cin(t_2377), .o(t_7665), .co(t_7666), .cout(t_7667));
compressor_4_2 u2_2638(.a(t_2404), .b(t_2401), .c(t_2398), .d(t_2395), .cin(t_2392), .o(t_7668), .co(t_7669), .cout(t_7670));
compressor_4_2 u2_2639(.a(t_2454), .b(t_2451), .c(t_2448), .d(t_7652), .cin(t_7655), .o(t_7671), .co(t_7672), .cout(t_7673));
compressor_4_2 u2_2640(.a(t_2463), .b(t_2460), .c(t_2457), .d(t_7658), .cin(t_7661), .o(t_7674), .co(t_7675), .cout(t_7676));
compressor_4_2 u2_2641(.a(t_2472), .b(t_2469), .c(t_2466), .d(t_7664), .cin(t_7667), .o(t_7677), .co(t_7678), .cout(t_7679));
compressor_4_2 u2_2642(.a(t_2484), .b(t_2481), .c(t_2478), .d(t_2475), .cin(t_7670), .o(t_7680), .co(t_7681), .cout(t_7682));
compressor_4_2 u2_2643(.a(t_2413), .b(t_2410), .c(t_2407), .d(t_2490), .cin(t_2487), .o(t_7683), .co(t_7684), .cout(t_7685));
compressor_4_2 u2_2644(.a(t_2428), .b(t_2425), .c(t_2422), .d(t_2419), .cin(t_2416), .o(t_7686), .co(t_7687), .cout(t_7688));
compressor_4_2 u2_2645(.a(t_2443), .b(t_2440), .c(t_2437), .d(t_2434), .cin(t_2431), .o(t_7689), .co(t_7690), .cout(t_7691));
compressor_4_2 u2_2646(.a(t_2498), .b(t_2495), .c(t_2492), .d(t_7673), .cin(t_7676), .o(t_7692), .co(t_7693), .cout(t_7694));
compressor_4_2 u2_2647(.a(t_2507), .b(t_2504), .c(t_2501), .d(t_7679), .cin(t_7682), .o(t_7695), .co(t_7696), .cout(t_7697));
compressor_4_2 u2_2648(.a(t_2516), .b(t_2513), .c(t_2510), .d(t_7685), .cin(t_7688), .o(t_7698), .co(t_7699), .cout(t_7700));
compressor_4_2 u2_2649(.a(t_2528), .b(t_2525), .c(t_2522), .d(t_2519), .cin(t_7691), .o(t_7701), .co(t_7702), .cout(t_7703));
compressor_4_2 u2_2650(.a(t_2455), .b(t_2452), .c(t_2449), .d(t_2534), .cin(t_2531), .o(t_7704), .co(t_7705), .cout(t_7706));
compressor_4_2 u2_2651(.a(t_2470), .b(t_2467), .c(t_2464), .d(t_2461), .cin(t_2458), .o(t_7707), .co(t_7708), .cout(t_7709));
compressor_4_2 u2_2652(.a(t_2485), .b(t_2482), .c(t_2479), .d(t_2476), .cin(t_2473), .o(t_7710), .co(t_7711), .cout(t_7712));
compressor_4_2 u2_2653(.a(t_2539), .b(t_2536), .c(s_114_58), .d(t_7694), .cin(t_7697), .o(t_7713), .co(t_7714), .cout(t_7715));
compressor_4_2 u2_2654(.a(t_2548), .b(t_2545), .c(t_2542), .d(t_7700), .cin(t_7703), .o(t_7716), .co(t_7717), .cout(t_7718));
compressor_4_2 u2_2655(.a(t_2557), .b(t_2554), .c(t_2551), .d(t_7706), .cin(t_7709), .o(t_7719), .co(t_7720), .cout(t_7721));
compressor_4_2 u2_2656(.a(t_2569), .b(t_2566), .c(t_2563), .d(t_2560), .cin(t_7712), .o(t_7722), .co(t_7723), .cout(t_7724));
compressor_4_2 u2_2657(.a(t_2496), .b(t_2493), .c(t_2578), .d(t_2575), .cin(t_2572), .o(t_7725), .co(t_7726), .cout(t_7727));
compressor_4_2 u2_2658(.a(t_2511), .b(t_2508), .c(t_2505), .d(t_2502), .cin(t_2499), .o(t_7728), .co(t_7729), .cout(t_7730));
compressor_4_2 u2_2659(.a(t_2526), .b(t_2523), .c(t_2520), .d(t_2517), .cin(t_2514), .o(t_7731), .co(t_7732), .cout(t_7733));
half_adder u0_2660(.a(t_2532), .b(t_2529), .o(t_7734), .cout(t_7735));
compressor_4_2 u2_2661(.a(t_2586), .b(t_2583), .c(t_2580), .d(t_7715), .cin(t_7718), .o(t_7736), .co(t_7737), .cout(t_7738));
compressor_4_2 u2_2662(.a(t_2595), .b(t_2592), .c(t_2589), .d(t_7721), .cin(t_7724), .o(t_7739), .co(t_7740), .cout(t_7741));
compressor_4_2 u2_2663(.a(t_2604), .b(t_2601), .c(t_2598), .d(t_7727), .cin(t_7730), .o(t_7742), .co(t_7743), .cout(t_7744));
compressor_4_2 u2_2664(.a(t_2613), .b(t_2610), .c(t_2607), .d(t_7733), .cin(t_7735), .o(t_7745), .co(t_7746), .cout(t_7747));
compressor_4_2 u2_2665(.a(t_2540), .b(t_2537), .c(t_2622), .d(t_2619), .cin(t_2616), .o(t_7748), .co(t_7749), .cout(t_7750));
compressor_4_2 u2_2666(.a(t_2555), .b(t_2552), .c(t_2549), .d(t_2546), .cin(t_2543), .o(t_7751), .co(t_7752), .cout(t_7753));
compressor_4_2 u2_2667(.a(t_2570), .b(t_2567), .c(t_2564), .d(t_2561), .cin(t_2558), .o(t_7754), .co(t_7755), .cout(t_7756));
half_adder u0_2668(.a(t_2576), .b(t_2573), .o(t_7757), .cout(t_7758));
compressor_4_2 u2_2669(.a(t_2630), .b(t_2627), .c(t_2624), .d(t_7738), .cin(t_7741), .o(t_7759), .co(t_7760), .cout(t_7761));
compressor_4_2 u2_2670(.a(t_2639), .b(t_2636), .c(t_2633), .d(t_7744), .cin(t_7747), .o(t_7762), .co(t_7763), .cout(t_7764));
compressor_4_2 u2_2671(.a(t_2648), .b(t_2645), .c(t_2642), .d(t_7750), .cin(t_7753), .o(t_7765), .co(t_7766), .cout(t_7767));
compressor_4_2 u2_2672(.a(t_2657), .b(t_2654), .c(t_2651), .d(t_7756), .cin(t_7758), .o(t_7768), .co(t_7769), .cout(t_7770));
compressor_4_2 u2_2673(.a(t_2584), .b(t_2581), .c(t_2666), .d(t_2663), .cin(t_2660), .o(t_7771), .co(t_7772), .cout(t_7773));
compressor_4_2 u2_2674(.a(t_2599), .b(t_2596), .c(t_2593), .d(t_2590), .cin(t_2587), .o(t_7774), .co(t_7775), .cout(t_7776));
compressor_4_2 u2_2675(.a(t_2614), .b(t_2611), .c(t_2608), .d(t_2605), .cin(t_2602), .o(t_7777), .co(t_7778), .cout(t_7779));
half_adder u0_2676(.a(t_2620), .b(t_2617), .o(t_7780), .cout(t_7781));
compressor_4_2 u2_2677(.a(t_2672), .b(t_2669), .c(s_117_58), .d(t_7761), .cin(t_7764), .o(t_7782), .co(t_7783), .cout(t_7784));
compressor_4_2 u2_2678(.a(t_2681), .b(t_2678), .c(t_2675), .d(t_7767), .cin(t_7770), .o(t_7785), .co(t_7786), .cout(t_7787));
compressor_4_2 u2_2679(.a(t_2690), .b(t_2687), .c(t_2684), .d(t_7773), .cin(t_7776), .o(t_7788), .co(t_7789), .cout(t_7790));
compressor_4_2 u2_2680(.a(t_2699), .b(t_2696), .c(t_2693), .d(t_7779), .cin(t_7781), .o(t_7791), .co(t_7792), .cout(t_7793));
compressor_4_2 u2_2681(.a(t_2625), .b(t_2711), .c(t_2708), .d(t_2705), .cin(t_2702), .o(t_7794), .co(t_7795), .cout(t_7796));
compressor_4_2 u2_2682(.a(t_2640), .b(t_2637), .c(t_2634), .d(t_2631), .cin(t_2628), .o(t_7797), .co(t_7798), .cout(t_7799));
compressor_4_2 u2_2683(.a(t_2655), .b(t_2652), .c(t_2649), .d(t_2646), .cin(t_2643), .o(t_7800), .co(t_7801), .cout(t_7802));
compressor_3_2 u1_2684(.a(t_2664), .b(t_2661), .cin(t_2658), .o(t_7803), .cout(t_7804));
compressor_4_2 u2_2685(.a(t_2716), .b(t_2713), .c(s_118_60), .d(t_7784), .cin(t_7787), .o(t_7805), .co(t_7806), .cout(t_7807));
compressor_4_2 u2_2686(.a(t_2725), .b(t_2722), .c(t_2719), .d(t_7790), .cin(t_7793), .o(t_7808), .co(t_7809), .cout(t_7810));
compressor_4_2 u2_2687(.a(t_2734), .b(t_2731), .c(t_2728), .d(t_7796), .cin(t_7799), .o(t_7811), .co(t_7812), .cout(t_7813));
compressor_4_2 u2_2688(.a(t_2743), .b(t_2740), .c(t_2737), .d(t_7802), .cin(t_7804), .o(t_7814), .co(t_7815), .cout(t_7816));
compressor_4_2 u2_2689(.a(t_2670), .b(t_2755), .c(t_2752), .d(t_2749), .cin(t_2746), .o(t_7817), .co(t_7818), .cout(t_7819));
compressor_4_2 u2_2690(.a(t_2685), .b(t_2682), .c(t_2679), .d(t_2676), .cin(t_2673), .o(t_7820), .co(t_7821), .cout(t_7822));
compressor_4_2 u2_2691(.a(t_2700), .b(t_2697), .c(t_2694), .d(t_2691), .cin(t_2688), .o(t_7823), .co(t_7824), .cout(t_7825));
compressor_3_2 u1_2692(.a(t_2709), .b(t_2706), .cin(t_2703), .o(t_7826), .cout(t_7827));
compressor_4_2 u2_2693(.a(t_2764), .b(t_2761), .c(t_2758), .d(t_7807), .cin(t_7810), .o(t_7828), .co(t_7829), .cout(t_7830));
compressor_4_2 u2_2694(.a(t_2773), .b(t_2770), .c(t_2767), .d(t_7813), .cin(t_7816), .o(t_7831), .co(t_7832), .cout(t_7833));
compressor_4_2 u2_2695(.a(t_2782), .b(t_2779), .c(t_2776), .d(t_7819), .cin(t_7822), .o(t_7834), .co(t_7835), .cout(t_7836));
compressor_4_2 u2_2696(.a(t_2791), .b(t_2788), .c(t_2785), .d(t_7825), .cin(t_7827), .o(t_7837), .co(t_7838), .cout(t_7839));
compressor_4_2 u2_2697(.a(t_2717), .b(t_2714), .c(t_2800), .d(t_2797), .cin(t_2794), .o(t_7840), .co(t_7841), .cout(t_7842));
compressor_4_2 u2_2698(.a(t_2732), .b(t_2729), .c(t_2726), .d(t_2723), .cin(t_2720), .o(t_7843), .co(t_7844), .cout(t_7845));
compressor_4_2 u2_2699(.a(t_2747), .b(t_2744), .c(t_2741), .d(t_2738), .cin(t_2735), .o(t_7846), .co(t_7847), .cout(t_7848));
compressor_3_2 u1_2700(.a(t_2756), .b(t_2753), .cin(t_2750), .o(t_7849), .cout(t_7850));
compressor_4_2 u2_2701(.a(t_2809), .b(t_2806), .c(t_2803), .d(t_7830), .cin(t_7833), .o(t_7851), .co(t_7852), .cout(t_7853));
compressor_4_2 u2_2702(.a(t_2818), .b(t_2815), .c(t_2812), .d(t_7836), .cin(t_7839), .o(t_7854), .co(t_7855), .cout(t_7856));
compressor_4_2 u2_2703(.a(t_2827), .b(t_2824), .c(t_2821), .d(t_7842), .cin(t_7845), .o(t_7857), .co(t_7858), .cout(t_7859));
compressor_4_2 u2_2704(.a(t_2836), .b(t_2833), .c(t_2830), .d(t_7848), .cin(t_7850), .o(t_7860), .co(t_7861), .cout(t_7862));
compressor_4_2 u2_2705(.a(t_2759), .b(t_2848), .c(t_2845), .d(t_2842), .cin(t_2839), .o(t_7863), .co(t_7864), .cout(t_7865));
compressor_4_2 u2_2706(.a(t_2774), .b(t_2771), .c(t_2768), .d(t_2765), .cin(t_2762), .o(t_7866), .co(t_7867), .cout(t_7868));
compressor_4_2 u2_2707(.a(t_2789), .b(t_2786), .c(t_2783), .d(t_2780), .cin(t_2777), .o(t_7869), .co(t_7870), .cout(t_7871));
compressor_3_2 u1_2708(.a(t_2798), .b(t_2795), .cin(t_2792), .o(t_7872), .cout(t_7873));
compressor_4_2 u2_2709(.a(t_2856), .b(t_2853), .c(t_2850), .d(t_7853), .cin(t_7856), .o(t_7874), .co(t_7875), .cout(t_7876));
compressor_4_2 u2_2710(.a(t_2865), .b(t_2862), .c(t_2859), .d(t_7859), .cin(t_7862), .o(t_7877), .co(t_7878), .cout(t_7879));
compressor_4_2 u2_2711(.a(t_2874), .b(t_2871), .c(t_2868), .d(t_7865), .cin(t_7868), .o(t_7880), .co(t_7881), .cout(t_7882));
compressor_4_2 u2_2712(.a(t_2883), .b(t_2880), .c(t_2877), .d(t_7871), .cin(t_7873), .o(t_7883), .co(t_7884), .cout(t_7885));
compressor_4_2 u2_2713(.a(t_2804), .b(t_2895), .c(t_2892), .d(t_2889), .cin(t_2886), .o(t_7886), .co(t_7887), .cout(t_7888));
compressor_4_2 u2_2714(.a(t_2819), .b(t_2816), .c(t_2813), .d(t_2810), .cin(t_2807), .o(t_7889), .co(t_7890), .cout(t_7891));
compressor_4_2 u2_2715(.a(t_2834), .b(t_2831), .c(t_2828), .d(t_2825), .cin(t_2822), .o(t_7892), .co(t_7893), .cout(t_7894));
compressor_3_2 u1_2716(.a(t_2843), .b(t_2840), .cin(t_2837), .o(t_7895), .cout(t_7896));
compressor_4_2 u2_2717(.a(t_2900), .b(t_2897), .c(s_122_62), .d(t_7876), .cin(t_7879), .o(t_7897), .co(t_7898), .cout(t_7899));
compressor_4_2 u2_2718(.a(t_2909), .b(t_2906), .c(t_2903), .d(t_7882), .cin(t_7885), .o(t_7900), .co(t_7901), .cout(t_7902));
compressor_4_2 u2_2719(.a(t_2918), .b(t_2915), .c(t_2912), .d(t_7888), .cin(t_7891), .o(t_7903), .co(t_7904), .cout(t_7905));
compressor_4_2 u2_2720(.a(t_2927), .b(t_2924), .c(t_2921), .d(t_7894), .cin(t_7896), .o(t_7906), .co(t_7907), .cout(t_7908));
compressor_4_2 u2_2721(.a(t_2942), .b(t_2939), .c(t_2936), .d(t_2933), .cin(t_2930), .o(t_7909), .co(t_7910), .cout(t_7911));
compressor_4_2 u2_2722(.a(t_2863), .b(t_2860), .c(t_2857), .d(t_2854), .cin(t_2851), .o(t_7912), .co(t_7913), .cout(t_7914));
compressor_4_2 u2_2723(.a(t_2878), .b(t_2875), .c(t_2872), .d(t_2869), .cin(t_2866), .o(t_7915), .co(t_7916), .cout(t_7917));
compressor_4_2 u2_2724(.a(t_2893), .b(t_2890), .c(t_2887), .d(t_2884), .cin(t_2881), .o(t_7918), .co(t_7919), .cout(t_7920));
compressor_4_2 u2_2725(.a(t_2950), .b(t_2947), .c(t_2944), .d(t_7899), .cin(t_7902), .o(t_7921), .co(t_7922), .cout(t_7923));
compressor_4_2 u2_2726(.a(t_2959), .b(t_2956), .c(t_2953), .d(t_7905), .cin(t_7908), .o(t_7924), .co(t_7925), .cout(t_7926));
compressor_4_2 u2_2727(.a(t_2968), .b(t_2965), .c(t_2962), .d(t_7911), .cin(t_7914), .o(t_7927), .co(t_7928), .cout(t_7929));
compressor_4_2 u2_2728(.a(t_2977), .b(t_2974), .c(t_2971), .d(t_7917), .cin(t_7920), .o(t_7930), .co(t_7931), .cout(t_7932));
compressor_4_2 u2_2729(.a(t_2898), .b(t_2989), .c(t_2986), .d(t_2983), .cin(t_2980), .o(t_7933), .co(t_7934), .cout(t_7935));
compressor_4_2 u2_2730(.a(t_2913), .b(t_2910), .c(t_2907), .d(t_2904), .cin(t_2901), .o(t_7936), .co(t_7937), .cout(t_7938));
compressor_4_2 u2_2731(.a(t_2928), .b(t_2925), .c(t_2922), .d(t_2919), .cin(t_2916), .o(t_7939), .co(t_7940), .cout(t_7941));
compressor_3_2 u1_2732(.a(t_2937), .b(t_2934), .cin(t_2931), .o(t_7942), .cout(t_7943));
compressor_4_2 u2_2733(.a(t_2997), .b(t_2994), .c(t_2991), .d(t_7923), .cin(t_7926), .o(t_7944), .co(t_7945), .cout(t_7946));
compressor_4_2 u2_2734(.a(t_3006), .b(t_3003), .c(t_3000), .d(t_7929), .cin(t_7932), .o(t_7947), .co(t_7948), .cout(t_7949));
compressor_4_2 u2_2735(.a(t_3015), .b(t_3012), .c(t_3009), .d(t_7935), .cin(t_7938), .o(t_7950), .co(t_7951), .cout(t_7952));
compressor_4_2 u2_2736(.a(t_3024), .b(t_3021), .c(t_3018), .d(t_7941), .cin(t_7943), .o(t_7953), .co(t_7954), .cout(t_7955));
compressor_4_2 u2_2737(.a(t_2945), .b(t_3036), .c(t_3033), .d(t_3030), .cin(t_3027), .o(t_7956), .co(t_7957), .cout(t_7958));
compressor_4_2 u2_2738(.a(t_2960), .b(t_2957), .c(t_2954), .d(t_2951), .cin(t_2948), .o(t_7959), .co(t_7960), .cout(t_7961));
compressor_4_2 u2_2739(.a(t_2975), .b(t_2972), .c(t_2969), .d(t_2966), .cin(t_2963), .o(t_7962), .co(t_7963), .cout(t_7964));
compressor_3_2 u1_2740(.a(t_2984), .b(t_2981), .cin(t_2978), .o(t_7965), .cout(t_7966));
compressor_4_2 u2_2741(.a(t_3042), .b(t_3039), .c(s_125_62), .d(t_7946), .cin(t_7949), .o(t_7967), .co(t_7968), .cout(t_7969));
compressor_4_2 u2_2742(.a(t_3051), .b(t_3048), .c(t_3045), .d(t_7952), .cin(t_7955), .o(t_7970), .co(t_7971), .cout(t_7972));
compressor_4_2 u2_2743(.a(t_3060), .b(t_3057), .c(t_3054), .d(t_7958), .cin(t_7961), .o(t_7973), .co(t_7974), .cout(t_7975));
compressor_4_2 u2_2744(.a(t_3069), .b(t_3066), .c(t_3063), .d(t_7964), .cin(t_7966), .o(t_7976), .co(t_7977), .cout(t_7978));
compressor_4_2 u2_2745(.a(t_3084), .b(t_3081), .c(t_3078), .d(t_3075), .cin(t_3072), .o(t_7979), .co(t_7980), .cout(t_7981));
compressor_4_2 u2_2746(.a(t_3004), .b(t_3001), .c(t_2998), .d(t_2995), .cin(t_2992), .o(t_7982), .co(t_7983), .cout(t_7984));
compressor_4_2 u2_2747(.a(t_3019), .b(t_3016), .c(t_3013), .d(t_3010), .cin(t_3007), .o(t_7985), .co(t_7986), .cout(t_7987));
compressor_4_2 u2_2748(.a(t_3034), .b(t_3031), .c(t_3028), .d(t_3025), .cin(t_3022), .o(t_7988), .co(t_7989), .cout(t_7990));
compressor_4_2 u2_2749(.a(t_3089), .b(t_3086), .c(s_126_64), .d(t_7969), .cin(t_7972), .o(t_7991), .co(t_7992), .cout(t_7993));
compressor_4_2 u2_2750(.a(t_3098), .b(t_3095), .c(t_3092), .d(t_7975), .cin(t_7978), .o(t_7994), .co(t_7995), .cout(t_7996));
compressor_4_2 u2_2751(.a(t_3107), .b(t_3104), .c(t_3101), .d(t_7981), .cin(t_7984), .o(t_7997), .co(t_7998), .cout(t_7999));
compressor_4_2 u2_2752(.a(t_3116), .b(t_3113), .c(t_3110), .d(t_7987), .cin(t_7990), .o(t_8000), .co(t_8001), .cout(t_8002));
compressor_4_2 u2_2753(.a(t_3131), .b(t_3128), .c(t_3125), .d(t_3122), .cin(t_3119), .o(t_8003), .co(t_8004), .cout(t_8005));
compressor_4_2 u2_2754(.a(t_3052), .b(t_3049), .c(t_3046), .d(t_3043), .cin(t_3040), .o(t_8006), .co(t_8007), .cout(t_8008));
compressor_4_2 u2_2755(.a(t_3067), .b(t_3064), .c(t_3061), .d(t_3058), .cin(t_3055), .o(t_8009), .co(t_8010), .cout(t_8011));
compressor_4_2 u2_2756(.a(t_3082), .b(t_3079), .c(t_3076), .d(t_3073), .cin(t_3070), .o(t_8012), .co(t_8013), .cout(t_8014));
compressor_4_2 u2_2757(.a(t_3140), .b(t_3137), .c(t_3134), .d(t_7993), .cin(t_7996), .o(t_8015), .co(t_8016), .cout(t_8017));
compressor_4_2 u2_2758(.a(t_3149), .b(t_3146), .c(t_3143), .d(t_7999), .cin(t_8002), .o(t_8018), .co(t_8019), .cout(t_8020));
compressor_4_2 u2_2759(.a(t_3158), .b(t_3155), .c(t_3152), .d(t_8005), .cin(t_8008), .o(t_8021), .co(t_8022), .cout(t_8023));
compressor_4_2 u2_2760(.a(t_3167), .b(t_3164), .c(t_3161), .d(t_8011), .cin(t_8014), .o(t_8024), .co(t_8025), .cout(t_8026));
compressor_4_2 u2_2761(.a(t_3087), .b(t_3179), .c(t_3176), .d(t_3173), .cin(t_3170), .o(t_8027), .co(t_8028), .cout(t_8029));
compressor_4_2 u2_2762(.a(t_3102), .b(t_3099), .c(t_3096), .d(t_3093), .cin(t_3090), .o(t_8030), .co(t_8031), .cout(t_8032));
compressor_4_2 u2_2763(.a(t_3117), .b(t_3114), .c(t_3111), .d(t_3108), .cin(t_3105), .o(t_8033), .co(t_8034), .cout(t_8035));
compressor_4_2 u2_2764(.a(t_3132), .b(t_3129), .c(t_3126), .d(t_3123), .cin(t_3120), .o(t_8036), .co(t_8037), .cout(t_8038));
compressor_4_2 u2_2765(.a(t_3185), .b(t_3182), .c(s_128_64), .d(t_8017), .cin(t_8020), .o(t_8039), .co(t_8040), .cout(t_8041));
compressor_4_2 u2_2766(.a(t_3194), .b(t_3191), .c(t_3188), .d(t_8023), .cin(t_8026), .o(t_8042), .co(t_8043), .cout(t_8044));
compressor_4_2 u2_2767(.a(t_3203), .b(t_3200), .c(t_3197), .d(t_8029), .cin(t_8032), .o(t_8045), .co(t_8046), .cout(t_8047));
compressor_4_2 u2_2768(.a(t_3212), .b(t_3209), .c(t_3206), .d(t_8035), .cin(t_8038), .o(t_8048), .co(t_8049), .cout(t_8050));
compressor_4_2 u2_2769(.a(t_3227), .b(t_3224), .c(t_3221), .d(t_3218), .cin(t_3215), .o(t_8051), .co(t_8052), .cout(t_8053));
compressor_4_2 u2_2770(.a(t_3147), .b(t_3144), .c(t_3141), .d(t_3138), .cin(t_3135), .o(t_8054), .co(t_8055), .cout(t_8056));
compressor_4_2 u2_2771(.a(t_3162), .b(t_3159), .c(t_3156), .d(t_3153), .cin(t_3150), .o(t_8057), .co(t_8058), .cout(t_8059));
compressor_4_2 u2_2772(.a(t_3177), .b(t_3174), .c(t_3171), .d(t_3168), .cin(t_3165), .o(t_8060), .co(t_8061), .cout(t_8062));
compressor_4_2 u2_2773(.a(t_3233), .b(t_3230), .c(s_129_64), .d(t_8041), .cin(t_8044), .o(t_8063), .co(t_8064), .cout(t_8065));
compressor_4_2 u2_2774(.a(t_3242), .b(t_3239), .c(t_3236), .d(t_8047), .cin(t_8050), .o(t_8066), .co(t_8067), .cout(t_8068));
compressor_4_2 u2_2775(.a(t_3251), .b(t_3248), .c(t_3245), .d(t_8053), .cin(t_8056), .o(t_8069), .co(t_8070), .cout(t_8071));
compressor_4_2 u2_2776(.a(t_3260), .b(t_3257), .c(t_3254), .d(t_8059), .cin(t_8062), .o(t_8072), .co(t_8073), .cout(t_8074));
compressor_4_2 u2_2777(.a(t_3275), .b(t_3272), .c(t_3269), .d(t_3266), .cin(t_3263), .o(t_8075), .co(t_8076), .cout(t_8077));
compressor_4_2 u2_2778(.a(t_3195), .b(t_3192), .c(t_3189), .d(t_3186), .cin(t_3183), .o(t_8078), .co(t_8079), .cout(t_8080));
compressor_4_2 u2_2779(.a(t_3210), .b(t_3207), .c(t_3204), .d(t_3201), .cin(t_3198), .o(t_8081), .co(t_8082), .cout(t_8083));
compressor_4_2 u2_2780(.a(t_3225), .b(t_3222), .c(t_3219), .d(t_3216), .cin(t_3213), .o(t_8084), .co(t_8085), .cout(t_8086));
compressor_4_2 u2_2781(.a(t_3284), .b(t_3281), .c(t_3278), .d(t_8065), .cin(t_8068), .o(t_8087), .co(t_8088), .cout(t_8089));
compressor_4_2 u2_2782(.a(t_3293), .b(t_3290), .c(t_3287), .d(t_8071), .cin(t_8074), .o(t_8090), .co(t_8091), .cout(t_8092));
compressor_4_2 u2_2783(.a(t_3302), .b(t_3299), .c(t_3296), .d(t_8077), .cin(t_8080), .o(t_8093), .co(t_8094), .cout(t_8095));
compressor_4_2 u2_2784(.a(t_3311), .b(t_3308), .c(t_3305), .d(t_8083), .cin(t_8086), .o(t_8096), .co(t_8097), .cout(t_8098));
compressor_4_2 u2_2785(.a(t_3231), .b(t_3323), .c(t_3320), .d(t_3317), .cin(t_3314), .o(t_8099), .co(t_8100), .cout(t_8101));
compressor_4_2 u2_2786(.a(t_3246), .b(t_3243), .c(t_3240), .d(t_3237), .cin(t_3234), .o(t_8102), .co(t_8103), .cout(t_8104));
compressor_4_2 u2_2787(.a(t_3261), .b(t_3258), .c(t_3255), .d(t_3252), .cin(t_3249), .o(t_8105), .co(t_8106), .cout(t_8107));
compressor_4_2 u2_2788(.a(t_3276), .b(t_3273), .c(t_3270), .d(t_3267), .cin(t_3264), .o(t_8108), .co(t_8109), .cout(t_8110));
compressor_4_2 u2_2789(.a(t_3332), .b(t_3329), .c(t_3326), .d(t_8089), .cin(t_8092), .o(t_8111), .co(t_8112), .cout(t_8113));
compressor_4_2 u2_2790(.a(t_3341), .b(t_3338), .c(t_3335), .d(t_8095), .cin(t_8098), .o(t_8114), .co(t_8115), .cout(t_8116));
compressor_4_2 u2_2791(.a(t_3350), .b(t_3347), .c(t_3344), .d(t_8101), .cin(t_8104), .o(t_8117), .co(t_8118), .cout(t_8119));
compressor_4_2 u2_2792(.a(t_3359), .b(t_3356), .c(t_3353), .d(t_8107), .cin(t_8110), .o(t_8120), .co(t_8121), .cout(t_8122));
compressor_4_2 u2_2793(.a(t_3279), .b(t_3371), .c(t_3368), .d(t_3365), .cin(t_3362), .o(t_8123), .co(t_8124), .cout(t_8125));
compressor_4_2 u2_2794(.a(t_3294), .b(t_3291), .c(t_3288), .d(t_3285), .cin(t_3282), .o(t_8126), .co(t_8127), .cout(t_8128));
compressor_4_2 u2_2795(.a(t_3309), .b(t_3306), .c(t_3303), .d(t_3300), .cin(t_3297), .o(t_8129), .co(t_8130), .cout(t_8131));
compressor_4_2 u2_2796(.a(t_3324), .b(t_3321), .c(t_3318), .d(t_3315), .cin(t_3312), .o(t_8132), .co(t_8133), .cout(t_8134));
compressor_4_2 u2_2797(.a(t_3377), .b(t_3374), .c(s_132_62), .d(t_8113), .cin(t_8116), .o(t_8135), .co(t_8136), .cout(t_8137));
compressor_4_2 u2_2798(.a(t_3386), .b(t_3383), .c(t_3380), .d(t_8119), .cin(t_8122), .o(t_8138), .co(t_8139), .cout(t_8140));
compressor_4_2 u2_2799(.a(t_3395), .b(t_3392), .c(t_3389), .d(t_8125), .cin(t_8128), .o(t_8141), .co(t_8142), .cout(t_8143));
compressor_4_2 u2_2800(.a(t_3404), .b(t_3401), .c(t_3398), .d(t_8131), .cin(t_8134), .o(t_8144), .co(t_8145), .cout(t_8146));
compressor_4_2 u2_2801(.a(t_3419), .b(t_3416), .c(t_3413), .d(t_3410), .cin(t_3407), .o(t_8147), .co(t_8148), .cout(t_8149));
compressor_4_2 u2_2802(.a(t_3339), .b(t_3336), .c(t_3333), .d(t_3330), .cin(t_3327), .o(t_8150), .co(t_8151), .cout(t_8152));
compressor_4_2 u2_2803(.a(t_3354), .b(t_3351), .c(t_3348), .d(t_3345), .cin(t_3342), .o(t_8153), .co(t_8154), .cout(t_8155));
compressor_4_2 u2_2804(.a(t_3369), .b(t_3366), .c(t_3363), .d(t_3360), .cin(t_3357), .o(t_8156), .co(t_8157), .cout(t_8158));
compressor_4_2 u2_2805(.a(t_3424), .b(t_3421), .c(s_133_62), .d(t_8137), .cin(t_8140), .o(t_8159), .co(t_8160), .cout(t_8161));
compressor_4_2 u2_2806(.a(t_3433), .b(t_3430), .c(t_3427), .d(t_8143), .cin(t_8146), .o(t_8162), .co(t_8163), .cout(t_8164));
compressor_4_2 u2_2807(.a(t_3442), .b(t_3439), .c(t_3436), .d(t_8149), .cin(t_8152), .o(t_8165), .co(t_8166), .cout(t_8167));
compressor_4_2 u2_2808(.a(t_3451), .b(t_3448), .c(t_3445), .d(t_8155), .cin(t_8158), .o(t_8168), .co(t_8169), .cout(t_8170));
compressor_4_2 u2_2809(.a(t_3466), .b(t_3463), .c(t_3460), .d(t_3457), .cin(t_3454), .o(t_8171), .co(t_8172), .cout(t_8173));
compressor_4_2 u2_2810(.a(t_3387), .b(t_3384), .c(t_3381), .d(t_3378), .cin(t_3375), .o(t_8174), .co(t_8175), .cout(t_8176));
compressor_4_2 u2_2811(.a(t_3402), .b(t_3399), .c(t_3396), .d(t_3393), .cin(t_3390), .o(t_8177), .co(t_8178), .cout(t_8179));
compressor_4_2 u2_2812(.a(t_3417), .b(t_3414), .c(t_3411), .d(t_3408), .cin(t_3405), .o(t_8180), .co(t_8181), .cout(t_8182));
compressor_4_2 u2_2813(.a(t_3474), .b(t_3471), .c(t_3468), .d(t_8161), .cin(t_8164), .o(t_8183), .co(t_8184), .cout(t_8185));
compressor_4_2 u2_2814(.a(t_3483), .b(t_3480), .c(t_3477), .d(t_8167), .cin(t_8170), .o(t_8186), .co(t_8187), .cout(t_8188));
compressor_4_2 u2_2815(.a(t_3492), .b(t_3489), .c(t_3486), .d(t_8173), .cin(t_8176), .o(t_8189), .co(t_8190), .cout(t_8191));
compressor_4_2 u2_2816(.a(t_3501), .b(t_3498), .c(t_3495), .d(t_8179), .cin(t_8182), .o(t_8192), .co(t_8193), .cout(t_8194));
compressor_4_2 u2_2817(.a(t_3422), .b(t_3513), .c(t_3510), .d(t_3507), .cin(t_3504), .o(t_8195), .co(t_8196), .cout(t_8197));
compressor_4_2 u2_2818(.a(t_3437), .b(t_3434), .c(t_3431), .d(t_3428), .cin(t_3425), .o(t_8198), .co(t_8199), .cout(t_8200));
compressor_4_2 u2_2819(.a(t_3452), .b(t_3449), .c(t_3446), .d(t_3443), .cin(t_3440), .o(t_8201), .co(t_8202), .cout(t_8203));
compressor_3_2 u1_2820(.a(t_3461), .b(t_3458), .cin(t_3455), .o(t_8204), .cout(t_8205));
compressor_4_2 u2_2821(.a(t_3521), .b(t_3518), .c(t_3515), .d(t_8185), .cin(t_8188), .o(t_8206), .co(t_8207), .cout(t_8208));
compressor_4_2 u2_2822(.a(t_3530), .b(t_3527), .c(t_3524), .d(t_8191), .cin(t_8194), .o(t_8209), .co(t_8210), .cout(t_8211));
compressor_4_2 u2_2823(.a(t_3539), .b(t_3536), .c(t_3533), .d(t_8197), .cin(t_8200), .o(t_8212), .co(t_8213), .cout(t_8214));
compressor_4_2 u2_2824(.a(t_3548), .b(t_3545), .c(t_3542), .d(t_8203), .cin(t_8205), .o(t_8215), .co(t_8216), .cout(t_8217));
compressor_4_2 u2_2825(.a(t_3469), .b(t_3560), .c(t_3557), .d(t_3554), .cin(t_3551), .o(t_8218), .co(t_8219), .cout(t_8220));
compressor_4_2 u2_2826(.a(t_3484), .b(t_3481), .c(t_3478), .d(t_3475), .cin(t_3472), .o(t_8221), .co(t_8222), .cout(t_8223));
compressor_4_2 u2_2827(.a(t_3499), .b(t_3496), .c(t_3493), .d(t_3490), .cin(t_3487), .o(t_8224), .co(t_8225), .cout(t_8226));
compressor_3_2 u1_2828(.a(t_3508), .b(t_3505), .cin(t_3502), .o(t_8227), .cout(t_8228));
compressor_4_2 u2_2829(.a(t_3568), .b(t_3565), .c(t_3562), .d(t_8208), .cin(t_8211), .o(t_8229), .co(t_8230), .cout(t_8231));
compressor_4_2 u2_2830(.a(t_3577), .b(t_3574), .c(t_3571), .d(t_8214), .cin(t_8217), .o(t_8232), .co(t_8233), .cout(t_8234));
compressor_4_2 u2_2831(.a(t_3586), .b(t_3583), .c(t_3580), .d(t_8220), .cin(t_8223), .o(t_8235), .co(t_8236), .cout(t_8237));
compressor_4_2 u2_2832(.a(t_3595), .b(t_3592), .c(t_3589), .d(t_8226), .cin(t_8228), .o(t_8238), .co(t_8239), .cout(t_8240));
compressor_4_2 u2_2833(.a(t_3516), .b(t_3607), .c(t_3604), .d(t_3601), .cin(t_3598), .o(t_8241), .co(t_8242), .cout(t_8243));
compressor_4_2 u2_2834(.a(t_3531), .b(t_3528), .c(t_3525), .d(t_3522), .cin(t_3519), .o(t_8244), .co(t_8245), .cout(t_8246));
compressor_4_2 u2_2835(.a(t_3546), .b(t_3543), .c(t_3540), .d(t_3537), .cin(t_3534), .o(t_8247), .co(t_8248), .cout(t_8249));
compressor_3_2 u1_2836(.a(t_3555), .b(t_3552), .cin(t_3549), .o(t_8250), .cout(t_8251));
compressor_4_2 u2_2837(.a(t_3615), .b(t_3612), .c(t_3609), .d(t_8231), .cin(t_8234), .o(t_8252), .co(t_8253), .cout(t_8254));
compressor_4_2 u2_2838(.a(t_3624), .b(t_3621), .c(t_3618), .d(t_8237), .cin(t_8240), .o(t_8255), .co(t_8256), .cout(t_8257));
compressor_4_2 u2_2839(.a(t_3633), .b(t_3630), .c(t_3627), .d(t_8243), .cin(t_8246), .o(t_8258), .co(t_8259), .cout(t_8260));
compressor_4_2 u2_2840(.a(t_3642), .b(t_3639), .c(t_3636), .d(t_8249), .cin(t_8251), .o(t_8261), .co(t_8262), .cout(t_8263));
compressor_4_2 u2_2841(.a(t_3563), .b(t_3654), .c(t_3651), .d(t_3648), .cin(t_3645), .o(t_8264), .co(t_8265), .cout(t_8266));
compressor_4_2 u2_2842(.a(t_3578), .b(t_3575), .c(t_3572), .d(t_3569), .cin(t_3566), .o(t_8267), .co(t_8268), .cout(t_8269));
compressor_4_2 u2_2843(.a(t_3593), .b(t_3590), .c(t_3587), .d(t_3584), .cin(t_3581), .o(t_8270), .co(t_8271), .cout(t_8272));
compressor_3_2 u1_2844(.a(t_3602), .b(t_3599), .cin(t_3596), .o(t_8273), .cout(t_8274));
compressor_4_2 u2_2845(.a(t_3659), .b(t_3656), .c(s_138_59), .d(t_8254), .cin(t_8257), .o(t_8275), .co(t_8276), .cout(t_8277));
compressor_4_2 u2_2846(.a(t_3668), .b(t_3665), .c(t_3662), .d(t_8260), .cin(t_8263), .o(t_8278), .co(t_8279), .cout(t_8280));
compressor_4_2 u2_2847(.a(t_3677), .b(t_3674), .c(t_3671), .d(t_8266), .cin(t_8269), .o(t_8281), .co(t_8282), .cout(t_8283));
compressor_4_2 u2_2848(.a(t_3686), .b(t_3683), .c(t_3680), .d(t_8272), .cin(t_8274), .o(t_8284), .co(t_8285), .cout(t_8286));
compressor_4_2 u2_2849(.a(t_3610), .b(t_3698), .c(t_3695), .d(t_3692), .cin(t_3689), .o(t_8287), .co(t_8288), .cout(t_8289));
compressor_4_2 u2_2850(.a(t_3625), .b(t_3622), .c(t_3619), .d(t_3616), .cin(t_3613), .o(t_8290), .co(t_8291), .cout(t_8292));
compressor_4_2 u2_2851(.a(t_3640), .b(t_3637), .c(t_3634), .d(t_3631), .cin(t_3628), .o(t_8293), .co(t_8294), .cout(t_8295));
compressor_3_2 u1_2852(.a(t_3649), .b(t_3646), .cin(t_3643), .o(t_8296), .cout(t_8297));
compressor_4_2 u2_2853(.a(t_3707), .b(t_3704), .c(t_3701), .d(t_8277), .cin(t_8280), .o(t_8298), .co(t_8299), .cout(t_8300));
compressor_4_2 u2_2854(.a(t_3716), .b(t_3713), .c(t_3710), .d(t_8283), .cin(t_8286), .o(t_8301), .co(t_8302), .cout(t_8303));
compressor_4_2 u2_2855(.a(t_3725), .b(t_3722), .c(t_3719), .d(t_8289), .cin(t_8292), .o(t_8304), .co(t_8305), .cout(t_8306));
compressor_4_2 u2_2856(.a(t_3734), .b(t_3731), .c(t_3728), .d(t_8295), .cin(t_8297), .o(t_8307), .co(t_8308), .cout(t_8309));
compressor_4_2 u2_2857(.a(t_3660), .b(t_3657), .c(t_3743), .d(t_3740), .cin(t_3737), .o(t_8310), .co(t_8311), .cout(t_8312));
compressor_4_2 u2_2858(.a(t_3675), .b(t_3672), .c(t_3669), .d(t_3666), .cin(t_3663), .o(t_8313), .co(t_8314), .cout(t_8315));
compressor_4_2 u2_2859(.a(t_3690), .b(t_3687), .c(t_3684), .d(t_3681), .cin(t_3678), .o(t_8316), .co(t_8317), .cout(t_8318));
compressor_3_2 u1_2860(.a(t_3699), .b(t_3696), .cin(t_3693), .o(t_8319), .cout(t_8320));
compressor_4_2 u2_2861(.a(t_3749), .b(t_3746), .c(s_140_58), .d(t_8300), .cin(t_8303), .o(t_8321), .co(t_8322), .cout(t_8323));
compressor_4_2 u2_2862(.a(t_3758), .b(t_3755), .c(t_3752), .d(t_8306), .cin(t_8309), .o(t_8324), .co(t_8325), .cout(t_8326));
compressor_4_2 u2_2863(.a(t_3767), .b(t_3764), .c(t_3761), .d(t_8312), .cin(t_8315), .o(t_8327), .co(t_8328), .cout(t_8329));
compressor_4_2 u2_2864(.a(t_3776), .b(t_3773), .c(t_3770), .d(t_8318), .cin(t_8320), .o(t_8330), .co(t_8331), .cout(t_8332));
compressor_4_2 u2_2865(.a(t_3702), .b(t_3788), .c(t_3785), .d(t_3782), .cin(t_3779), .o(t_8333), .co(t_8334), .cout(t_8335));
compressor_4_2 u2_2866(.a(t_3717), .b(t_3714), .c(t_3711), .d(t_3708), .cin(t_3705), .o(t_8336), .co(t_8337), .cout(t_8338));
compressor_4_2 u2_2867(.a(t_3732), .b(t_3729), .c(t_3726), .d(t_3723), .cin(t_3720), .o(t_8339), .co(t_8340), .cout(t_8341));
compressor_3_2 u1_2868(.a(t_3741), .b(t_3738), .cin(t_3735), .o(t_8342), .cout(t_8343));
compressor_4_2 u2_2869(.a(t_3793), .b(t_3790), .c(s_141_58), .d(t_8323), .cin(t_8326), .o(t_8344), .co(t_8345), .cout(t_8346));
compressor_4_2 u2_2870(.a(t_3802), .b(t_3799), .c(t_3796), .d(t_8329), .cin(t_8332), .o(t_8347), .co(t_8348), .cout(t_8349));
compressor_4_2 u2_2871(.a(t_3811), .b(t_3808), .c(t_3805), .d(t_8335), .cin(t_8338), .o(t_8350), .co(t_8351), .cout(t_8352));
compressor_4_2 u2_2872(.a(t_3820), .b(t_3817), .c(t_3814), .d(t_8341), .cin(t_8343), .o(t_8353), .co(t_8354), .cout(t_8355));
compressor_4_2 u2_2873(.a(t_3747), .b(t_3832), .c(t_3829), .d(t_3826), .cin(t_3823), .o(t_8356), .co(t_8357), .cout(t_8358));
compressor_4_2 u2_2874(.a(t_3762), .b(t_3759), .c(t_3756), .d(t_3753), .cin(t_3750), .o(t_8359), .co(t_8360), .cout(t_8361));
compressor_4_2 u2_2875(.a(t_3777), .b(t_3774), .c(t_3771), .d(t_3768), .cin(t_3765), .o(t_8362), .co(t_8363), .cout(t_8364));
compressor_3_2 u1_2876(.a(t_3786), .b(t_3783), .cin(t_3780), .o(t_8365), .cout(t_8366));
compressor_4_2 u2_2877(.a(t_3840), .b(t_3837), .c(t_3834), .d(t_8346), .cin(t_8349), .o(t_8367), .co(t_8368), .cout(t_8369));
compressor_4_2 u2_2878(.a(t_3849), .b(t_3846), .c(t_3843), .d(t_8352), .cin(t_8355), .o(t_8370), .co(t_8371), .cout(t_8372));
compressor_4_2 u2_2879(.a(t_3858), .b(t_3855), .c(t_3852), .d(t_8358), .cin(t_8361), .o(t_8373), .co(t_8374), .cout(t_8375));
compressor_4_2 u2_2880(.a(t_3867), .b(t_3864), .c(t_3861), .d(t_8364), .cin(t_8366), .o(t_8376), .co(t_8377), .cout(t_8378));
compressor_4_2 u2_2881(.a(t_3794), .b(t_3791), .c(t_3876), .d(t_3873), .cin(t_3870), .o(t_8379), .co(t_8380), .cout(t_8381));
compressor_4_2 u2_2882(.a(t_3809), .b(t_3806), .c(t_3803), .d(t_3800), .cin(t_3797), .o(t_8382), .co(t_8383), .cout(t_8384));
compressor_4_2 u2_2883(.a(t_3824), .b(t_3821), .c(t_3818), .d(t_3815), .cin(t_3812), .o(t_8385), .co(t_8386), .cout(t_8387));
half_adder u0_2884(.a(t_3830), .b(t_3827), .o(t_8388), .cout(t_8389));
compressor_4_2 u2_2885(.a(t_3884), .b(t_3881), .c(t_3878), .d(t_8369), .cin(t_8372), .o(t_8390), .co(t_8391), .cout(t_8392));
compressor_4_2 u2_2886(.a(t_3893), .b(t_3890), .c(t_3887), .d(t_8375), .cin(t_8378), .o(t_8393), .co(t_8394), .cout(t_8395));
compressor_4_2 u2_2887(.a(t_3902), .b(t_3899), .c(t_3896), .d(t_8381), .cin(t_8384), .o(t_8396), .co(t_8397), .cout(t_8398));
compressor_4_2 u2_2888(.a(t_3911), .b(t_3908), .c(t_3905), .d(t_8387), .cin(t_8389), .o(t_8399), .co(t_8400), .cout(t_8401));
compressor_4_2 u2_2889(.a(t_3838), .b(t_3835), .c(t_3920), .d(t_3917), .cin(t_3914), .o(t_8402), .co(t_8403), .cout(t_8404));
compressor_4_2 u2_2890(.a(t_3853), .b(t_3850), .c(t_3847), .d(t_3844), .cin(t_3841), .o(t_8405), .co(t_8406), .cout(t_8407));
compressor_4_2 u2_2891(.a(t_3868), .b(t_3865), .c(t_3862), .d(t_3859), .cin(t_3856), .o(t_8408), .co(t_8409), .cout(t_8410));
half_adder u0_2892(.a(t_3874), .b(t_3871), .o(t_8411), .cout(t_8412));
compressor_4_2 u2_2893(.a(t_3928), .b(t_3925), .c(t_3922), .d(t_8392), .cin(t_8395), .o(t_8413), .co(t_8414), .cout(t_8415));
compressor_4_2 u2_2894(.a(t_3937), .b(t_3934), .c(t_3931), .d(t_8398), .cin(t_8401), .o(t_8416), .co(t_8417), .cout(t_8418));
compressor_4_2 u2_2895(.a(t_3946), .b(t_3943), .c(t_3940), .d(t_8404), .cin(t_8407), .o(t_8419), .co(t_8420), .cout(t_8421));
compressor_4_2 u2_2896(.a(t_3955), .b(t_3952), .c(t_3949), .d(t_8410), .cin(t_8412), .o(t_8422), .co(t_8423), .cout(t_8424));
compressor_4_2 u2_2897(.a(t_3882), .b(t_3879), .c(t_3964), .d(t_3961), .cin(t_3958), .o(t_8425), .co(t_8426), .cout(t_8427));
compressor_4_2 u2_2898(.a(t_3897), .b(t_3894), .c(t_3891), .d(t_3888), .cin(t_3885), .o(t_8428), .co(t_8429), .cout(t_8430));
compressor_4_2 u2_2899(.a(t_3912), .b(t_3909), .c(t_3906), .d(t_3903), .cin(t_3900), .o(t_8431), .co(t_8432), .cout(t_8433));
half_adder u0_2900(.a(t_3918), .b(t_3915), .o(t_8434), .cout(t_8435));
compressor_4_2 u2_2901(.a(t_3972), .b(t_3969), .c(t_3966), .d(t_8415), .cin(t_8418), .o(t_8436), .co(t_8437), .cout(t_8438));
compressor_4_2 u2_2902(.a(t_3981), .b(t_3978), .c(t_3975), .d(t_8421), .cin(t_8424), .o(t_8439), .co(t_8440), .cout(t_8441));
compressor_4_2 u2_2903(.a(t_3990), .b(t_3987), .c(t_3984), .d(t_8427), .cin(t_8430), .o(t_8442), .co(t_8443), .cout(t_8444));
compressor_4_2 u2_2904(.a(t_3999), .b(t_3996), .c(t_3993), .d(t_8433), .cin(t_8435), .o(t_8445), .co(t_8446), .cout(t_8447));
compressor_4_2 u2_2905(.a(t_3926), .b(t_3923), .c(t_4008), .d(t_4005), .cin(t_4002), .o(t_8448), .co(t_8449), .cout(t_8450));
compressor_4_2 u2_2906(.a(t_3941), .b(t_3938), .c(t_3935), .d(t_3932), .cin(t_3929), .o(t_8451), .co(t_8452), .cout(t_8453));
compressor_4_2 u2_2907(.a(t_3956), .b(t_3953), .c(t_3950), .d(t_3947), .cin(t_3944), .o(t_8454), .co(t_8455), .cout(t_8456));
half_adder u0_2908(.a(t_3962), .b(t_3959), .o(t_8457), .cout(t_8458));
compressor_4_2 u2_2909(.a(t_4013), .b(t_4010), .c(s_146_55), .d(t_8438), .cin(t_8441), .o(t_8459), .co(t_8460), .cout(t_8461));
compressor_4_2 u2_2910(.a(t_4022), .b(t_4019), .c(t_4016), .d(t_8444), .cin(t_8447), .o(t_8462), .co(t_8463), .cout(t_8464));
compressor_4_2 u2_2911(.a(t_4031), .b(t_4028), .c(t_4025), .d(t_8450), .cin(t_8453), .o(t_8465), .co(t_8466), .cout(t_8467));
compressor_4_2 u2_2912(.a(t_4040), .b(t_4037), .c(t_4034), .d(t_8456), .cin(t_8458), .o(t_8468), .co(t_8469), .cout(t_8470));
compressor_4_2 u2_2913(.a(t_3970), .b(t_3967), .c(t_4049), .d(t_4046), .cin(t_4043), .o(t_8471), .co(t_8472), .cout(t_8473));
compressor_4_2 u2_2914(.a(t_3985), .b(t_3982), .c(t_3979), .d(t_3976), .cin(t_3973), .o(t_8474), .co(t_8475), .cout(t_8476));
compressor_4_2 u2_2915(.a(t_4000), .b(t_3997), .c(t_3994), .d(t_3991), .cin(t_3988), .o(t_8477), .co(t_8478), .cout(t_8479));
half_adder u0_2916(.a(t_4006), .b(t_4003), .o(t_8480), .cout(t_8481));
compressor_4_2 u2_2917(.a(t_4058), .b(t_4055), .c(t_4052), .d(t_8461), .cin(t_8464), .o(t_8482), .co(t_8483), .cout(t_8484));
compressor_4_2 u2_2918(.a(t_4067), .b(t_4064), .c(t_4061), .d(t_8467), .cin(t_8470), .o(t_8485), .co(t_8486), .cout(t_8487));
compressor_4_2 u2_2919(.a(t_4076), .b(t_4073), .c(t_4070), .d(t_8473), .cin(t_8476), .o(t_8488), .co(t_8489), .cout(t_8490));
compressor_4_2 u2_2920(.a(t_4085), .b(t_4082), .c(t_4079), .d(t_8479), .cin(t_8481), .o(t_8491), .co(t_8492), .cout(t_8493));
compressor_4_2 u2_2921(.a(t_4017), .b(t_4014), .c(t_4011), .d(t_4091), .cin(t_4088), .o(t_8494), .co(t_8495), .cout(t_8496));
compressor_4_2 u2_2922(.a(t_4032), .b(t_4029), .c(t_4026), .d(t_4023), .cin(t_4020), .o(t_8497), .co(t_8498), .cout(t_8499));
compressor_4_2 u2_2923(.a(t_4047), .b(t_4044), .c(t_4041), .d(t_4038), .cin(t_4035), .o(t_8500), .co(t_8501), .cout(t_8502));
compressor_4_2 u2_2924(.a(t_4097), .b(t_4094), .c(s_148_54), .d(t_8484), .cin(t_8487), .o(t_8503), .co(t_8504), .cout(t_8505));
compressor_4_2 u2_2925(.a(t_4106), .b(t_4103), .c(t_4100), .d(t_8490), .cin(t_8493), .o(t_8506), .co(t_8507), .cout(t_8508));
compressor_4_2 u2_2926(.a(t_4115), .b(t_4112), .c(t_4109), .d(t_8496), .cin(t_8499), .o(t_8509), .co(t_8510), .cout(t_8511));
compressor_4_2 u2_2927(.a(t_4127), .b(t_4124), .c(t_4121), .d(t_4118), .cin(t_8502), .o(t_8512), .co(t_8513), .cout(t_8514));
compressor_4_2 u2_2928(.a(t_4059), .b(t_4056), .c(t_4053), .d(t_4133), .cin(t_4130), .o(t_8515), .co(t_8516), .cout(t_8517));
compressor_4_2 u2_2929(.a(t_4074), .b(t_4071), .c(t_4068), .d(t_4065), .cin(t_4062), .o(t_8518), .co(t_8519), .cout(t_8520));
compressor_4_2 u2_2930(.a(t_4089), .b(t_4086), .c(t_4083), .d(t_4080), .cin(t_4077), .o(t_8521), .co(t_8522), .cout(t_8523));
compressor_4_2 u2_2931(.a(t_4138), .b(t_4135), .c(s_149_54), .d(t_8505), .cin(t_8508), .o(t_8524), .co(t_8525), .cout(t_8526));
compressor_4_2 u2_2932(.a(t_4147), .b(t_4144), .c(t_4141), .d(t_8511), .cin(t_8514), .o(t_8527), .co(t_8528), .cout(t_8529));
compressor_4_2 u2_2933(.a(t_4156), .b(t_4153), .c(t_4150), .d(t_8517), .cin(t_8520), .o(t_8530), .co(t_8531), .cout(t_8532));
compressor_4_2 u2_2934(.a(t_4168), .b(t_4165), .c(t_4162), .d(t_4159), .cin(t_8523), .o(t_8533), .co(t_8534), .cout(t_8535));
compressor_4_2 u2_2935(.a(t_4101), .b(t_4098), .c(t_4095), .d(t_4174), .cin(t_4171), .o(t_8536), .co(t_8537), .cout(t_8538));
compressor_4_2 u2_2936(.a(t_4116), .b(t_4113), .c(t_4110), .d(t_4107), .cin(t_4104), .o(t_8539), .co(t_8540), .cout(t_8541));
compressor_4_2 u2_2937(.a(t_4131), .b(t_4128), .c(t_4125), .d(t_4122), .cin(t_4119), .o(t_8542), .co(t_8543), .cout(t_8544));
compressor_4_2 u2_2938(.a(t_4182), .b(t_4179), .c(t_4176), .d(t_8526), .cin(t_8529), .o(t_8545), .co(t_8546), .cout(t_8547));
compressor_4_2 u2_2939(.a(t_4191), .b(t_4188), .c(t_4185), .d(t_8532), .cin(t_8535), .o(t_8548), .co(t_8549), .cout(t_8550));
compressor_4_2 u2_2940(.a(t_4200), .b(t_4197), .c(t_4194), .d(t_8538), .cin(t_8541), .o(t_8551), .co(t_8552), .cout(t_8553));
compressor_4_2 u2_2941(.a(t_4212), .b(t_4209), .c(t_4206), .d(t_4203), .cin(t_8544), .o(t_8554), .co(t_8555), .cout(t_8556));
compressor_4_2 u2_2942(.a(t_4145), .b(t_4142), .c(t_4139), .d(t_4136), .cin(t_4215), .o(t_8557), .co(t_8558), .cout(t_8559));
compressor_4_2 u2_2943(.a(t_4160), .b(t_4157), .c(t_4154), .d(t_4151), .cin(t_4148), .o(t_8560), .co(t_8561), .cout(t_8562));
compressor_3_2 u1_2944(.a(t_4169), .b(t_4166), .cin(t_4163), .o(t_8563), .cout(t_8564));
compressor_4_2 u2_2945(.a(t_4223), .b(t_4220), .c(t_4217), .d(t_8547), .cin(t_8550), .o(t_8565), .co(t_8566), .cout(t_8567));
compressor_4_2 u2_2946(.a(t_4232), .b(t_4229), .c(t_4226), .d(t_8553), .cin(t_8556), .o(t_8568), .co(t_8569), .cout(t_8570));
compressor_4_2 u2_2947(.a(t_4241), .b(t_4238), .c(t_4235), .d(t_8559), .cin(t_8562), .o(t_8571), .co(t_8572), .cout(t_8573));
compressor_4_2 u2_2948(.a(t_4253), .b(t_4250), .c(t_4247), .d(t_4244), .cin(t_8564), .o(t_8574), .co(t_8575), .cout(t_8576));
compressor_4_2 u2_2949(.a(t_4186), .b(t_4183), .c(t_4180), .d(t_4177), .cin(t_4256), .o(t_8577), .co(t_8578), .cout(t_8579));
compressor_4_2 u2_2950(.a(t_4201), .b(t_4198), .c(t_4195), .d(t_4192), .cin(t_4189), .o(t_8580), .co(t_8581), .cout(t_8582));
compressor_3_2 u1_2951(.a(t_4210), .b(t_4207), .cin(t_4204), .o(t_8583), .cout(t_8584));
compressor_4_2 u2_2952(.a(t_4264), .b(t_4261), .c(t_4258), .d(t_8567), .cin(t_8570), .o(t_8585), .co(t_8586), .cout(t_8587));
compressor_4_2 u2_2953(.a(t_4273), .b(t_4270), .c(t_4267), .d(t_8573), .cin(t_8576), .o(t_8588), .co(t_8589), .cout(t_8590));
compressor_4_2 u2_2954(.a(t_4282), .b(t_4279), .c(t_4276), .d(t_8579), .cin(t_8582), .o(t_8591), .co(t_8592), .cout(t_8593));
compressor_4_2 u2_2955(.a(t_4294), .b(t_4291), .c(t_4288), .d(t_4285), .cin(t_8584), .o(t_8594), .co(t_8595), .cout(t_8596));
compressor_4_2 u2_2956(.a(t_4227), .b(t_4224), .c(t_4221), .d(t_4218), .cin(t_4297), .o(t_8597), .co(t_8598), .cout(t_8599));
compressor_4_2 u2_2957(.a(t_4242), .b(t_4239), .c(t_4236), .d(t_4233), .cin(t_4230), .o(t_8600), .co(t_8601), .cout(t_8602));
compressor_3_2 u1_2958(.a(t_4251), .b(t_4248), .cin(t_4245), .o(t_8603), .cout(t_8604));
compressor_4_2 u2_2959(.a(t_4305), .b(t_4302), .c(t_4299), .d(t_8587), .cin(t_8590), .o(t_8605), .co(t_8606), .cout(t_8607));
compressor_4_2 u2_2960(.a(t_4314), .b(t_4311), .c(t_4308), .d(t_8593), .cin(t_8596), .o(t_8608), .co(t_8609), .cout(t_8610));
compressor_4_2 u2_2961(.a(t_4323), .b(t_4320), .c(t_4317), .d(t_8599), .cin(t_8602), .o(t_8611), .co(t_8612), .cout(t_8613));
compressor_4_2 u2_2962(.a(t_4335), .b(t_4332), .c(t_4329), .d(t_4326), .cin(t_8604), .o(t_8614), .co(t_8615), .cout(t_8616));
compressor_4_2 u2_2963(.a(t_4268), .b(t_4265), .c(t_4262), .d(t_4259), .cin(t_4338), .o(t_8617), .co(t_8618), .cout(t_8619));
compressor_4_2 u2_2964(.a(t_4283), .b(t_4280), .c(t_4277), .d(t_4274), .cin(t_4271), .o(t_8620), .co(t_8621), .cout(t_8622));
compressor_3_2 u1_2965(.a(t_4292), .b(t_4289), .cin(t_4286), .o(t_8623), .cout(t_8624));
compressor_4_2 u2_2966(.a(t_4343), .b(t_4340), .c(s_154_51), .d(t_8607), .cin(t_8610), .o(t_8625), .co(t_8626), .cout(t_8627));
compressor_4_2 u2_2967(.a(t_4352), .b(t_4349), .c(t_4346), .d(t_8613), .cin(t_8616), .o(t_8628), .co(t_8629), .cout(t_8630));
compressor_4_2 u2_2968(.a(t_4361), .b(t_4358), .c(t_4355), .d(t_8619), .cin(t_8622), .o(t_8631), .co(t_8632), .cout(t_8633));
compressor_4_2 u2_2969(.a(t_4373), .b(t_4370), .c(t_4367), .d(t_4364), .cin(t_8624), .o(t_8634), .co(t_8635), .cout(t_8636));
compressor_4_2 u2_2970(.a(t_4309), .b(t_4306), .c(t_4303), .d(t_4300), .cin(t_4376), .o(t_8637), .co(t_8638), .cout(t_8639));
compressor_4_2 u2_2971(.a(t_4324), .b(t_4321), .c(t_4318), .d(t_4315), .cin(t_4312), .o(t_8640), .co(t_8641), .cout(t_8642));
compressor_3_2 u1_2972(.a(t_4333), .b(t_4330), .cin(t_4327), .o(t_8643), .cout(t_8644));
compressor_4_2 u2_2973(.a(t_4385), .b(t_4382), .c(t_4379), .d(t_8627), .cin(t_8630), .o(t_8645), .co(t_8646), .cout(t_8647));
compressor_4_2 u2_2974(.a(t_4394), .b(t_4391), .c(t_4388), .d(t_8633), .cin(t_8636), .o(t_8648), .co(t_8649), .cout(t_8650));
compressor_4_2 u2_2975(.a(t_4403), .b(t_4400), .c(t_4397), .d(t_8639), .cin(t_8642), .o(t_8651), .co(t_8652), .cout(t_8653));
compressor_4_2 u2_2976(.a(t_4415), .b(t_4412), .c(t_4409), .d(t_4406), .cin(t_8644), .o(t_8654), .co(t_8655), .cout(t_8656));
compressor_4_2 u2_2977(.a(t_4353), .b(t_4350), .c(t_4347), .d(t_4344), .cin(t_4341), .o(t_8657), .co(t_8658), .cout(t_8659));
compressor_4_2 u2_2978(.a(t_4368), .b(t_4365), .c(t_4362), .d(t_4359), .cin(t_4356), .o(t_8660), .co(t_8661), .cout(t_8662));
compressor_3_2 u1_2979(.a(t_4377), .b(t_4374), .cin(t_4371), .o(t_8663), .cout(t_8664));
compressor_4_2 u2_2980(.a(t_4421), .b(t_4418), .c(s_156_50), .d(t_8647), .cin(t_8650), .o(t_8665), .co(t_8666), .cout(t_8667));
compressor_4_2 u2_2981(.a(t_4430), .b(t_4427), .c(t_4424), .d(t_8653), .cin(t_8656), .o(t_8668), .co(t_8669), .cout(t_8670));
compressor_4_2 u2_2982(.a(t_4439), .b(t_4436), .c(t_4433), .d(t_8659), .cin(t_8662), .o(t_8671), .co(t_8672), .cout(t_8673));
compressor_4_2 u2_2983(.a(t_4451), .b(t_4448), .c(t_4445), .d(t_4442), .cin(t_8664), .o(t_8674), .co(t_8675), .cout(t_8676));
compressor_4_2 u2_2984(.a(t_4389), .b(t_4386), .c(t_4383), .d(t_4380), .cin(t_4454), .o(t_8677), .co(t_8678), .cout(t_8679));
compressor_4_2 u2_2985(.a(t_4404), .b(t_4401), .c(t_4398), .d(t_4395), .cin(t_4392), .o(t_8680), .co(t_8681), .cout(t_8682));
compressor_3_2 u1_2986(.a(t_4413), .b(t_4410), .cin(t_4407), .o(t_8683), .cout(t_8684));
compressor_4_2 u2_2987(.a(t_4459), .b(t_4456), .c(s_157_50), .d(t_8667), .cin(t_8670), .o(t_8685), .co(t_8686), .cout(t_8687));
compressor_4_2 u2_2988(.a(t_4468), .b(t_4465), .c(t_4462), .d(t_8673), .cin(t_8676), .o(t_8688), .co(t_8689), .cout(t_8690));
compressor_4_2 u2_2989(.a(t_4477), .b(t_4474), .c(t_4471), .d(t_8679), .cin(t_8682), .o(t_8691), .co(t_8692), .cout(t_8693));
compressor_4_2 u2_2990(.a(t_4489), .b(t_4486), .c(t_4483), .d(t_4480), .cin(t_8684), .o(t_8694), .co(t_8695), .cout(t_8696));
compressor_4_2 u2_2991(.a(t_4428), .b(t_4425), .c(t_4422), .d(t_4419), .cin(t_4492), .o(t_8697), .co(t_8698), .cout(t_8699));
compressor_4_2 u2_2992(.a(t_4443), .b(t_4440), .c(t_4437), .d(t_4434), .cin(t_4431), .o(t_8700), .co(t_8701), .cout(t_8702));
compressor_3_2 u1_2993(.a(t_4452), .b(t_4449), .cin(t_4446), .o(t_8703), .cout(t_8704));
compressor_4_2 u2_2994(.a(t_4500), .b(t_4497), .c(t_4494), .d(t_8687), .cin(t_8690), .o(t_8705), .co(t_8706), .cout(t_8707));
compressor_4_2 u2_2995(.a(t_4509), .b(t_4506), .c(t_4503), .d(t_8693), .cin(t_8696), .o(t_8708), .co(t_8709), .cout(t_8710));
compressor_4_2 u2_2996(.a(t_4518), .b(t_4515), .c(t_4512), .d(t_8699), .cin(t_8702), .o(t_8711), .co(t_8712), .cout(t_8713));
compressor_4_2 u2_2997(.a(t_4530), .b(t_4527), .c(t_4524), .d(t_4521), .cin(t_8704), .o(t_8714), .co(t_8715), .cout(t_8716));
compressor_4_2 u2_2998(.a(t_4469), .b(t_4466), .c(t_4463), .d(t_4460), .cin(t_4457), .o(t_8717), .co(t_8718), .cout(t_8719));
compressor_4_2 u2_2999(.a(t_4484), .b(t_4481), .c(t_4478), .d(t_4475), .cin(t_4472), .o(t_8720), .co(t_8721), .cout(t_8722));
half_adder u0_3000(.a(t_4490), .b(t_4487), .o(t_8723), .cout(t_8724));
compressor_4_2 u2_3001(.a(t_4538), .b(t_4535), .c(t_4532), .d(t_8707), .cin(t_8710), .o(t_8725), .co(t_8726), .cout(t_8727));
compressor_4_2 u2_3002(.a(t_4547), .b(t_4544), .c(t_4541), .d(t_8713), .cin(t_8716), .o(t_8728), .co(t_8729), .cout(t_8730));
compressor_4_2 u2_3003(.a(t_4556), .b(t_4553), .c(t_4550), .d(t_8719), .cin(t_8722), .o(t_8731), .co(t_8732), .cout(t_8733));
compressor_4_2 u2_3004(.a(t_4568), .b(t_4565), .c(t_4562), .d(t_4559), .cin(t_8724), .o(t_8734), .co(t_8735), .cout(t_8736));
compressor_4_2 u2_3005(.a(t_4507), .b(t_4504), .c(t_4501), .d(t_4498), .cin(t_4495), .o(t_8737), .co(t_8738), .cout(t_8739));
compressor_4_2 u2_3006(.a(t_4522), .b(t_4519), .c(t_4516), .d(t_4513), .cin(t_4510), .o(t_8740), .co(t_8741), .cout(t_8742));
half_adder u0_3007(.a(t_4528), .b(t_4525), .o(t_8743), .cout(t_8744));
compressor_4_2 u2_3008(.a(t_4576), .b(t_4573), .c(t_4570), .d(t_8727), .cin(t_8730), .o(t_8745), .co(t_8746), .cout(t_8747));
compressor_4_2 u2_3009(.a(t_4585), .b(t_4582), .c(t_4579), .d(t_8733), .cin(t_8736), .o(t_8748), .co(t_8749), .cout(t_8750));
compressor_4_2 u2_3010(.a(t_4594), .b(t_4591), .c(t_4588), .d(t_8739), .cin(t_8742), .o(t_8751), .co(t_8752), .cout(t_8753));
compressor_4_2 u2_3011(.a(t_4606), .b(t_4603), .c(t_4600), .d(t_4597), .cin(t_8744), .o(t_8754), .co(t_8755), .cout(t_8756));
compressor_4_2 u2_3012(.a(t_4545), .b(t_4542), .c(t_4539), .d(t_4536), .cin(t_4533), .o(t_8757), .co(t_8758), .cout(t_8759));
compressor_4_2 u2_3013(.a(t_4560), .b(t_4557), .c(t_4554), .d(t_4551), .cin(t_4548), .o(t_8760), .co(t_8761), .cout(t_8762));
half_adder u0_3014(.a(t_4566), .b(t_4563), .o(t_8763), .cout(t_8764));
compressor_4_2 u2_3015(.a(t_4614), .b(t_4611), .c(t_4608), .d(t_8747), .cin(t_8750), .o(t_8765), .co(t_8766), .cout(t_8767));
compressor_4_2 u2_3016(.a(t_4623), .b(t_4620), .c(t_4617), .d(t_8753), .cin(t_8756), .o(t_8768), .co(t_8769), .cout(t_8770));
compressor_4_2 u2_3017(.a(t_4632), .b(t_4629), .c(t_4626), .d(t_8759), .cin(t_8762), .o(t_8771), .co(t_8772), .cout(t_8773));
compressor_4_2 u2_3018(.a(t_4644), .b(t_4641), .c(t_4638), .d(t_4635), .cin(t_8764), .o(t_8774), .co(t_8775), .cout(t_8776));
compressor_4_2 u2_3019(.a(t_4583), .b(t_4580), .c(t_4577), .d(t_4574), .cin(t_4571), .o(t_8777), .co(t_8778), .cout(t_8779));
compressor_4_2 u2_3020(.a(t_4598), .b(t_4595), .c(t_4592), .d(t_4589), .cin(t_4586), .o(t_8780), .co(t_8781), .cout(t_8782));
half_adder u0_3021(.a(t_4604), .b(t_4601), .o(t_8783), .cout(t_8784));
compressor_4_2 u2_3022(.a(t_4649), .b(t_4646), .c(s_162_47), .d(t_8767), .cin(t_8770), .o(t_8785), .co(t_8786), .cout(t_8787));
compressor_4_2 u2_3023(.a(t_4658), .b(t_4655), .c(t_4652), .d(t_8773), .cin(t_8776), .o(t_8788), .co(t_8789), .cout(t_8790));
compressor_4_2 u2_3024(.a(t_4667), .b(t_4664), .c(t_4661), .d(t_8779), .cin(t_8782), .o(t_8791), .co(t_8792), .cout(t_8793));
compressor_4_2 u2_3025(.a(t_4679), .b(t_4676), .c(t_4673), .d(t_4670), .cin(t_8784), .o(t_8794), .co(t_8795), .cout(t_8796));
compressor_4_2 u2_3026(.a(t_4621), .b(t_4618), .c(t_4615), .d(t_4612), .cin(t_4609), .o(t_8797), .co(t_8798), .cout(t_8799));
compressor_4_2 u2_3027(.a(t_4636), .b(t_4633), .c(t_4630), .d(t_4627), .cin(t_4624), .o(t_8800), .co(t_8801), .cout(t_8802));
half_adder u0_3028(.a(t_4642), .b(t_4639), .o(t_8803), .cout(t_8804));
compressor_4_2 u2_3029(.a(t_4688), .b(t_4685), .c(t_4682), .d(t_8787), .cin(t_8790), .o(t_8805), .co(t_8806), .cout(t_8807));
compressor_4_2 u2_3030(.a(t_4697), .b(t_4694), .c(t_4691), .d(t_8793), .cin(t_8796), .o(t_8808), .co(t_8809), .cout(t_8810));
compressor_4_2 u2_3031(.a(t_4706), .b(t_4703), .c(t_4700), .d(t_8799), .cin(t_8802), .o(t_8811), .co(t_8812), .cout(t_8813));
compressor_4_2 u2_3032(.a(t_4647), .b(t_4715), .c(t_4712), .d(t_4709), .cin(t_8804), .o(t_8814), .co(t_8815), .cout(t_8816));
compressor_4_2 u2_3033(.a(t_4662), .b(t_4659), .c(t_4656), .d(t_4653), .cin(t_4650), .o(t_8817), .co(t_8818), .cout(t_8819));
compressor_4_2 u2_3034(.a(t_4677), .b(t_4674), .c(t_4671), .d(t_4668), .cin(t_4665), .o(t_8820), .co(t_8821), .cout(t_8822));
compressor_4_2 u2_3035(.a(t_4721), .b(t_4718), .c(s_164_46), .d(t_8807), .cin(t_8810), .o(t_8823), .co(t_8824), .cout(t_8825));
compressor_4_2 u2_3036(.a(t_4730), .b(t_4727), .c(t_4724), .d(t_8813), .cin(t_8816), .o(t_8826), .co(t_8827), .cout(t_8828));
compressor_4_2 u2_3037(.a(t_4739), .b(t_4736), .c(t_4733), .d(t_8819), .cin(t_8822), .o(t_8829), .co(t_8830), .cout(t_8831));
compressor_4_2 u2_3038(.a(t_4683), .b(t_4751), .c(t_4748), .d(t_4745), .cin(t_4742), .o(t_8832), .co(t_8833), .cout(t_8834));
compressor_4_2 u2_3039(.a(t_4698), .b(t_4695), .c(t_4692), .d(t_4689), .cin(t_4686), .o(t_8835), .co(t_8836), .cout(t_8837));
compressor_4_2 u2_3040(.a(t_4713), .b(t_4710), .c(t_4707), .d(t_4704), .cin(t_4701), .o(t_8838), .co(t_8839), .cout(t_8840));
compressor_4_2 u2_3041(.a(t_4756), .b(t_4753), .c(s_165_46), .d(t_8825), .cin(t_8828), .o(t_8841), .co(t_8842), .cout(t_8843));
compressor_4_2 u2_3042(.a(t_4765), .b(t_4762), .c(t_4759), .d(t_8831), .cin(t_8834), .o(t_8844), .co(t_8845), .cout(t_8846));
compressor_4_2 u2_3043(.a(t_4774), .b(t_4771), .c(t_4768), .d(t_8837), .cin(t_8840), .o(t_8847), .co(t_8848), .cout(t_8849));
compressor_4_2 u2_3044(.a(t_4719), .b(t_4786), .c(t_4783), .d(t_4780), .cin(t_4777), .o(t_8850), .co(t_8851), .cout(t_8852));
compressor_4_2 u2_3045(.a(t_4734), .b(t_4731), .c(t_4728), .d(t_4725), .cin(t_4722), .o(t_8853), .co(t_8854), .cout(t_8855));
compressor_4_2 u2_3046(.a(t_4749), .b(t_4746), .c(t_4743), .d(t_4740), .cin(t_4737), .o(t_8856), .co(t_8857), .cout(t_8858));
compressor_4_2 u2_3047(.a(t_4794), .b(t_4791), .c(t_4788), .d(t_8843), .cin(t_8846), .o(t_8859), .co(t_8860), .cout(t_8861));
compressor_4_2 u2_3048(.a(t_4803), .b(t_4800), .c(t_4797), .d(t_8849), .cin(t_8852), .o(t_8862), .co(t_8863), .cout(t_8864));
compressor_4_2 u2_3049(.a(t_4812), .b(t_4809), .c(t_4806), .d(t_8855), .cin(t_8858), .o(t_8865), .co(t_8866), .cout(t_8867));
compressor_4_2 u2_3050(.a(t_4757), .b(t_4754), .c(t_4821), .d(t_4818), .cin(t_4815), .o(t_8868), .co(t_8869), .cout(t_8870));
compressor_4_2 u2_3051(.a(t_4772), .b(t_4769), .c(t_4766), .d(t_4763), .cin(t_4760), .o(t_8871), .co(t_8872), .cout(t_8873));
compressor_3_2 u1_3052(.a(t_4781), .b(t_4778), .cin(t_4775), .o(t_8874), .cout(t_8875));
compressor_4_2 u2_3053(.a(t_4829), .b(t_4826), .c(t_4823), .d(t_8861), .cin(t_8864), .o(t_8876), .co(t_8877), .cout(t_8878));
compressor_4_2 u2_3054(.a(t_4838), .b(t_4835), .c(t_4832), .d(t_8867), .cin(t_8870), .o(t_8879), .co(t_8880), .cout(t_8881));
compressor_4_2 u2_3055(.a(t_4847), .b(t_4844), .c(t_4841), .d(t_8873), .cin(t_8875), .o(t_8882), .co(t_8883), .cout(t_8884));
compressor_4_2 u2_3056(.a(t_4792), .b(t_4789), .c(t_4856), .d(t_4853), .cin(t_4850), .o(t_8885), .co(t_8886), .cout(t_8887));
compressor_4_2 u2_3057(.a(t_4807), .b(t_4804), .c(t_4801), .d(t_4798), .cin(t_4795), .o(t_8888), .co(t_8889), .cout(t_8890));
compressor_3_2 u1_3058(.a(t_4816), .b(t_4813), .cin(t_4810), .o(t_8891), .cout(t_8892));
compressor_4_2 u2_3059(.a(t_4864), .b(t_4861), .c(t_4858), .d(t_8878), .cin(t_8881), .o(t_8893), .co(t_8894), .cout(t_8895));
compressor_4_2 u2_3060(.a(t_4873), .b(t_4870), .c(t_4867), .d(t_8884), .cin(t_8887), .o(t_8896), .co(t_8897), .cout(t_8898));
compressor_4_2 u2_3061(.a(t_4882), .b(t_4879), .c(t_4876), .d(t_8890), .cin(t_8892), .o(t_8899), .co(t_8900), .cout(t_8901));
compressor_4_2 u2_3062(.a(t_4827), .b(t_4824), .c(t_4891), .d(t_4888), .cin(t_4885), .o(t_8902), .co(t_8903), .cout(t_8904));
compressor_4_2 u2_3063(.a(t_4842), .b(t_4839), .c(t_4836), .d(t_4833), .cin(t_4830), .o(t_8905), .co(t_8906), .cout(t_8907));
compressor_3_2 u1_3064(.a(t_4851), .b(t_4848), .cin(t_4845), .o(t_8908), .cout(t_8909));
compressor_4_2 u2_3065(.a(t_4899), .b(t_4896), .c(t_4893), .d(t_8895), .cin(t_8898), .o(t_8910), .co(t_8911), .cout(t_8912));
compressor_4_2 u2_3066(.a(t_4908), .b(t_4905), .c(t_4902), .d(t_8901), .cin(t_8904), .o(t_8913), .co(t_8914), .cout(t_8915));
compressor_4_2 u2_3067(.a(t_4917), .b(t_4914), .c(t_4911), .d(t_8907), .cin(t_8909), .o(t_8916), .co(t_8917), .cout(t_8918));
compressor_4_2 u2_3068(.a(t_4862), .b(t_4859), .c(t_4926), .d(t_4923), .cin(t_4920), .o(t_8919), .co(t_8920), .cout(t_8921));
compressor_4_2 u2_3069(.a(t_4877), .b(t_4874), .c(t_4871), .d(t_4868), .cin(t_4865), .o(t_8922), .co(t_8923), .cout(t_8924));
compressor_3_2 u1_3070(.a(t_4886), .b(t_4883), .cin(t_4880), .o(t_8925), .cout(t_8926));
compressor_4_2 u2_3071(.a(t_4931), .b(t_4928), .c(s_170_43), .d(t_8912), .cin(t_8915), .o(t_8927), .co(t_8928), .cout(t_8929));
compressor_4_2 u2_3072(.a(t_4940), .b(t_4937), .c(t_4934), .d(t_8918), .cin(t_8921), .o(t_8930), .co(t_8931), .cout(t_8932));
compressor_4_2 u2_3073(.a(t_4949), .b(t_4946), .c(t_4943), .d(t_8924), .cin(t_8926), .o(t_8933), .co(t_8934), .cout(t_8935));
compressor_4_2 u2_3074(.a(t_4897), .b(t_4894), .c(t_4958), .d(t_4955), .cin(t_4952), .o(t_8936), .co(t_8937), .cout(t_8938));
compressor_4_2 u2_3075(.a(t_4912), .b(t_4909), .c(t_4906), .d(t_4903), .cin(t_4900), .o(t_8939), .co(t_8940), .cout(t_8941));
compressor_3_2 u1_3076(.a(t_4921), .b(t_4918), .cin(t_4915), .o(t_8942), .cout(t_8943));
compressor_4_2 u2_3077(.a(t_4967), .b(t_4964), .c(t_4961), .d(t_8929), .cin(t_8932), .o(t_8944), .co(t_8945), .cout(t_8946));
compressor_4_2 u2_3078(.a(t_4976), .b(t_4973), .c(t_4970), .d(t_8935), .cin(t_8938), .o(t_8947), .co(t_8948), .cout(t_8949));
compressor_4_2 u2_3079(.a(t_4985), .b(t_4982), .c(t_4979), .d(t_8941), .cin(t_8943), .o(t_8950), .co(t_8951), .cout(t_8952));
compressor_4_2 u2_3080(.a(t_4935), .b(t_4932), .c(t_4929), .d(t_4991), .cin(t_4988), .o(t_8953), .co(t_8954), .cout(t_8955));
compressor_4_2 u2_3081(.a(t_4950), .b(t_4947), .c(t_4944), .d(t_4941), .cin(t_4938), .o(t_8956), .co(t_8957), .cout(t_8958));
compressor_3_2 u1_3082(.a(t_4959), .b(t_4956), .cin(t_4953), .o(t_8959), .cout(t_8960));
compressor_4_2 u2_3083(.a(t_4997), .b(t_4994), .c(s_172_42), .d(t_8946), .cin(t_8949), .o(t_8961), .co(t_8962), .cout(t_8963));
compressor_4_2 u2_3084(.a(t_5006), .b(t_5003), .c(t_5000), .d(t_8952), .cin(t_8955), .o(t_8964), .co(t_8965), .cout(t_8966));
compressor_4_2 u2_3085(.a(t_5015), .b(t_5012), .c(t_5009), .d(t_8958), .cin(t_8960), .o(t_8967), .co(t_8968), .cout(t_8969));
compressor_4_2 u2_3086(.a(t_4965), .b(t_4962), .c(t_5024), .d(t_5021), .cin(t_5018), .o(t_8970), .co(t_8971), .cout(t_8972));
compressor_4_2 u2_3087(.a(t_4980), .b(t_4977), .c(t_4974), .d(t_4971), .cin(t_4968), .o(t_8973), .co(t_8974), .cout(t_8975));
compressor_3_2 u1_3088(.a(t_4989), .b(t_4986), .cin(t_4983), .o(t_8976), .cout(t_8977));
compressor_4_2 u2_3089(.a(t_5029), .b(t_5026), .c(s_173_42), .d(t_8963), .cin(t_8966), .o(t_8978), .co(t_8979), .cout(t_8980));
compressor_4_2 u2_3090(.a(t_5038), .b(t_5035), .c(t_5032), .d(t_8969), .cin(t_8972), .o(t_8981), .co(t_8982), .cout(t_8983));
compressor_4_2 u2_3091(.a(t_5047), .b(t_5044), .c(t_5041), .d(t_8975), .cin(t_8977), .o(t_8984), .co(t_8985), .cout(t_8986));
compressor_4_2 u2_3092(.a(t_4998), .b(t_4995), .c(t_5056), .d(t_5053), .cin(t_5050), .o(t_8987), .co(t_8988), .cout(t_8989));
compressor_4_2 u2_3093(.a(t_5013), .b(t_5010), .c(t_5007), .d(t_5004), .cin(t_5001), .o(t_8990), .co(t_8991), .cout(t_8992));
compressor_3_2 u1_3094(.a(t_5022), .b(t_5019), .cin(t_5016), .o(t_8993), .cout(t_8994));
compressor_4_2 u2_3095(.a(t_5064), .b(t_5061), .c(t_5058), .d(t_8980), .cin(t_8983), .o(t_8995), .co(t_8996), .cout(t_8997));
compressor_4_2 u2_3096(.a(t_5073), .b(t_5070), .c(t_5067), .d(t_8986), .cin(t_8989), .o(t_8998), .co(t_8999), .cout(t_9000));
compressor_4_2 u2_3097(.a(t_5082), .b(t_5079), .c(t_5076), .d(t_8992), .cin(t_8994), .o(t_9001), .co(t_9002), .cout(t_9003));
compressor_4_2 u2_3098(.a(t_5033), .b(t_5030), .c(t_5027), .d(t_5088), .cin(t_5085), .o(t_9004), .co(t_9005), .cout(t_9006));
compressor_4_2 u2_3099(.a(t_5048), .b(t_5045), .c(t_5042), .d(t_5039), .cin(t_5036), .o(t_9007), .co(t_9008), .cout(t_9009));
half_adder u0_3100(.a(t_5054), .b(t_5051), .o(t_9010), .cout(t_9011));
compressor_4_2 u2_3101(.a(t_5096), .b(t_5093), .c(t_5090), .d(t_8997), .cin(t_9000), .o(t_9012), .co(t_9013), .cout(t_9014));
compressor_4_2 u2_3102(.a(t_5105), .b(t_5102), .c(t_5099), .d(t_9003), .cin(t_9006), .o(t_9015), .co(t_9016), .cout(t_9017));
compressor_4_2 u2_3103(.a(t_5114), .b(t_5111), .c(t_5108), .d(t_9009), .cin(t_9011), .o(t_9018), .co(t_9019), .cout(t_9020));
compressor_4_2 u2_3104(.a(t_5065), .b(t_5062), .c(t_5059), .d(t_5120), .cin(t_5117), .o(t_9021), .co(t_9022), .cout(t_9023));
compressor_4_2 u2_3105(.a(t_5080), .b(t_5077), .c(t_5074), .d(t_5071), .cin(t_5068), .o(t_9024), .co(t_9025), .cout(t_9026));
half_adder u0_3106(.a(t_5086), .b(t_5083), .o(t_9027), .cout(t_9028));
compressor_4_2 u2_3107(.a(t_5128), .b(t_5125), .c(t_5122), .d(t_9014), .cin(t_9017), .o(t_9029), .co(t_9030), .cout(t_9031));
compressor_4_2 u2_3108(.a(t_5137), .b(t_5134), .c(t_5131), .d(t_9020), .cin(t_9023), .o(t_9032), .co(t_9033), .cout(t_9034));
compressor_4_2 u2_3109(.a(t_5146), .b(t_5143), .c(t_5140), .d(t_9026), .cin(t_9028), .o(t_9035), .co(t_9036), .cout(t_9037));
compressor_4_2 u2_3110(.a(t_5097), .b(t_5094), .c(t_5091), .d(t_5152), .cin(t_5149), .o(t_9038), .co(t_9039), .cout(t_9040));
compressor_4_2 u2_3111(.a(t_5112), .b(t_5109), .c(t_5106), .d(t_5103), .cin(t_5100), .o(t_9041), .co(t_9042), .cout(t_9043));
half_adder u0_3112(.a(t_5118), .b(t_5115), .o(t_9044), .cout(t_9045));
compressor_4_2 u2_3113(.a(t_5160), .b(t_5157), .c(t_5154), .d(t_9031), .cin(t_9034), .o(t_9046), .co(t_9047), .cout(t_9048));
compressor_4_2 u2_3114(.a(t_5169), .b(t_5166), .c(t_5163), .d(t_9037), .cin(t_9040), .o(t_9049), .co(t_9050), .cout(t_9051));
compressor_4_2 u2_3115(.a(t_5178), .b(t_5175), .c(t_5172), .d(t_9043), .cin(t_9045), .o(t_9052), .co(t_9053), .cout(t_9054));
compressor_4_2 u2_3116(.a(t_5129), .b(t_5126), .c(t_5123), .d(t_5184), .cin(t_5181), .o(t_9055), .co(t_9056), .cout(t_9057));
compressor_4_2 u2_3117(.a(t_5144), .b(t_5141), .c(t_5138), .d(t_5135), .cin(t_5132), .o(t_9058), .co(t_9059), .cout(t_9060));
half_adder u0_3118(.a(t_5150), .b(t_5147), .o(t_9061), .cout(t_9062));
compressor_4_2 u2_3119(.a(t_5189), .b(t_5186), .c(s_178_39), .d(t_9048), .cin(t_9051), .o(t_9063), .co(t_9064), .cout(t_9065));
compressor_4_2 u2_3120(.a(t_5198), .b(t_5195), .c(t_5192), .d(t_9054), .cin(t_9057), .o(t_9066), .co(t_9067), .cout(t_9068));
compressor_4_2 u2_3121(.a(t_5207), .b(t_5204), .c(t_5201), .d(t_9060), .cin(t_9062), .o(t_9069), .co(t_9070), .cout(t_9071));
compressor_4_2 u2_3122(.a(t_5161), .b(t_5158), .c(t_5155), .d(t_5213), .cin(t_5210), .o(t_9072), .co(t_9073), .cout(t_9074));
compressor_4_2 u2_3123(.a(t_5176), .b(t_5173), .c(t_5170), .d(t_5167), .cin(t_5164), .o(t_9075), .co(t_9076), .cout(t_9077));
half_adder u0_3124(.a(t_5182), .b(t_5179), .o(t_9078), .cout(t_9079));
compressor_4_2 u2_3125(.a(t_5222), .b(t_5219), .c(t_5216), .d(t_9065), .cin(t_9068), .o(t_9080), .co(t_9081), .cout(t_9082));
compressor_4_2 u2_3126(.a(t_5231), .b(t_5228), .c(t_5225), .d(t_9071), .cin(t_9074), .o(t_9083), .co(t_9084), .cout(t_9085));
compressor_4_2 u2_3127(.a(t_5240), .b(t_5237), .c(t_5234), .d(t_9077), .cin(t_9079), .o(t_9086), .co(t_9087), .cout(t_9088));
compressor_4_2 u2_3128(.a(t_5196), .b(t_5193), .c(t_5190), .d(t_5187), .cin(t_5243), .o(t_9089), .co(t_9090), .cout(t_9091));
compressor_4_2 u2_3129(.a(t_5211), .b(t_5208), .c(t_5205), .d(t_5202), .cin(t_5199), .o(t_9092), .co(t_9093), .cout(t_9094));
compressor_4_2 u2_3130(.a(t_5249), .b(t_5246), .c(s_180_38), .d(t_9082), .cin(t_9085), .o(t_9095), .co(t_9096), .cout(t_9097));
compressor_4_2 u2_3131(.a(t_5258), .b(t_5255), .c(t_5252), .d(t_9088), .cin(t_9091), .o(t_9098), .co(t_9099), .cout(t_9100));
compressor_4_2 u2_3132(.a(t_5270), .b(t_5267), .c(t_5264), .d(t_5261), .cin(t_9094), .o(t_9101), .co(t_9102), .cout(t_9103));
compressor_4_2 u2_3133(.a(t_5226), .b(t_5223), .c(t_5220), .d(t_5217), .cin(t_5273), .o(t_9104), .co(t_9105), .cout(t_9106));
compressor_4_2 u2_3134(.a(t_5241), .b(t_5238), .c(t_5235), .d(t_5232), .cin(t_5229), .o(t_9107), .co(t_9108), .cout(t_9109));
compressor_4_2 u2_3135(.a(t_5278), .b(t_5275), .c(s_181_38), .d(t_9097), .cin(t_9100), .o(t_9110), .co(t_9111), .cout(t_9112));
compressor_4_2 u2_3136(.a(t_5287), .b(t_5284), .c(t_5281), .d(t_9103), .cin(t_9106), .o(t_9113), .co(t_9114), .cout(t_9115));
compressor_4_2 u2_3137(.a(t_5299), .b(t_5296), .c(t_5293), .d(t_5290), .cin(t_9109), .o(t_9116), .co(t_9117), .cout(t_9118));
compressor_4_2 u2_3138(.a(t_5256), .b(t_5253), .c(t_5250), .d(t_5247), .cin(t_5302), .o(t_9119), .co(t_9120), .cout(t_9121));
compressor_4_2 u2_3139(.a(t_5271), .b(t_5268), .c(t_5265), .d(t_5262), .cin(t_5259), .o(t_9122), .co(t_9123), .cout(t_9124));
compressor_4_2 u2_3140(.a(t_5310), .b(t_5307), .c(t_5304), .d(t_9112), .cin(t_9115), .o(t_9125), .co(t_9126), .cout(t_9127));
compressor_4_2 u2_3141(.a(t_5319), .b(t_5316), .c(t_5313), .d(t_9118), .cin(t_9121), .o(t_9128), .co(t_9129), .cout(t_9130));
compressor_4_2 u2_3142(.a(t_5331), .b(t_5328), .c(t_5325), .d(t_5322), .cin(t_9124), .o(t_9131), .co(t_9132), .cout(t_9133));
compressor_4_2 u2_3143(.a(t_5288), .b(t_5285), .c(t_5282), .d(t_5279), .cin(t_5276), .o(t_9134), .co(t_9135), .cout(t_9136));
compressor_3_2 u1_3144(.a(t_5297), .b(t_5294), .cin(t_5291), .o(t_9137), .cout(t_9138));
compressor_4_2 u2_3145(.a(t_5339), .b(t_5336), .c(t_5333), .d(t_9127), .cin(t_9130), .o(t_9139), .co(t_9140), .cout(t_9141));
compressor_4_2 u2_3146(.a(t_5348), .b(t_5345), .c(t_5342), .d(t_9133), .cin(t_9136), .o(t_9142), .co(t_9143), .cout(t_9144));
compressor_4_2 u2_3147(.a(t_5360), .b(t_5357), .c(t_5354), .d(t_5351), .cin(t_9138), .o(t_9145), .co(t_9146), .cout(t_9147));
compressor_4_2 u2_3148(.a(t_5317), .b(t_5314), .c(t_5311), .d(t_5308), .cin(t_5305), .o(t_9148), .co(t_9149), .cout(t_9150));
compressor_3_2 u1_3149(.a(t_5326), .b(t_5323), .cin(t_5320), .o(t_9151), .cout(t_9152));
compressor_4_2 u2_3150(.a(t_5368), .b(t_5365), .c(t_5362), .d(t_9141), .cin(t_9144), .o(t_9153), .co(t_9154), .cout(t_9155));
compressor_4_2 u2_3151(.a(t_5377), .b(t_5374), .c(t_5371), .d(t_9147), .cin(t_9150), .o(t_9156), .co(t_9157), .cout(t_9158));
compressor_4_2 u2_3152(.a(t_5389), .b(t_5386), .c(t_5383), .d(t_5380), .cin(t_9152), .o(t_9159), .co(t_9160), .cout(t_9161));
compressor_4_2 u2_3153(.a(t_5346), .b(t_5343), .c(t_5340), .d(t_5337), .cin(t_5334), .o(t_9162), .co(t_9163), .cout(t_9164));
compressor_3_2 u1_3154(.a(t_5355), .b(t_5352), .cin(t_5349), .o(t_9165), .cout(t_9166));
compressor_4_2 u2_3155(.a(t_5397), .b(t_5394), .c(t_5391), .d(t_9155), .cin(t_9158), .o(t_9167), .co(t_9168), .cout(t_9169));
compressor_4_2 u2_3156(.a(t_5406), .b(t_5403), .c(t_5400), .d(t_9161), .cin(t_9164), .o(t_9170), .co(t_9171), .cout(t_9172));
compressor_4_2 u2_3157(.a(t_5418), .b(t_5415), .c(t_5412), .d(t_5409), .cin(t_9166), .o(t_9173), .co(t_9174), .cout(t_9175));
compressor_4_2 u2_3158(.a(t_5375), .b(t_5372), .c(t_5369), .d(t_5366), .cin(t_5363), .o(t_9176), .co(t_9177), .cout(t_9178));
compressor_3_2 u1_3159(.a(t_5384), .b(t_5381), .cin(t_5378), .o(t_9179), .cout(t_9180));
compressor_4_2 u2_3160(.a(t_5423), .b(t_5420), .c(s_186_35), .d(t_9169), .cin(t_9172), .o(t_9181), .co(t_9182), .cout(t_9183));
compressor_4_2 u2_3161(.a(t_5432), .b(t_5429), .c(t_5426), .d(t_9175), .cin(t_9178), .o(t_9184), .co(t_9185), .cout(t_9186));
compressor_4_2 u2_3162(.a(t_5444), .b(t_5441), .c(t_5438), .d(t_5435), .cin(t_9180), .o(t_9187), .co(t_9188), .cout(t_9189));
compressor_4_2 u2_3163(.a(t_5404), .b(t_5401), .c(t_5398), .d(t_5395), .cin(t_5392), .o(t_9190), .co(t_9191), .cout(t_9192));
compressor_3_2 u1_3164(.a(t_5413), .b(t_5410), .cin(t_5407), .o(t_9193), .cout(t_9194));
compressor_4_2 u2_3165(.a(t_5453), .b(t_5450), .c(t_5447), .d(t_9183), .cin(t_9186), .o(t_9195), .co(t_9196), .cout(t_9197));
compressor_4_2 u2_3166(.a(t_5462), .b(t_5459), .c(t_5456), .d(t_9189), .cin(t_9192), .o(t_9198), .co(t_9199), .cout(t_9200));
compressor_4_2 u2_3167(.a(t_5421), .b(t_5471), .c(t_5468), .d(t_5465), .cin(t_9194), .o(t_9201), .co(t_9202), .cout(t_9203));
compressor_4_2 u2_3168(.a(t_5436), .b(t_5433), .c(t_5430), .d(t_5427), .cin(t_5424), .o(t_9204), .co(t_9205), .cout(t_9206));
compressor_3_2 u1_3169(.a(t_5445), .b(t_5442), .cin(t_5439), .o(t_9207), .cout(t_9208));
compressor_4_2 u2_3170(.a(t_5477), .b(t_5474), .c(s_188_34), .d(t_9197), .cin(t_9200), .o(t_9209), .co(t_9210), .cout(t_9211));
compressor_4_2 u2_3171(.a(t_5486), .b(t_5483), .c(t_5480), .d(t_9203), .cin(t_9206), .o(t_9212), .co(t_9213), .cout(t_9214));
compressor_4_2 u2_3172(.a(t_5498), .b(t_5495), .c(t_5492), .d(t_5489), .cin(t_9208), .o(t_9215), .co(t_9216), .cout(t_9217));
compressor_4_2 u2_3173(.a(t_5460), .b(t_5457), .c(t_5454), .d(t_5451), .cin(t_5448), .o(t_9218), .co(t_9219), .cout(t_9220));
compressor_3_2 u1_3174(.a(t_5469), .b(t_5466), .cin(t_5463), .o(t_9221), .cout(t_9222));
compressor_4_2 u2_3175(.a(t_5503), .b(t_5500), .c(s_189_34), .d(t_9211), .cin(t_9214), .o(t_9223), .co(t_9224), .cout(t_9225));
compressor_4_2 u2_3176(.a(t_5512), .b(t_5509), .c(t_5506), .d(t_9217), .cin(t_9220), .o(t_9226), .co(t_9227), .cout(t_9228));
compressor_4_2 u2_3177(.a(t_5524), .b(t_5521), .c(t_5518), .d(t_5515), .cin(t_9222), .o(t_9229), .co(t_9230), .cout(t_9231));
compressor_4_2 u2_3178(.a(t_5487), .b(t_5484), .c(t_5481), .d(t_5478), .cin(t_5475), .o(t_9232), .co(t_9233), .cout(t_9234));
compressor_3_2 u1_3179(.a(t_5496), .b(t_5493), .cin(t_5490), .o(t_9235), .cout(t_9236));
compressor_4_2 u2_3180(.a(t_5532), .b(t_5529), .c(t_5526), .d(t_9225), .cin(t_9228), .o(t_9237), .co(t_9238), .cout(t_9239));
compressor_4_2 u2_3181(.a(t_5541), .b(t_5538), .c(t_5535), .d(t_9231), .cin(t_9234), .o(t_9240), .co(t_9241), .cout(t_9242));
compressor_4_2 u2_3182(.a(t_5501), .b(t_5550), .c(t_5547), .d(t_5544), .cin(t_9236), .o(t_9243), .co(t_9244), .cout(t_9245));
compressor_4_2 u2_3183(.a(t_5516), .b(t_5513), .c(t_5510), .d(t_5507), .cin(t_5504), .o(t_9246), .co(t_9247), .cout(t_9248));
half_adder u0_3184(.a(t_5522), .b(t_5519), .o(t_9249), .cout(t_9250));
compressor_4_2 u2_3185(.a(t_5558), .b(t_5555), .c(t_5552), .d(t_9239), .cin(t_9242), .o(t_9251), .co(t_9252), .cout(t_9253));
compressor_4_2 u2_3186(.a(t_5567), .b(t_5564), .c(t_5561), .d(t_9245), .cin(t_9248), .o(t_9254), .co(t_9255), .cout(t_9256));
compressor_4_2 u2_3187(.a(t_5527), .b(t_5576), .c(t_5573), .d(t_5570), .cin(t_9250), .o(t_9257), .co(t_9258), .cout(t_9259));
compressor_4_2 u2_3188(.a(t_5542), .b(t_5539), .c(t_5536), .d(t_5533), .cin(t_5530), .o(t_9260), .co(t_9261), .cout(t_9262));
half_adder u0_3189(.a(t_5548), .b(t_5545), .o(t_9263), .cout(t_9264));
compressor_4_2 u2_3190(.a(t_5584), .b(t_5581), .c(t_5578), .d(t_9253), .cin(t_9256), .o(t_9265), .co(t_9266), .cout(t_9267));
compressor_4_2 u2_3191(.a(t_5593), .b(t_5590), .c(t_5587), .d(t_9259), .cin(t_9262), .o(t_9268), .co(t_9269), .cout(t_9270));
compressor_4_2 u2_3192(.a(t_5553), .b(t_5602), .c(t_5599), .d(t_5596), .cin(t_9264), .o(t_9271), .co(t_9272), .cout(t_9273));
compressor_4_2 u2_3193(.a(t_5568), .b(t_5565), .c(t_5562), .d(t_5559), .cin(t_5556), .o(t_9274), .co(t_9275), .cout(t_9276));
half_adder u0_3194(.a(t_5574), .b(t_5571), .o(t_9277), .cout(t_9278));
compressor_4_2 u2_3195(.a(t_5610), .b(t_5607), .c(t_5604), .d(t_9267), .cin(t_9270), .o(t_9279), .co(t_9280), .cout(t_9281));
compressor_4_2 u2_3196(.a(t_5619), .b(t_5616), .c(t_5613), .d(t_9273), .cin(t_9276), .o(t_9282), .co(t_9283), .cout(t_9284));
compressor_4_2 u2_3197(.a(t_5579), .b(t_5628), .c(t_5625), .d(t_5622), .cin(t_9278), .o(t_9285), .co(t_9286), .cout(t_9287));
compressor_4_2 u2_3198(.a(t_5594), .b(t_5591), .c(t_5588), .d(t_5585), .cin(t_5582), .o(t_9288), .co(t_9289), .cout(t_9290));
half_adder u0_3199(.a(t_5600), .b(t_5597), .o(t_9291), .cout(t_9292));
compressor_4_2 u2_3200(.a(t_5633), .b(t_5630), .c(s_194_31), .d(t_9281), .cin(t_9284), .o(t_9293), .co(t_9294), .cout(t_9295));
compressor_4_2 u2_3201(.a(t_5642), .b(t_5639), .c(t_5636), .d(t_9287), .cin(t_9290), .o(t_9296), .co(t_9297), .cout(t_9298));
compressor_4_2 u2_3202(.a(t_5605), .b(t_5651), .c(t_5648), .d(t_5645), .cin(t_9292), .o(t_9299), .co(t_9300), .cout(t_9301));
compressor_4_2 u2_3203(.a(t_5620), .b(t_5617), .c(t_5614), .d(t_5611), .cin(t_5608), .o(t_9302), .co(t_9303), .cout(t_9304));
half_adder u0_3204(.a(t_5626), .b(t_5623), .o(t_9305), .cout(t_9306));
compressor_4_2 u2_3205(.a(t_5660), .b(t_5657), .c(t_5654), .d(t_9295), .cin(t_9298), .o(t_9307), .co(t_9308), .cout(t_9309));
compressor_4_2 u2_3206(.a(t_5669), .b(t_5666), .c(t_5663), .d(t_9301), .cin(t_9304), .o(t_9310), .co(t_9311), .cout(t_9312));
compressor_4_2 u2_3207(.a(t_5634), .b(t_5631), .c(t_5675), .d(t_5672), .cin(t_9306), .o(t_9313), .co(t_9314), .cout(t_9315));
compressor_4_2 u2_3208(.a(t_5649), .b(t_5646), .c(t_5643), .d(t_5640), .cin(t_5637), .o(t_9316), .co(t_9317), .cout(t_9318));
compressor_4_2 u2_3209(.a(t_5681), .b(t_5678), .c(s_196_30), .d(t_9309), .cin(t_9312), .o(t_9319), .co(t_9320), .cout(t_9321));
compressor_4_2 u2_3210(.a(t_5690), .b(t_5687), .c(t_5684), .d(t_9315), .cin(t_9318), .o(t_9322), .co(t_9323), .cout(t_9324));
compressor_4_2 u2_3211(.a(t_5658), .b(t_5655), .c(t_5699), .d(t_5696), .cin(t_5693), .o(t_9325), .co(t_9326), .cout(t_9327));
compressor_4_2 u2_3212(.a(t_5673), .b(t_5670), .c(t_5667), .d(t_5664), .cin(t_5661), .o(t_9328), .co(t_9329), .cout(t_9330));
compressor_4_2 u2_3213(.a(t_5704), .b(t_5701), .c(s_197_30), .d(t_9321), .cin(t_9324), .o(t_9331), .co(t_9332), .cout(t_9333));
compressor_4_2 u2_3214(.a(t_5713), .b(t_5710), .c(t_5707), .d(t_9327), .cin(t_9330), .o(t_9334), .co(t_9335), .cout(t_9336));
compressor_4_2 u2_3215(.a(t_5682), .b(t_5679), .c(t_5722), .d(t_5719), .cin(t_5716), .o(t_9337), .co(t_9338), .cout(t_9339));
compressor_4_2 u2_3216(.a(t_5697), .b(t_5694), .c(t_5691), .d(t_5688), .cin(t_5685), .o(t_9340), .co(t_9341), .cout(t_9342));
compressor_4_2 u2_3217(.a(t_5730), .b(t_5727), .c(t_5724), .d(t_9333), .cin(t_9336), .o(t_9343), .co(t_9344), .cout(t_9345));
compressor_4_2 u2_3218(.a(t_5739), .b(t_5736), .c(t_5733), .d(t_9339), .cin(t_9342), .o(t_9346), .co(t_9347), .cout(t_9348));
compressor_4_2 u2_3219(.a(t_5708), .b(t_5705), .c(t_5702), .d(t_5745), .cin(t_5742), .o(t_9349), .co(t_9350), .cout(t_9351));
compressor_3_2 u1_3220(.a(t_5717), .b(t_5714), .cin(t_5711), .o(t_9352), .cout(t_9353));
compressor_4_2 u2_3221(.a(t_5753), .b(t_5750), .c(t_5747), .d(t_9345), .cin(t_9348), .o(t_9354), .co(t_9355), .cout(t_9356));
compressor_4_2 u2_3222(.a(t_5762), .b(t_5759), .c(t_5756), .d(t_9351), .cin(t_9353), .o(t_9357), .co(t_9358), .cout(t_9359));
compressor_4_2 u2_3223(.a(t_5731), .b(t_5728), .c(t_5725), .d(t_5768), .cin(t_5765), .o(t_9360), .co(t_9361), .cout(t_9362));
compressor_3_2 u1_3224(.a(t_5740), .b(t_5737), .cin(t_5734), .o(t_9363), .cout(t_9364));
compressor_4_2 u2_3225(.a(t_5776), .b(t_5773), .c(t_5770), .d(t_9356), .cin(t_9359), .o(t_9365), .co(t_9366), .cout(t_9367));
compressor_4_2 u2_3226(.a(t_5785), .b(t_5782), .c(t_5779), .d(t_9362), .cin(t_9364), .o(t_9368), .co(t_9369), .cout(t_9370));
compressor_4_2 u2_3227(.a(t_5754), .b(t_5751), .c(t_5748), .d(t_5791), .cin(t_5788), .o(t_9371), .co(t_9372), .cout(t_9373));
compressor_3_2 u1_3228(.a(t_5763), .b(t_5760), .cin(t_5757), .o(t_9374), .cout(t_9375));
compressor_4_2 u2_3229(.a(t_5799), .b(t_5796), .c(t_5793), .d(t_9367), .cin(t_9370), .o(t_9376), .co(t_9377), .cout(t_9378));
compressor_4_2 u2_3230(.a(t_5808), .b(t_5805), .c(t_5802), .d(t_9373), .cin(t_9375), .o(t_9379), .co(t_9380), .cout(t_9381));
compressor_4_2 u2_3231(.a(t_5777), .b(t_5774), .c(t_5771), .d(t_5814), .cin(t_5811), .o(t_9382), .co(t_9383), .cout(t_9384));
compressor_3_2 u1_3232(.a(t_5786), .b(t_5783), .cin(t_5780), .o(t_9385), .cout(t_9386));
compressor_4_2 u2_3233(.a(t_5819), .b(t_5816), .c(s_202_27), .d(t_9378), .cin(t_9381), .o(t_9387), .co(t_9388), .cout(t_9389));
compressor_4_2 u2_3234(.a(t_5828), .b(t_5825), .c(t_5822), .d(t_9384), .cin(t_9386), .o(t_9390), .co(t_9391), .cout(t_9392));
compressor_4_2 u2_3235(.a(t_5800), .b(t_5797), .c(t_5794), .d(t_5834), .cin(t_5831), .o(t_9393), .co(t_9394), .cout(t_9395));
compressor_3_2 u1_3236(.a(t_5809), .b(t_5806), .cin(t_5803), .o(t_9396), .cout(t_9397));
compressor_4_2 u2_3237(.a(t_5843), .b(t_5840), .c(t_5837), .d(t_9389), .cin(t_9392), .o(t_9398), .co(t_9399), .cout(t_9400));
compressor_4_2 u2_3238(.a(t_5852), .b(t_5849), .c(t_5846), .d(t_9395), .cin(t_9397), .o(t_9401), .co(t_9402), .cout(t_9403));
compressor_4_2 u2_3239(.a(t_5826), .b(t_5823), .c(t_5820), .d(t_5817), .cin(t_5855), .o(t_9404), .co(t_9405), .cout(t_9406));
compressor_3_2 u1_3240(.a(t_5835), .b(t_5832), .cin(t_5829), .o(t_9407), .cout(t_9408));
compressor_4_2 u2_3241(.a(t_5861), .b(t_5858), .c(s_204_26), .d(t_9400), .cin(t_9403), .o(t_9409), .co(t_9410), .cout(t_9411));
compressor_4_2 u2_3242(.a(t_5870), .b(t_5867), .c(t_5864), .d(t_9406), .cin(t_9408), .o(t_9412), .co(t_9413), .cout(t_9414));
compressor_4_2 u2_3243(.a(t_5844), .b(t_5841), .c(t_5838), .d(t_5876), .cin(t_5873), .o(t_9415), .co(t_9416), .cout(t_9417));
compressor_3_2 u1_3244(.a(t_5853), .b(t_5850), .cin(t_5847), .o(t_9418), .cout(t_9419));
compressor_4_2 u2_3245(.a(t_5881), .b(t_5878), .c(s_205_26), .d(t_9411), .cin(t_9414), .o(t_9420), .co(t_9421), .cout(t_9422));
compressor_4_2 u2_3246(.a(t_5890), .b(t_5887), .c(t_5884), .d(t_9417), .cin(t_9419), .o(t_9423), .co(t_9424), .cout(t_9425));
compressor_4_2 u2_3247(.a(t_5865), .b(t_5862), .c(t_5859), .d(t_5896), .cin(t_5893), .o(t_9426), .co(t_9427), .cout(t_9428));
compressor_3_2 u1_3248(.a(t_5874), .b(t_5871), .cin(t_5868), .o(t_9429), .cout(t_9430));
compressor_4_2 u2_3249(.a(t_5904), .b(t_5901), .c(t_5898), .d(t_9422), .cin(t_9425), .o(t_9431), .co(t_9432), .cout(t_9433));
compressor_4_2 u2_3250(.a(t_5913), .b(t_5910), .c(t_5907), .d(t_9428), .cin(t_9430), .o(t_9434), .co(t_9435), .cout(t_9436));
compressor_4_2 u2_3251(.a(t_5888), .b(t_5885), .c(t_5882), .d(t_5879), .cin(t_5916), .o(t_9437), .co(t_9438), .cout(t_9439));
half_adder u0_3252(.a(t_5894), .b(t_5891), .o(t_9440), .cout(t_9441));
compressor_4_2 u2_3253(.a(t_5924), .b(t_5921), .c(t_5918), .d(t_9433), .cin(t_9436), .o(t_9442), .co(t_9443), .cout(t_9444));
compressor_4_2 u2_3254(.a(t_5933), .b(t_5930), .c(t_5927), .d(t_9439), .cin(t_9441), .o(t_9445), .co(t_9446), .cout(t_9447));
compressor_4_2 u2_3255(.a(t_5908), .b(t_5905), .c(t_5902), .d(t_5899), .cin(t_5936), .o(t_9448), .co(t_9449), .cout(t_9450));
half_adder u0_3256(.a(t_5914), .b(t_5911), .o(t_9451), .cout(t_9452));
compressor_4_2 u2_3257(.a(t_5944), .b(t_5941), .c(t_5938), .d(t_9444), .cin(t_9447), .o(t_9453), .co(t_9454), .cout(t_9455));
compressor_4_2 u2_3258(.a(t_5953), .b(t_5950), .c(t_5947), .d(t_9450), .cin(t_9452), .o(t_9456), .co(t_9457), .cout(t_9458));
compressor_4_2 u2_3259(.a(t_5928), .b(t_5925), .c(t_5922), .d(t_5919), .cin(t_5956), .o(t_9459), .co(t_9460), .cout(t_9461));
half_adder u0_3260(.a(t_5934), .b(t_5931), .o(t_9462), .cout(t_9463));
compressor_4_2 u2_3261(.a(t_5964), .b(t_5961), .c(t_5958), .d(t_9455), .cin(t_9458), .o(t_9464), .co(t_9465), .cout(t_9466));
compressor_4_2 u2_3262(.a(t_5973), .b(t_5970), .c(t_5967), .d(t_9461), .cin(t_9463), .o(t_9467), .co(t_9468), .cout(t_9469));
compressor_4_2 u2_3263(.a(t_5948), .b(t_5945), .c(t_5942), .d(t_5939), .cin(t_5976), .o(t_9470), .co(t_9471), .cout(t_9472));
half_adder u0_3264(.a(t_5954), .b(t_5951), .o(t_9473), .cout(t_9474));
compressor_4_2 u2_3265(.a(t_5981), .b(t_5978), .c(s_210_23), .d(t_9466), .cin(t_9469), .o(t_9475), .co(t_9476), .cout(t_9477));
compressor_4_2 u2_3266(.a(t_5990), .b(t_5987), .c(t_5984), .d(t_9472), .cin(t_9474), .o(t_9478), .co(t_9479), .cout(t_9480));
compressor_4_2 u2_3267(.a(t_5968), .b(t_5965), .c(t_5962), .d(t_5959), .cin(t_5993), .o(t_9481), .co(t_9482), .cout(t_9483));
half_adder u0_3268(.a(t_5974), .b(t_5971), .o(t_9484), .cout(t_9485));
compressor_4_2 u2_3269(.a(t_6002), .b(t_5999), .c(t_5996), .d(t_9477), .cin(t_9480), .o(t_9486), .co(t_9487), .cout(t_9488));
compressor_4_2 u2_3270(.a(t_6011), .b(t_6008), .c(t_6005), .d(t_9483), .cin(t_9485), .o(t_9489), .co(t_9490), .cout(t_9491));
compressor_4_2 u2_3271(.a(t_5991), .b(t_5988), .c(t_5985), .d(t_5982), .cin(t_5979), .o(t_9492), .co(t_9493), .cout(t_9494));
compressor_4_2 u2_3272(.a(t_6017), .b(t_6014), .c(s_212_22), .d(t_9488), .cin(t_9491), .o(t_9495), .co(t_9496), .cout(t_9497));
compressor_4_2 u2_3273(.a(t_6029), .b(t_6026), .c(t_6023), .d(t_6020), .cin(t_9494), .o(t_9498), .co(t_9499), .cout(t_9500));
compressor_4_2 u2_3274(.a(t_6009), .b(t_6006), .c(t_6003), .d(t_6000), .cin(t_5997), .o(t_9501), .co(t_9502), .cout(t_9503));
compressor_4_2 u2_3275(.a(t_6034), .b(t_6031), .c(s_213_22), .d(t_9497), .cin(t_9500), .o(t_9504), .co(t_9505), .cout(t_9506));
compressor_4_2 u2_3276(.a(t_6046), .b(t_6043), .c(t_6040), .d(t_6037), .cin(t_9503), .o(t_9507), .co(t_9508), .cout(t_9509));
compressor_4_2 u2_3277(.a(t_6027), .b(t_6024), .c(t_6021), .d(t_6018), .cin(t_6015), .o(t_9510), .co(t_9511), .cout(t_9512));
compressor_4_2 u2_3278(.a(t_6054), .b(t_6051), .c(t_6048), .d(t_9506), .cin(t_9509), .o(t_9513), .co(t_9514), .cout(t_9515));
compressor_4_2 u2_3279(.a(t_6032), .b(t_6063), .c(t_6060), .d(t_6057), .cin(t_9512), .o(t_9516), .co(t_9517), .cout(t_9518));
compressor_3_2 u1_3280(.a(t_6041), .b(t_6038), .cin(t_6035), .o(t_9519), .cout(t_9520));
compressor_4_2 u2_3281(.a(t_6071), .b(t_6068), .c(t_6065), .d(t_9515), .cin(t_9518), .o(t_9521), .co(t_9522), .cout(t_9523));
compressor_4_2 u2_3282(.a(t_6049), .b(t_6080), .c(t_6077), .d(t_6074), .cin(t_9520), .o(t_9524), .co(t_9525), .cout(t_9526));
compressor_3_2 u1_3283(.a(t_6058), .b(t_6055), .cin(t_6052), .o(t_9527), .cout(t_9528));
compressor_4_2 u2_3284(.a(t_6088), .b(t_6085), .c(t_6082), .d(t_9523), .cin(t_9526), .o(t_9529), .co(t_9530), .cout(t_9531));
compressor_4_2 u2_3285(.a(t_6066), .b(t_6097), .c(t_6094), .d(t_6091), .cin(t_9528), .o(t_9532), .co(t_9533), .cout(t_9534));
compressor_3_2 u1_3286(.a(t_6075), .b(t_6072), .cin(t_6069), .o(t_9535), .cout(t_9536));
compressor_4_2 u2_3287(.a(t_6105), .b(t_6102), .c(t_6099), .d(t_9531), .cin(t_9534), .o(t_9537), .co(t_9538), .cout(t_9539));
compressor_4_2 u2_3288(.a(t_6083), .b(t_6114), .c(t_6111), .d(t_6108), .cin(t_9536), .o(t_9540), .co(t_9541), .cout(t_9542));
compressor_3_2 u1_3289(.a(t_6092), .b(t_6089), .cin(t_6086), .o(t_9543), .cout(t_9544));
compressor_4_2 u2_3290(.a(t_6119), .b(t_6116), .c(s_218_19), .d(t_9539), .cin(t_9542), .o(t_9545), .co(t_9546), .cout(t_9547));
compressor_4_2 u2_3291(.a(t_6100), .b(t_6128), .c(t_6125), .d(t_6122), .cin(t_9544), .o(t_9548), .co(t_9549), .cout(t_9550));
compressor_3_2 u1_3292(.a(t_6109), .b(t_6106), .cin(t_6103), .o(t_9551), .cout(t_9552));
compressor_4_2 u2_3293(.a(t_6137), .b(t_6134), .c(t_6131), .d(t_9547), .cin(t_9550), .o(t_9553), .co(t_9554), .cout(t_9555));
compressor_4_2 u2_3294(.a(t_6120), .b(t_6117), .c(t_6143), .d(t_6140), .cin(t_9552), .o(t_9556), .co(t_9557), .cout(t_9558));
compressor_3_2 u1_3295(.a(t_6129), .b(t_6126), .cin(t_6123), .o(t_9559), .cout(t_9560));
compressor_4_2 u2_3296(.a(t_6149), .b(t_6146), .c(s_220_18), .d(t_9555), .cin(t_9558), .o(t_9561), .co(t_9562), .cout(t_9563));
compressor_4_2 u2_3297(.a(t_6132), .b(t_6158), .c(t_6155), .d(t_6152), .cin(t_9560), .o(t_9564), .co(t_9565), .cout(t_9566));
compressor_3_2 u1_3298(.a(t_6141), .b(t_6138), .cin(t_6135), .o(t_9567), .cout(t_9568));
compressor_4_2 u2_3299(.a(t_6163), .b(t_6160), .c(s_221_18), .d(t_9563), .cin(t_9566), .o(t_9569), .co(t_9570), .cout(t_9571));
compressor_4_2 u2_3300(.a(t_6147), .b(t_6172), .c(t_6169), .d(t_6166), .cin(t_9568), .o(t_9572), .co(t_9573), .cout(t_9574));
compressor_3_2 u1_3301(.a(t_6156), .b(t_6153), .cin(t_6150), .o(t_9575), .cout(t_9576));
compressor_4_2 u2_3302(.a(t_6180), .b(t_6177), .c(t_6174), .d(t_9571), .cin(t_9574), .o(t_9577), .co(t_9578), .cout(t_9579));
compressor_4_2 u2_3303(.a(t_6164), .b(t_6161), .c(t_6186), .d(t_6183), .cin(t_9576), .o(t_9580), .co(t_9581), .cout(t_9582));
half_adder u0_3304(.a(t_6170), .b(t_6167), .o(t_9583), .cout(t_9584));
compressor_4_2 u2_3305(.a(t_6194), .b(t_6191), .c(t_6188), .d(t_9579), .cin(t_9582), .o(t_9585), .co(t_9586), .cout(t_9587));
compressor_4_2 u2_3306(.a(t_6178), .b(t_6175), .c(t_6200), .d(t_6197), .cin(t_9584), .o(t_9588), .co(t_9589), .cout(t_9590));
half_adder u0_3307(.a(t_6184), .b(t_6181), .o(t_9591), .cout(t_9592));
compressor_4_2 u2_3308(.a(t_6208), .b(t_6205), .c(t_6202), .d(t_9587), .cin(t_9590), .o(t_9593), .co(t_9594), .cout(t_9595));
compressor_4_2 u2_3309(.a(t_6192), .b(t_6189), .c(t_6214), .d(t_6211), .cin(t_9592), .o(t_9596), .co(t_9597), .cout(t_9598));
half_adder u0_3310(.a(t_6198), .b(t_6195), .o(t_9599), .cout(t_9600));
compressor_4_2 u2_3311(.a(t_6222), .b(t_6219), .c(t_6216), .d(t_9595), .cin(t_9598), .o(t_9601), .co(t_9602), .cout(t_9603));
compressor_4_2 u2_3312(.a(t_6206), .b(t_6203), .c(t_6228), .d(t_6225), .cin(t_9600), .o(t_9604), .co(t_9605), .cout(t_9606));
half_adder u0_3313(.a(t_6212), .b(t_6209), .o(t_9607), .cout(t_9608));
compressor_4_2 u2_3314(.a(t_6233), .b(t_6230), .c(s_226_15), .d(t_9603), .cin(t_9606), .o(t_9609), .co(t_9610), .cout(t_9611));
compressor_4_2 u2_3315(.a(t_6220), .b(t_6217), .c(t_6239), .d(t_6236), .cin(t_9608), .o(t_9612), .co(t_9613), .cout(t_9614));
half_adder u0_3316(.a(t_6226), .b(t_6223), .o(t_9615), .cout(t_9616));
compressor_4_2 u2_3317(.a(t_6248), .b(t_6245), .c(t_6242), .d(t_9611), .cin(t_9614), .o(t_9617), .co(t_9618), .cout(t_9619));
compressor_4_2 u2_3318(.a(t_6237), .b(t_6234), .c(t_6231), .d(t_6251), .cin(t_9616), .o(t_9620), .co(t_9621), .cout(t_9622));
compressor_4_2 u2_3319(.a(t_6257), .b(t_6254), .c(s_228_14), .d(t_9619), .cin(t_9622), .o(t_9623), .co(t_9624), .cout(t_9625));
compressor_4_2 u2_3320(.a(t_6249), .b(t_6246), .c(t_6243), .d(t_6263), .cin(t_6260), .o(t_9626), .co(t_9627), .cout(t_9628));
compressor_4_2 u2_3321(.a(t_6268), .b(t_6265), .c(s_229_14), .d(t_9625), .cin(t_9628), .o(t_9629), .co(t_9630), .cout(t_9631));
compressor_4_2 u2_3322(.a(t_6261), .b(t_6258), .c(t_6255), .d(t_6274), .cin(t_6271), .o(t_9632), .co(t_9633), .cout(t_9634));
compressor_4_2 u2_3323(.a(t_6282), .b(t_6279), .c(t_6276), .d(t_9631), .cin(t_9634), .o(t_9635), .co(t_9636), .cout(t_9637));
compressor_3_2 u1_3324(.a(t_6269), .b(t_6266), .cin(t_6285), .o(t_9638), .cout(t_9639));
compressor_4_2 u2_3325(.a(t_6293), .b(t_6290), .c(t_6287), .d(t_9637), .cin(t_9639), .o(t_9640), .co(t_9641), .cout(t_9642));
compressor_3_2 u1_3326(.a(t_6280), .b(t_6277), .cin(t_6296), .o(t_9643), .cout(t_9644));
compressor_4_2 u2_3327(.a(t_6304), .b(t_6301), .c(t_6298), .d(t_9642), .cin(t_9644), .o(t_9645), .co(t_9646), .cout(t_9647));
compressor_3_2 u1_3328(.a(t_6291), .b(t_6288), .cin(t_6307), .o(t_9648), .cout(t_9649));
compressor_4_2 u2_3329(.a(t_6315), .b(t_6312), .c(t_6309), .d(t_9647), .cin(t_9649), .o(t_9650), .co(t_9651), .cout(t_9652));
compressor_3_2 u1_3330(.a(t_6302), .b(t_6299), .cin(t_6318), .o(t_9653), .cout(t_9654));
compressor_4_2 u2_3331(.a(t_6323), .b(t_6320), .c(s_234_11), .d(t_9652), .cin(t_9654), .o(t_9655), .co(t_9656), .cout(t_9657));
compressor_3_2 u1_3332(.a(t_6313), .b(t_6310), .cin(t_6326), .o(t_9658), .cout(t_9659));
compressor_4_2 u2_3333(.a(t_6335), .b(t_6332), .c(t_6329), .d(t_9657), .cin(t_9659), .o(t_9660), .co(t_9661), .cout(t_9662));
compressor_3_2 u1_3334(.a(t_6327), .b(t_6324), .cin(t_6321), .o(t_9663), .cout(t_9664));
compressor_4_2 u2_3335(.a(t_6341), .b(t_6338), .c(s_236_10), .d(t_9662), .cin(t_9664), .o(t_9665), .co(t_9666), .cout(t_9667));
compressor_3_2 u1_3336(.a(t_6333), .b(t_6330), .cin(t_6344), .o(t_9668), .cout(t_9669));
compressor_4_2 u2_3337(.a(t_6349), .b(t_6346), .c(s_237_10), .d(t_9667), .cin(t_9669), .o(t_9670), .co(t_9671), .cout(t_9672));
compressor_3_2 u1_3338(.a(t_6342), .b(t_6339), .cin(t_6352), .o(t_9673), .cout(t_9674));
compressor_4_2 u2_3339(.a(t_6360), .b(t_6357), .c(t_6354), .d(t_9672), .cin(t_9674), .o(t_9675), .co(t_9676), .cout(t_9677));
half_adder u0_3340(.a(t_6350), .b(t_6347), .o(t_9678), .cout(t_9679));
compressor_4_2 u2_3341(.a(t_6368), .b(t_6365), .c(t_6362), .d(t_9677), .cin(t_9679), .o(t_9680), .co(t_9681), .cout(t_9682));
half_adder u0_3342(.a(t_6358), .b(t_6355), .o(t_9683), .cout(t_9684));
compressor_4_2 u2_3343(.a(t_6376), .b(t_6373), .c(t_6370), .d(t_9682), .cin(t_9684), .o(t_9685), .co(t_9686), .cout(t_9687));
half_adder u0_3344(.a(t_6366), .b(t_6363), .o(t_9688), .cout(t_9689));
compressor_4_2 u2_3345(.a(t_6384), .b(t_6381), .c(t_6378), .d(t_9687), .cin(t_9689), .o(t_9690), .co(t_9691), .cout(t_9692));
half_adder u0_3346(.a(t_6374), .b(t_6371), .o(t_9693), .cout(t_9694));
compressor_4_2 u2_3347(.a(t_6389), .b(t_6386), .c(s_242_7), .d(t_9692), .cin(t_9694), .o(t_9695), .co(t_9696), .cout(t_9697));
half_adder u0_3348(.a(t_6382), .b(t_6379), .o(t_9698), .cout(t_9699));
compressor_4_2 u2_3349(.a(t_6387), .b(t_6395), .c(t_6392), .d(t_9697), .cin(t_9699), .o(t_9700), .co(t_9701), .cout(t_9702));
compressor_4_2 u2_3350(.a(t_6393), .b(t_6401), .c(t_6398), .d(s_244_6), .cin(t_9702), .o(t_9703), .co(t_9704), .cout(t_9705));
compressor_4_2 u2_3351(.a(t_6399), .b(t_6406), .c(t_6403), .d(s_245_6), .cin(t_9705), .o(t_9706), .co(t_9707), .cout(t_9708));
compressor_3_2 u1_3352(.a(t_6411), .b(t_6408), .cin(t_9708), .o(t_9709), .cout(t_9710));
compressor_3_2 u1_3353(.a(t_6409), .b(t_6416), .cin(t_6413), .o(t_9711), .cout(t_9712));
compressor_3_2 u1_3354(.a(t_6414), .b(t_6421), .cin(t_6418), .o(t_9713), .cout(t_9714));
compressor_3_2 u1_3355(.a(t_6419), .b(t_6426), .cin(t_6423), .o(t_9715), .cout(t_9716));
compressor_3_2 u1_3356(.a(t_6424), .b(t_6428), .cin(s_250_3), .o(t_9717), .cout(t_9718));
half_adder u0_3357(.a(t_6429), .b(t_6431), .o(t_9719), .cout(t_9720));
compressor_3_2 u1_3358(.a(t_6432), .b(t_6434), .cin(s_252_2), .o(t_9721), .cout(t_9722));
half_adder u0_3359(.a(t_6435), .b(t_6436), .o(t_9723), .cout(t_9724));
half_adder u0_3360(.a(t_6437), .b(t_6438), .o(t_9725), .cout(t_9726));
half_adder u0_3361(.a(t_6439), .b(t_6440), .o(t_9727), .cout());

/* u0_3362 Output nets */
wire t_9728,   t_9729;
/* u0_3363 Output nets */
wire t_9730,   t_9731;
/* u0_3364 Output nets */
wire t_9732,   t_9733;
/* u0_3365 Output nets */
wire t_9734,   t_9735;
/* u0_3366 Output nets */
wire t_9736,   t_9737;
/* u0_3367 Output nets */
wire t_9738,   t_9739;
/* u1_3368 Output nets */
wire t_9740,   t_9741;
/* u0_3369 Output nets */
wire t_9742,   t_9743;
/* u0_3370 Output nets */
wire t_9744,   t_9745;
/* u0_3371 Output nets */
wire t_9746,   t_9747;
/* u0_3372 Output nets */
wire t_9748,   t_9749;
/* u1_3373 Output nets */
wire t_9750,   t_9751;
/* u1_3374 Output nets */
wire t_9752,   t_9753;
/* u1_3375 Output nets */
wire t_9754,   t_9755;
/* u1_3376 Output nets */
wire t_9756,   t_9757;
/* u1_3377 Output nets */
wire t_9758,   t_9759;
/* u2_3378 Output nets */
wire t_9760,   t_9761,   t_9762;
/* u1_3379 Output nets */
wire t_9763,   t_9764;
/* u1_3380 Output nets */
wire t_9765,   t_9766;
/* u2_3381 Output nets */
wire t_9767,   t_9768,   t_9769;
/* u2_3382 Output nets */
wire t_9770,   t_9771,   t_9772;
/* u1_3383 Output nets */
wire t_9773,   t_9774;
/* u2_3384 Output nets */
wire t_9775,   t_9776,   t_9777;
/* u2_3385 Output nets */
wire t_9778,   t_9779,   t_9780;
/* u2_3386 Output nets */
wire t_9781,   t_9782,   t_9783;
/* u2_3387 Output nets */
wire t_9784,   t_9785,   t_9786;
/* u2_3388 Output nets */
wire t_9787,   t_9788,   t_9789;
/* u2_3389 Output nets */
wire t_9790,   t_9791,   t_9792;
/* u2_3390 Output nets */
wire t_9793,   t_9794,   t_9795;
/* u2_3391 Output nets */
wire t_9796,   t_9797,   t_9798;
/* u2_3392 Output nets */
wire t_9799,   t_9800,   t_9801;
/* u2_3393 Output nets */
wire t_9802,   t_9803,   t_9804;
/* u2_3394 Output nets */
wire t_9805,   t_9806,   t_9807;
/* u0_3395 Output nets */
wire t_9808,   t_9809;
/* u2_3396 Output nets */
wire t_9810,   t_9811,   t_9812;
/* u0_3397 Output nets */
wire t_9813,   t_9814;
/* u2_3398 Output nets */
wire t_9815,   t_9816,   t_9817;
/* u0_3399 Output nets */
wire t_9818,   t_9819;
/* u2_3400 Output nets */
wire t_9820,   t_9821,   t_9822;
/* u1_3401 Output nets */
wire t_9823,   t_9824;
/* u2_3402 Output nets */
wire t_9825,   t_9826,   t_9827;
/* u1_3403 Output nets */
wire t_9828,   t_9829;
/* u2_3404 Output nets */
wire t_9830,   t_9831,   t_9832;
/* u0_3405 Output nets */
wire t_9833,   t_9834;
/* u2_3406 Output nets */
wire t_9835,   t_9836,   t_9837;
/* u1_3407 Output nets */
wire t_9838,   t_9839;
/* u2_3408 Output nets */
wire t_9840,   t_9841,   t_9842;
/* u1_3409 Output nets */
wire t_9843,   t_9844;
/* u2_3410 Output nets */
wire t_9845,   t_9846,   t_9847;
/* u1_3411 Output nets */
wire t_9848,   t_9849;
/* u2_3412 Output nets */
wire t_9850,   t_9851,   t_9852;
/* u1_3413 Output nets */
wire t_9853,   t_9854;
/* u2_3414 Output nets */
wire t_9855,   t_9856,   t_9857;
/* u1_3415 Output nets */
wire t_9858,   t_9859;
/* u2_3416 Output nets */
wire t_9860,   t_9861,   t_9862;
/* u1_3417 Output nets */
wire t_9863,   t_9864;
/* u2_3418 Output nets */
wire t_9865,   t_9866,   t_9867;
/* u1_3419 Output nets */
wire t_9868,   t_9869;
/* u2_3420 Output nets */
wire t_9870,   t_9871,   t_9872;
/* u1_3421 Output nets */
wire t_9873,   t_9874;
/* u2_3422 Output nets */
wire t_9875,   t_9876,   t_9877;
/* u1_3423 Output nets */
wire t_9878,   t_9879;
/* u2_3424 Output nets */
wire t_9880,   t_9881,   t_9882;
/* u1_3425 Output nets */
wire t_9883,   t_9884;
/* u2_3426 Output nets */
wire t_9885,   t_9886,   t_9887;
/* u2_3427 Output nets */
wire t_9888,   t_9889,   t_9890;
/* u2_3428 Output nets */
wire t_9891,   t_9892,   t_9893;
/* u1_3429 Output nets */
wire t_9894,   t_9895;
/* u2_3430 Output nets */
wire t_9896,   t_9897,   t_9898;
/* u1_3431 Output nets */
wire t_9899,   t_9900;
/* u2_3432 Output nets */
wire t_9901,   t_9902,   t_9903;
/* u2_3433 Output nets */
wire t_9904,   t_9905,   t_9906;
/* u2_3434 Output nets */
wire t_9907,   t_9908,   t_9909;
/* u2_3435 Output nets */
wire t_9910,   t_9911,   t_9912;
/* u2_3436 Output nets */
wire t_9913,   t_9914,   t_9915;
/* u1_3437 Output nets */
wire t_9916,   t_9917;
/* u2_3438 Output nets */
wire t_9918,   t_9919,   t_9920;
/* u2_3439 Output nets */
wire t_9921,   t_9922,   t_9923;
/* u2_3440 Output nets */
wire t_9924,   t_9925,   t_9926;
/* u2_3441 Output nets */
wire t_9927,   t_9928,   t_9929;
/* u2_3442 Output nets */
wire t_9930,   t_9931,   t_9932;
/* u2_3443 Output nets */
wire t_9933,   t_9934,   t_9935;
/* u2_3444 Output nets */
wire t_9936,   t_9937,   t_9938;
/* u2_3445 Output nets */
wire t_9939,   t_9940,   t_9941;
/* u2_3446 Output nets */
wire t_9942,   t_9943,   t_9944;
/* u2_3447 Output nets */
wire t_9945,   t_9946,   t_9947;
/* u2_3448 Output nets */
wire t_9948,   t_9949,   t_9950;
/* u2_3449 Output nets */
wire t_9951,   t_9952,   t_9953;
/* u2_3450 Output nets */
wire t_9954,   t_9955,   t_9956;
/* u2_3451 Output nets */
wire t_9957,   t_9958,   t_9959;
/* u2_3452 Output nets */
wire t_9960,   t_9961,   t_9962;
/* u2_3453 Output nets */
wire t_9963,   t_9964,   t_9965;
/* u2_3454 Output nets */
wire t_9966,   t_9967,   t_9968;
/* u2_3455 Output nets */
wire t_9969,   t_9970,   t_9971;
/* u2_3456 Output nets */
wire t_9972,   t_9973,   t_9974;
/* u2_3457 Output nets */
wire t_9975,   t_9976,   t_9977;
/* u2_3458 Output nets */
wire t_9978,   t_9979,   t_9980;
/* u2_3459 Output nets */
wire t_9981,   t_9982,   t_9983;
/* u0_3460 Output nets */
wire t_9984,   t_9985;
/* u2_3461 Output nets */
wire t_9986,   t_9987,   t_9988;
/* u2_3462 Output nets */
wire t_9989,   t_9990,   t_9991;
/* u0_3463 Output nets */
wire t_9992,   t_9993;
/* u2_3464 Output nets */
wire t_9994,   t_9995,   t_9996;
/* u2_3465 Output nets */
wire t_9997,   t_9998,   t_9999;
/* u0_3466 Output nets */
wire t_10000,  t_10001;
/* u2_3467 Output nets */
wire t_10002,  t_10003,  t_10004;
/* u2_3468 Output nets */
wire t_10005,  t_10006,  t_10007;
/* u1_3469 Output nets */
wire t_10008,  t_10009;
/* u2_3470 Output nets */
wire t_10010,  t_10011,  t_10012;
/* u2_3471 Output nets */
wire t_10013,  t_10014,  t_10015;
/* u1_3472 Output nets */
wire t_10016,  t_10017;
/* u2_3473 Output nets */
wire t_10018,  t_10019,  t_10020;
/* u2_3474 Output nets */
wire t_10021,  t_10022,  t_10023;
/* u0_3475 Output nets */
wire t_10024,  t_10025;
/* u2_3476 Output nets */
wire t_10026,  t_10027,  t_10028;
/* u2_3477 Output nets */
wire t_10029,  t_10030,  t_10031;
/* u1_3478 Output nets */
wire t_10032,  t_10033;
/* u2_3479 Output nets */
wire t_10034,  t_10035,  t_10036;
/* u2_3480 Output nets */
wire t_10037,  t_10038,  t_10039;
/* u1_3481 Output nets */
wire t_10040,  t_10041;
/* u2_3482 Output nets */
wire t_10042,  t_10043,  t_10044;
/* u2_3483 Output nets */
wire t_10045,  t_10046,  t_10047;
/* u1_3484 Output nets */
wire t_10048,  t_10049;
/* u2_3485 Output nets */
wire t_10050,  t_10051,  t_10052;
/* u2_3486 Output nets */
wire t_10053,  t_10054,  t_10055;
/* u1_3487 Output nets */
wire t_10056,  t_10057;
/* u2_3488 Output nets */
wire t_10058,  t_10059,  t_10060;
/* u2_3489 Output nets */
wire t_10061,  t_10062,  t_10063;
/* u1_3490 Output nets */
wire t_10064,  t_10065;
/* u2_3491 Output nets */
wire t_10066,  t_10067,  t_10068;
/* u2_3492 Output nets */
wire t_10069,  t_10070,  t_10071;
/* u1_3493 Output nets */
wire t_10072,  t_10073;
/* u2_3494 Output nets */
wire t_10074,  t_10075,  t_10076;
/* u2_3495 Output nets */
wire t_10077,  t_10078,  t_10079;
/* u1_3496 Output nets */
wire t_10080,  t_10081;
/* u2_3497 Output nets */
wire t_10082,  t_10083,  t_10084;
/* u2_3498 Output nets */
wire t_10085,  t_10086,  t_10087;
/* u1_3499 Output nets */
wire t_10088,  t_10089;
/* u2_3500 Output nets */
wire t_10090,  t_10091,  t_10092;
/* u2_3501 Output nets */
wire t_10093,  t_10094,  t_10095;
/* u1_3502 Output nets */
wire t_10096,  t_10097;
/* u2_3503 Output nets */
wire t_10098,  t_10099,  t_10100;
/* u2_3504 Output nets */
wire t_10101,  t_10102,  t_10103;
/* u1_3505 Output nets */
wire t_10104,  t_10105;
/* u2_3506 Output nets */
wire t_10106,  t_10107,  t_10108;
/* u2_3507 Output nets */
wire t_10109,  t_10110,  t_10111;
/* u2_3508 Output nets */
wire t_10112,  t_10113,  t_10114;
/* u2_3509 Output nets */
wire t_10115,  t_10116,  t_10117;
/* u2_3510 Output nets */
wire t_10118,  t_10119,  t_10120;
/* u1_3511 Output nets */
wire t_10121,  t_10122;
/* u2_3512 Output nets */
wire t_10123,  t_10124,  t_10125;
/* u2_3513 Output nets */
wire t_10126,  t_10127,  t_10128;
/* u1_3514 Output nets */
wire t_10129,  t_10130;
/* u2_3515 Output nets */
wire t_10131,  t_10132,  t_10133;
/* u2_3516 Output nets */
wire t_10134,  t_10135,  t_10136;
/* u2_3517 Output nets */
wire t_10137,  t_10138,  t_10139;
/* u2_3518 Output nets */
wire t_10140,  t_10141,  t_10142;
/* u2_3519 Output nets */
wire t_10143,  t_10144,  t_10145;
/* u2_3520 Output nets */
wire t_10146,  t_10147,  t_10148;
/* u2_3521 Output nets */
wire t_10149,  t_10150,  t_10151;
/* u2_3522 Output nets */
wire t_10152,  t_10153,  t_10154;
/* u1_3523 Output nets */
wire t_10155,  t_10156;
/* u2_3524 Output nets */
wire t_10157,  t_10158,  t_10159;
/* u2_3525 Output nets */
wire t_10160,  t_10161,  t_10162;
/* u2_3526 Output nets */
wire t_10163,  t_10164,  t_10165;
/* u2_3527 Output nets */
wire t_10166,  t_10167,  t_10168;
/* u2_3528 Output nets */
wire t_10169,  t_10170,  t_10171;
/* u2_3529 Output nets */
wire t_10172,  t_10173,  t_10174;
/* u2_3530 Output nets */
wire t_10175,  t_10176,  t_10177;
/* u2_3531 Output nets */
wire t_10178,  t_10179,  t_10180;
/* u2_3532 Output nets */
wire t_10181,  t_10182,  t_10183;
/* u2_3533 Output nets */
wire t_10184,  t_10185,  t_10186;
/* u2_3534 Output nets */
wire t_10187,  t_10188,  t_10189;
/* u2_3535 Output nets */
wire t_10190,  t_10191,  t_10192;
/* u2_3536 Output nets */
wire t_10193,  t_10194,  t_10195;
/* u2_3537 Output nets */
wire t_10196,  t_10197,  t_10198;
/* u2_3538 Output nets */
wire t_10199,  t_10200,  t_10201;
/* u2_3539 Output nets */
wire t_10202,  t_10203,  t_10204;
/* u2_3540 Output nets */
wire t_10205,  t_10206,  t_10207;
/* u2_3541 Output nets */
wire t_10208,  t_10209,  t_10210;
/* u2_3542 Output nets */
wire t_10211,  t_10212,  t_10213;
/* u2_3543 Output nets */
wire t_10214,  t_10215,  t_10216;
/* u2_3544 Output nets */
wire t_10217,  t_10218,  t_10219;
/* u2_3545 Output nets */
wire t_10220,  t_10221,  t_10222;
/* u2_3546 Output nets */
wire t_10223,  t_10224,  t_10225;
/* u2_3547 Output nets */
wire t_10226,  t_10227,  t_10228;
/* u2_3548 Output nets */
wire t_10229,  t_10230,  t_10231;
/* u2_3549 Output nets */
wire t_10232,  t_10233,  t_10234;
/* u2_3550 Output nets */
wire t_10235,  t_10236,  t_10237;
/* u2_3551 Output nets */
wire t_10238,  t_10239,  t_10240;
/* u2_3552 Output nets */
wire t_10241,  t_10242,  t_10243;
/* u2_3553 Output nets */
wire t_10244,  t_10245,  t_10246;
/* u2_3554 Output nets */
wire t_10247,  t_10248,  t_10249;
/* u2_3555 Output nets */
wire t_10250,  t_10251,  t_10252;
/* u2_3556 Output nets */
wire t_10253,  t_10254,  t_10255;
/* u0_3557 Output nets */
wire t_10256,  t_10257;
/* u2_3558 Output nets */
wire t_10258,  t_10259,  t_10260;
/* u2_3559 Output nets */
wire t_10261,  t_10262,  t_10263;
/* u2_3560 Output nets */
wire t_10264,  t_10265,  t_10266;
/* u0_3561 Output nets */
wire t_10267,  t_10268;
/* u2_3562 Output nets */
wire t_10269,  t_10270,  t_10271;
/* u2_3563 Output nets */
wire t_10272,  t_10273,  t_10274;
/* u2_3564 Output nets */
wire t_10275,  t_10276,  t_10277;
/* u0_3565 Output nets */
wire t_10278,  t_10279;
/* u2_3566 Output nets */
wire t_10280,  t_10281,  t_10282;
/* u2_3567 Output nets */
wire t_10283,  t_10284,  t_10285;
/* u2_3568 Output nets */
wire t_10286,  t_10287,  t_10288;
/* u1_3569 Output nets */
wire t_10289,  t_10290;
/* u2_3570 Output nets */
wire t_10291,  t_10292,  t_10293;
/* u2_3571 Output nets */
wire t_10294,  t_10295,  t_10296;
/* u2_3572 Output nets */
wire t_10297,  t_10298,  t_10299;
/* u1_3573 Output nets */
wire t_10300,  t_10301;
/* u2_3574 Output nets */
wire t_10302,  t_10303,  t_10304;
/* u2_3575 Output nets */
wire t_10305,  t_10306,  t_10307;
/* u2_3576 Output nets */
wire t_10308,  t_10309,  t_10310;
/* u0_3577 Output nets */
wire t_10311,  t_10312;
/* u2_3578 Output nets */
wire t_10313,  t_10314,  t_10315;
/* u2_3579 Output nets */
wire t_10316,  t_10317,  t_10318;
/* u2_3580 Output nets */
wire t_10319,  t_10320,  t_10321;
/* u1_3581 Output nets */
wire t_10322,  t_10323;
/* u2_3582 Output nets */
wire t_10324,  t_10325,  t_10326;
/* u2_3583 Output nets */
wire t_10327,  t_10328,  t_10329;
/* u2_3584 Output nets */
wire t_10330,  t_10331,  t_10332;
/* u1_3585 Output nets */
wire t_10333,  t_10334;
/* u2_3586 Output nets */
wire t_10335,  t_10336,  t_10337;
/* u2_3587 Output nets */
wire t_10338,  t_10339,  t_10340;
/* u2_3588 Output nets */
wire t_10341,  t_10342,  t_10343;
/* u1_3589 Output nets */
wire t_10344,  t_10345;
/* u2_3590 Output nets */
wire t_10346,  t_10347,  t_10348;
/* u2_3591 Output nets */
wire t_10349,  t_10350,  t_10351;
/* u2_3592 Output nets */
wire t_10352,  t_10353,  t_10354;
/* u1_3593 Output nets */
wire t_10355,  t_10356;
/* u2_3594 Output nets */
wire t_10357,  t_10358,  t_10359;
/* u2_3595 Output nets */
wire t_10360,  t_10361,  t_10362;
/* u2_3596 Output nets */
wire t_10363,  t_10364,  t_10365;
/* u1_3597 Output nets */
wire t_10366,  t_10367;
/* u2_3598 Output nets */
wire t_10368,  t_10369,  t_10370;
/* u2_3599 Output nets */
wire t_10371,  t_10372,  t_10373;
/* u2_3600 Output nets */
wire t_10374,  t_10375,  t_10376;
/* u1_3601 Output nets */
wire t_10377,  t_10378;
/* u2_3602 Output nets */
wire t_10379,  t_10380,  t_10381;
/* u2_3603 Output nets */
wire t_10382,  t_10383,  t_10384;
/* u2_3604 Output nets */
wire t_10385,  t_10386,  t_10387;
/* u1_3605 Output nets */
wire t_10388,  t_10389;
/* u2_3606 Output nets */
wire t_10390,  t_10391,  t_10392;
/* u2_3607 Output nets */
wire t_10393,  t_10394,  t_10395;
/* u2_3608 Output nets */
wire t_10396,  t_10397,  t_10398;
/* u1_3609 Output nets */
wire t_10399,  t_10400;
/* u2_3610 Output nets */
wire t_10401,  t_10402,  t_10403;
/* u2_3611 Output nets */
wire t_10404,  t_10405,  t_10406;
/* u2_3612 Output nets */
wire t_10407,  t_10408,  t_10409;
/* u1_3613 Output nets */
wire t_10410,  t_10411;
/* u2_3614 Output nets */
wire t_10412,  t_10413,  t_10414;
/* u2_3615 Output nets */
wire t_10415,  t_10416,  t_10417;
/* u2_3616 Output nets */
wire t_10418,  t_10419,  t_10420;
/* u1_3617 Output nets */
wire t_10421,  t_10422;
/* u2_3618 Output nets */
wire t_10423,  t_10424,  t_10425;
/* u2_3619 Output nets */
wire t_10426,  t_10427,  t_10428;
/* u2_3620 Output nets */
wire t_10429,  t_10430,  t_10431;
/* u2_3621 Output nets */
wire t_10432,  t_10433,  t_10434;
/* u2_3622 Output nets */
wire t_10435,  t_10436,  t_10437;
/* u2_3623 Output nets */
wire t_10438,  t_10439,  t_10440;
/* u2_3624 Output nets */
wire t_10441,  t_10442,  t_10443;
/* u1_3625 Output nets */
wire t_10444,  t_10445;
/* u2_3626 Output nets */
wire t_10446,  t_10447,  t_10448;
/* u2_3627 Output nets */
wire t_10449,  t_10450,  t_10451;
/* u2_3628 Output nets */
wire t_10452,  t_10453,  t_10454;
/* u1_3629 Output nets */
wire t_10455,  t_10456;
/* u2_3630 Output nets */
wire t_10457,  t_10458,  t_10459;
/* u2_3631 Output nets */
wire t_10460,  t_10461,  t_10462;
/* u2_3632 Output nets */
wire t_10463,  t_10464,  t_10465;
/* u2_3633 Output nets */
wire t_10466,  t_10467,  t_10468;
/* u2_3634 Output nets */
wire t_10469,  t_10470,  t_10471;
/* u2_3635 Output nets */
wire t_10472,  t_10473,  t_10474;
/* u2_3636 Output nets */
wire t_10475,  t_10476,  t_10477;
/* u2_3637 Output nets */
wire t_10478,  t_10479,  t_10480;
/* u2_3638 Output nets */
wire t_10481,  t_10482,  t_10483;
/* u2_3639 Output nets */
wire t_10484,  t_10485,  t_10486;
/* u2_3640 Output nets */
wire t_10487,  t_10488,  t_10489;
/* u1_3641 Output nets */
wire t_10490,  t_10491;
/* u2_3642 Output nets */
wire t_10492,  t_10493,  t_10494;
/* u2_3643 Output nets */
wire t_10495,  t_10496,  t_10497;
/* u2_3644 Output nets */
wire t_10498,  t_10499,  t_10500;
/* u2_3645 Output nets */
wire t_10501,  t_10502,  t_10503;
/* u2_3646 Output nets */
wire t_10504,  t_10505,  t_10506;
/* u2_3647 Output nets */
wire t_10507,  t_10508,  t_10509;
/* u2_3648 Output nets */
wire t_10510,  t_10511,  t_10512;
/* u2_3649 Output nets */
wire t_10513,  t_10514,  t_10515;
/* u2_3650 Output nets */
wire t_10516,  t_10517,  t_10518;
/* u2_3651 Output nets */
wire t_10519,  t_10520,  t_10521;
/* u2_3652 Output nets */
wire t_10522,  t_10523,  t_10524;
/* u2_3653 Output nets */
wire t_10525,  t_10526,  t_10527;
/* u2_3654 Output nets */
wire t_10528,  t_10529,  t_10530;
/* u2_3655 Output nets */
wire t_10531,  t_10532,  t_10533;
/* u2_3656 Output nets */
wire t_10534,  t_10535,  t_10536;
/* u2_3657 Output nets */
wire t_10537,  t_10538,  t_10539;
/* u2_3658 Output nets */
wire t_10540,  t_10541,  t_10542;
/* u2_3659 Output nets */
wire t_10543,  t_10544,  t_10545;
/* u2_3660 Output nets */
wire t_10546,  t_10547,  t_10548;
/* u2_3661 Output nets */
wire t_10549,  t_10550,  t_10551;
/* u2_3662 Output nets */
wire t_10552,  t_10553,  t_10554;
/* u2_3663 Output nets */
wire t_10555,  t_10556,  t_10557;
/* u2_3664 Output nets */
wire t_10558,  t_10559,  t_10560;
/* u2_3665 Output nets */
wire t_10561,  t_10562,  t_10563;
/* u2_3666 Output nets */
wire t_10564,  t_10565,  t_10566;
/* u2_3667 Output nets */
wire t_10567,  t_10568,  t_10569;
/* u2_3668 Output nets */
wire t_10570,  t_10571,  t_10572;
/* u2_3669 Output nets */
wire t_10573,  t_10574,  t_10575;
/* u2_3670 Output nets */
wire t_10576,  t_10577,  t_10578;
/* u2_3671 Output nets */
wire t_10579,  t_10580,  t_10581;
/* u2_3672 Output nets */
wire t_10582,  t_10583,  t_10584;
/* u2_3673 Output nets */
wire t_10585,  t_10586,  t_10587;
/* u2_3674 Output nets */
wire t_10588,  t_10589,  t_10590;
/* u2_3675 Output nets */
wire t_10591,  t_10592,  t_10593;
/* u2_3676 Output nets */
wire t_10594,  t_10595,  t_10596;
/* u2_3677 Output nets */
wire t_10597,  t_10598,  t_10599;
/* u2_3678 Output nets */
wire t_10600,  t_10601,  t_10602;
/* u2_3679 Output nets */
wire t_10603,  t_10604,  t_10605;
/* u2_3680 Output nets */
wire t_10606,  t_10607,  t_10608;
/* u2_3681 Output nets */
wire t_10609,  t_10610,  t_10611;
/* u2_3682 Output nets */
wire t_10612,  t_10613,  t_10614;
/* u2_3683 Output nets */
wire t_10615,  t_10616,  t_10617;
/* u2_3684 Output nets */
wire t_10618,  t_10619,  t_10620;
/* u2_3685 Output nets */
wire t_10621,  t_10622,  t_10623;
/* u2_3686 Output nets */
wire t_10624,  t_10625,  t_10626;
/* u2_3687 Output nets */
wire t_10627,  t_10628,  t_10629;
/* u2_3688 Output nets */
wire t_10630,  t_10631,  t_10632;
/* u2_3689 Output nets */
wire t_10633,  t_10634,  t_10635;
/* u2_3690 Output nets */
wire t_10636,  t_10637,  t_10638;
/* u2_3691 Output nets */
wire t_10639,  t_10640,  t_10641;
/* u2_3692 Output nets */
wire t_10642,  t_10643,  t_10644;
/* u2_3693 Output nets */
wire t_10645,  t_10646,  t_10647;
/* u2_3694 Output nets */
wire t_10648,  t_10649,  t_10650;
/* u2_3695 Output nets */
wire t_10651,  t_10652,  t_10653;
/* u2_3696 Output nets */
wire t_10654,  t_10655,  t_10656;
/* u2_3697 Output nets */
wire t_10657,  t_10658,  t_10659;
/* u2_3698 Output nets */
wire t_10660,  t_10661,  t_10662;
/* u2_3699 Output nets */
wire t_10663,  t_10664,  t_10665;
/* u2_3700 Output nets */
wire t_10666,  t_10667,  t_10668;
/* u2_3701 Output nets */
wire t_10669,  t_10670,  t_10671;
/* u2_3702 Output nets */
wire t_10672,  t_10673,  t_10674;
/* u2_3703 Output nets */
wire t_10675,  t_10676,  t_10677;
/* u2_3704 Output nets */
wire t_10678,  t_10679,  t_10680;
/* u2_3705 Output nets */
wire t_10681,  t_10682,  t_10683;
/* u2_3706 Output nets */
wire t_10684,  t_10685,  t_10686;
/* u2_3707 Output nets */
wire t_10687,  t_10688,  t_10689;
/* u2_3708 Output nets */
wire t_10690,  t_10691,  t_10692;
/* u1_3709 Output nets */
wire t_10693,  t_10694;
/* u2_3710 Output nets */
wire t_10695,  t_10696,  t_10697;
/* u2_3711 Output nets */
wire t_10698,  t_10699,  t_10700;
/* u2_3712 Output nets */
wire t_10701,  t_10702,  t_10703;
/* u2_3713 Output nets */
wire t_10704,  t_10705,  t_10706;
/* u2_3714 Output nets */
wire t_10707,  t_10708,  t_10709;
/* u2_3715 Output nets */
wire t_10710,  t_10711,  t_10712;
/* u2_3716 Output nets */
wire t_10713,  t_10714,  t_10715;
/* u1_3717 Output nets */
wire t_10716,  t_10717;
/* u2_3718 Output nets */
wire t_10718,  t_10719,  t_10720;
/* u2_3719 Output nets */
wire t_10721,  t_10722,  t_10723;
/* u2_3720 Output nets */
wire t_10724,  t_10725,  t_10726;
/* u1_3721 Output nets */
wire t_10727,  t_10728;
/* u2_3722 Output nets */
wire t_10729,  t_10730,  t_10731;
/* u2_3723 Output nets */
wire t_10732,  t_10733,  t_10734;
/* u2_3724 Output nets */
wire t_10735,  t_10736,  t_10737;
/* u1_3725 Output nets */
wire t_10738,  t_10739;
/* u2_3726 Output nets */
wire t_10740,  t_10741,  t_10742;
/* u2_3727 Output nets */
wire t_10743,  t_10744,  t_10745;
/* u2_3728 Output nets */
wire t_10746,  t_10747,  t_10748;
/* u1_3729 Output nets */
wire t_10749,  t_10750;
/* u2_3730 Output nets */
wire t_10751,  t_10752,  t_10753;
/* u2_3731 Output nets */
wire t_10754,  t_10755,  t_10756;
/* u2_3732 Output nets */
wire t_10757,  t_10758,  t_10759;
/* u1_3733 Output nets */
wire t_10760,  t_10761;
/* u2_3734 Output nets */
wire t_10762,  t_10763,  t_10764;
/* u2_3735 Output nets */
wire t_10765,  t_10766,  t_10767;
/* u2_3736 Output nets */
wire t_10768,  t_10769,  t_10770;
/* u1_3737 Output nets */
wire t_10771,  t_10772;
/* u2_3738 Output nets */
wire t_10773,  t_10774,  t_10775;
/* u2_3739 Output nets */
wire t_10776,  t_10777,  t_10778;
/* u2_3740 Output nets */
wire t_10779,  t_10780,  t_10781;
/* u1_3741 Output nets */
wire t_10782,  t_10783;
/* u2_3742 Output nets */
wire t_10784,  t_10785,  t_10786;
/* u2_3743 Output nets */
wire t_10787,  t_10788,  t_10789;
/* u2_3744 Output nets */
wire t_10790,  t_10791,  t_10792;
/* u1_3745 Output nets */
wire t_10793,  t_10794;
/* u2_3746 Output nets */
wire t_10795,  t_10796,  t_10797;
/* u2_3747 Output nets */
wire t_10798,  t_10799,  t_10800;
/* u2_3748 Output nets */
wire t_10801,  t_10802,  t_10803;
/* u1_3749 Output nets */
wire t_10804,  t_10805;
/* u2_3750 Output nets */
wire t_10806,  t_10807,  t_10808;
/* u2_3751 Output nets */
wire t_10809,  t_10810,  t_10811;
/* u2_3752 Output nets */
wire t_10812,  t_10813,  t_10814;
/* u1_3753 Output nets */
wire t_10815,  t_10816;
/* u2_3754 Output nets */
wire t_10817,  t_10818,  t_10819;
/* u2_3755 Output nets */
wire t_10820,  t_10821,  t_10822;
/* u2_3756 Output nets */
wire t_10823,  t_10824,  t_10825;
/* u1_3757 Output nets */
wire t_10826,  t_10827;
/* u2_3758 Output nets */
wire t_10828,  t_10829,  t_10830;
/* u2_3759 Output nets */
wire t_10831,  t_10832,  t_10833;
/* u2_3760 Output nets */
wire t_10834,  t_10835,  t_10836;
/* u1_3761 Output nets */
wire t_10837,  t_10838;
/* u2_3762 Output nets */
wire t_10839,  t_10840,  t_10841;
/* u2_3763 Output nets */
wire t_10842,  t_10843,  t_10844;
/* u2_3764 Output nets */
wire t_10845,  t_10846,  t_10847;
/* u1_3765 Output nets */
wire t_10848,  t_10849;
/* u2_3766 Output nets */
wire t_10850,  t_10851,  t_10852;
/* u2_3767 Output nets */
wire t_10853,  t_10854,  t_10855;
/* u2_3768 Output nets */
wire t_10856,  t_10857,  t_10858;
/* u1_3769 Output nets */
wire t_10859,  t_10860;
/* u2_3770 Output nets */
wire t_10861,  t_10862,  t_10863;
/* u2_3771 Output nets */
wire t_10864,  t_10865,  t_10866;
/* u2_3772 Output nets */
wire t_10867,  t_10868,  t_10869;
/* u0_3773 Output nets */
wire t_10870,  t_10871;
/* u2_3774 Output nets */
wire t_10872,  t_10873,  t_10874;
/* u2_3775 Output nets */
wire t_10875,  t_10876,  t_10877;
/* u2_3776 Output nets */
wire t_10878,  t_10879,  t_10880;
/* u1_3777 Output nets */
wire t_10881,  t_10882;
/* u2_3778 Output nets */
wire t_10883,  t_10884,  t_10885;
/* u2_3779 Output nets */
wire t_10886,  t_10887,  t_10888;
/* u2_3780 Output nets */
wire t_10889,  t_10890,  t_10891;
/* u0_3781 Output nets */
wire t_10892,  t_10893;
/* u2_3782 Output nets */
wire t_10894,  t_10895,  t_10896;
/* u2_3783 Output nets */
wire t_10897,  t_10898,  t_10899;
/* u2_3784 Output nets */
wire t_10900,  t_10901,  t_10902;
/* u0_3785 Output nets */
wire t_10903,  t_10904;
/* u2_3786 Output nets */
wire t_10905,  t_10906,  t_10907;
/* u2_3787 Output nets */
wire t_10908,  t_10909,  t_10910;
/* u2_3788 Output nets */
wire t_10911,  t_10912,  t_10913;
/* u0_3789 Output nets */
wire t_10914,  t_10915;
/* u2_3790 Output nets */
wire t_10916,  t_10917,  t_10918;
/* u2_3791 Output nets */
wire t_10919,  t_10920,  t_10921;
/* u2_3792 Output nets */
wire t_10922,  t_10923,  t_10924;
/* u0_3793 Output nets */
wire t_10925,  t_10926;
/* u2_3794 Output nets */
wire t_10927,  t_10928,  t_10929;
/* u2_3795 Output nets */
wire t_10930,  t_10931,  t_10932;
/* u2_3796 Output nets */
wire t_10933,  t_10934,  t_10935;
/* u0_3797 Output nets */
wire t_10936,  t_10937;
/* u2_3798 Output nets */
wire t_10938,  t_10939,  t_10940;
/* u2_3799 Output nets */
wire t_10941,  t_10942,  t_10943;
/* u2_3800 Output nets */
wire t_10944,  t_10945,  t_10946;
/* u0_3801 Output nets */
wire t_10947,  t_10948;
/* u2_3802 Output nets */
wire t_10949,  t_10950,  t_10951;
/* u2_3803 Output nets */
wire t_10952,  t_10953,  t_10954;
/* u2_3804 Output nets */
wire t_10955,  t_10956,  t_10957;
/* u0_3805 Output nets */
wire t_10958,  t_10959;
/* u2_3806 Output nets */
wire t_10960,  t_10961,  t_10962;
/* u2_3807 Output nets */
wire t_10963,  t_10964,  t_10965;
/* u2_3808 Output nets */
wire t_10966,  t_10967,  t_10968;
/* u0_3809 Output nets */
wire t_10969,  t_10970;
/* u2_3810 Output nets */
wire t_10971,  t_10972,  t_10973;
/* u2_3811 Output nets */
wire t_10974,  t_10975,  t_10976;
/* u2_3812 Output nets */
wire t_10977,  t_10978,  t_10979;
/* u2_3813 Output nets */
wire t_10980,  t_10981,  t_10982;
/* u2_3814 Output nets */
wire t_10983,  t_10984,  t_10985;
/* u2_3815 Output nets */
wire t_10986,  t_10987,  t_10988;
/* u2_3816 Output nets */
wire t_10989,  t_10990,  t_10991;
/* u2_3817 Output nets */
wire t_10992,  t_10993,  t_10994;
/* u2_3818 Output nets */
wire t_10995,  t_10996,  t_10997;
/* u2_3819 Output nets */
wire t_10998,  t_10999,  t_11000;
/* u2_3820 Output nets */
wire t_11001,  t_11002,  t_11003;
/* u2_3821 Output nets */
wire t_11004,  t_11005,  t_11006;
/* u2_3822 Output nets */
wire t_11007,  t_11008,  t_11009;
/* u2_3823 Output nets */
wire t_11010,  t_11011,  t_11012;
/* u2_3824 Output nets */
wire t_11013,  t_11014,  t_11015;
/* u2_3825 Output nets */
wire t_11016,  t_11017,  t_11018;
/* u2_3826 Output nets */
wire t_11019,  t_11020,  t_11021;
/* u2_3827 Output nets */
wire t_11022,  t_11023,  t_11024;
/* u2_3828 Output nets */
wire t_11025,  t_11026,  t_11027;
/* u2_3829 Output nets */
wire t_11028,  t_11029,  t_11030;
/* u1_3830 Output nets */
wire t_11031,  t_11032;
/* u2_3831 Output nets */
wire t_11033,  t_11034,  t_11035;
/* u2_3832 Output nets */
wire t_11036,  t_11037,  t_11038;
/* u2_3833 Output nets */
wire t_11039,  t_11040,  t_11041;
/* u2_3834 Output nets */
wire t_11042,  t_11043,  t_11044;
/* u2_3835 Output nets */
wire t_11045,  t_11046,  t_11047;
/* u1_3836 Output nets */
wire t_11048,  t_11049;
/* u2_3837 Output nets */
wire t_11050,  t_11051,  t_11052;
/* u2_3838 Output nets */
wire t_11053,  t_11054,  t_11055;
/* u1_3839 Output nets */
wire t_11056,  t_11057;
/* u2_3840 Output nets */
wire t_11058,  t_11059,  t_11060;
/* u2_3841 Output nets */
wire t_11061,  t_11062,  t_11063;
/* u1_3842 Output nets */
wire t_11064,  t_11065;
/* u2_3843 Output nets */
wire t_11066,  t_11067,  t_11068;
/* u2_3844 Output nets */
wire t_11069,  t_11070,  t_11071;
/* u1_3845 Output nets */
wire t_11072,  t_11073;
/* u2_3846 Output nets */
wire t_11074,  t_11075,  t_11076;
/* u2_3847 Output nets */
wire t_11077,  t_11078,  t_11079;
/* u1_3848 Output nets */
wire t_11080,  t_11081;
/* u2_3849 Output nets */
wire t_11082,  t_11083,  t_11084;
/* u2_3850 Output nets */
wire t_11085,  t_11086,  t_11087;
/* u1_3851 Output nets */
wire t_11088,  t_11089;
/* u2_3852 Output nets */
wire t_11090,  t_11091,  t_11092;
/* u2_3853 Output nets */
wire t_11093,  t_11094,  t_11095;
/* u1_3854 Output nets */
wire t_11096,  t_11097;
/* u2_3855 Output nets */
wire t_11098,  t_11099,  t_11100;
/* u2_3856 Output nets */
wire t_11101,  t_11102,  t_11103;
/* u1_3857 Output nets */
wire t_11104,  t_11105;
/* u2_3858 Output nets */
wire t_11106,  t_11107,  t_11108;
/* u2_3859 Output nets */
wire t_11109,  t_11110,  t_11111;
/* u1_3860 Output nets */
wire t_11112,  t_11113;
/* u2_3861 Output nets */
wire t_11114,  t_11115,  t_11116;
/* u2_3862 Output nets */
wire t_11117,  t_11118,  t_11119;
/* u1_3863 Output nets */
wire t_11120,  t_11121;
/* u2_3864 Output nets */
wire t_11122,  t_11123,  t_11124;
/* u2_3865 Output nets */
wire t_11125,  t_11126,  t_11127;
/* u1_3866 Output nets */
wire t_11128,  t_11129;
/* u2_3867 Output nets */
wire t_11130,  t_11131,  t_11132;
/* u2_3868 Output nets */
wire t_11133,  t_11134,  t_11135;
/* u1_3869 Output nets */
wire t_11136,  t_11137;
/* u2_3870 Output nets */
wire t_11138,  t_11139,  t_11140;
/* u2_3871 Output nets */
wire t_11141,  t_11142,  t_11143;
/* u1_3872 Output nets */
wire t_11144,  t_11145;
/* u2_3873 Output nets */
wire t_11146,  t_11147,  t_11148;
/* u2_3874 Output nets */
wire t_11149,  t_11150,  t_11151;
/* u1_3875 Output nets */
wire t_11152,  t_11153;
/* u2_3876 Output nets */
wire t_11154,  t_11155,  t_11156;
/* u2_3877 Output nets */
wire t_11157,  t_11158,  t_11159;
/* u0_3878 Output nets */
wire t_11160,  t_11161;
/* u2_3879 Output nets */
wire t_11162,  t_11163,  t_11164;
/* u2_3880 Output nets */
wire t_11165,  t_11166,  t_11167;
/* u1_3881 Output nets */
wire t_11168,  t_11169;
/* u2_3882 Output nets */
wire t_11170,  t_11171,  t_11172;
/* u2_3883 Output nets */
wire t_11173,  t_11174,  t_11175;
/* u0_3884 Output nets */
wire t_11176,  t_11177;
/* u2_3885 Output nets */
wire t_11178,  t_11179,  t_11180;
/* u2_3886 Output nets */
wire t_11181,  t_11182,  t_11183;
/* u0_3887 Output nets */
wire t_11184,  t_11185;
/* u2_3888 Output nets */
wire t_11186,  t_11187,  t_11188;
/* u2_3889 Output nets */
wire t_11189,  t_11190,  t_11191;
/* u0_3890 Output nets */
wire t_11192,  t_11193;
/* u2_3891 Output nets */
wire t_11194,  t_11195,  t_11196;
/* u2_3892 Output nets */
wire t_11197,  t_11198,  t_11199;
/* u0_3893 Output nets */
wire t_11200,  t_11201;
/* u2_3894 Output nets */
wire t_11202,  t_11203,  t_11204;
/* u2_3895 Output nets */
wire t_11205,  t_11206,  t_11207;
/* u0_3896 Output nets */
wire t_11208,  t_11209;
/* u2_3897 Output nets */
wire t_11210,  t_11211,  t_11212;
/* u2_3898 Output nets */
wire t_11213,  t_11214,  t_11215;
/* u0_3899 Output nets */
wire t_11216,  t_11217;
/* u2_3900 Output nets */
wire t_11218,  t_11219,  t_11220;
/* u2_3901 Output nets */
wire t_11221,  t_11222,  t_11223;
/* u0_3902 Output nets */
wire t_11224,  t_11225;
/* u2_3903 Output nets */
wire t_11226,  t_11227,  t_11228;
/* u2_3904 Output nets */
wire t_11229,  t_11230,  t_11231;
/* u0_3905 Output nets */
wire t_11232,  t_11233;
/* u2_3906 Output nets */
wire t_11234,  t_11235,  t_11236;
/* u2_3907 Output nets */
wire t_11237,  t_11238,  t_11239;
/* u2_3908 Output nets */
wire t_11240,  t_11241,  t_11242;
/* u2_3909 Output nets */
wire t_11243,  t_11244,  t_11245;
/* u2_3910 Output nets */
wire t_11246,  t_11247,  t_11248;
/* u2_3911 Output nets */
wire t_11249,  t_11250,  t_11251;
/* u2_3912 Output nets */
wire t_11252,  t_11253,  t_11254;
/* u2_3913 Output nets */
wire t_11255,  t_11256,  t_11257;
/* u2_3914 Output nets */
wire t_11258,  t_11259,  t_11260;
/* u2_3915 Output nets */
wire t_11261,  t_11262,  t_11263;
/* u2_3916 Output nets */
wire t_11264,  t_11265,  t_11266;
/* u2_3917 Output nets */
wire t_11267,  t_11268,  t_11269;
/* u2_3918 Output nets */
wire t_11270,  t_11271,  t_11272;
/* u1_3919 Output nets */
wire t_11273,  t_11274;
/* u2_3920 Output nets */
wire t_11275,  t_11276,  t_11277;
/* u2_3921 Output nets */
wire t_11278,  t_11279,  t_11280;
/* u2_3922 Output nets */
wire t_11281,  t_11282,  t_11283;
/* u1_3923 Output nets */
wire t_11284,  t_11285;
/* u2_3924 Output nets */
wire t_11286,  t_11287,  t_11288;
/* u1_3925 Output nets */
wire t_11289,  t_11290;
/* u2_3926 Output nets */
wire t_11291,  t_11292,  t_11293;
/* u1_3927 Output nets */
wire t_11294,  t_11295;
/* u2_3928 Output nets */
wire t_11296,  t_11297,  t_11298;
/* u1_3929 Output nets */
wire t_11299,  t_11300;
/* u2_3930 Output nets */
wire t_11301,  t_11302,  t_11303;
/* u1_3931 Output nets */
wire t_11304,  t_11305;
/* u2_3932 Output nets */
wire t_11306,  t_11307,  t_11308;
/* u1_3933 Output nets */
wire t_11309,  t_11310;
/* u2_3934 Output nets */
wire t_11311,  t_11312,  t_11313;
/* u1_3935 Output nets */
wire t_11314,  t_11315;
/* u2_3936 Output nets */
wire t_11316,  t_11317,  t_11318;
/* u1_3937 Output nets */
wire t_11319,  t_11320;
/* u2_3938 Output nets */
wire t_11321,  t_11322,  t_11323;
/* u1_3939 Output nets */
wire t_11324,  t_11325;
/* u2_3940 Output nets */
wire t_11326,  t_11327,  t_11328;
/* u1_3941 Output nets */
wire t_11329,  t_11330;
/* u2_3942 Output nets */
wire t_11331,  t_11332,  t_11333;
/* u1_3943 Output nets */
wire t_11334,  t_11335;
/* u2_3944 Output nets */
wire t_11336,  t_11337,  t_11338;
/* u1_3945 Output nets */
wire t_11339,  t_11340;
/* u2_3946 Output nets */
wire t_11341,  t_11342,  t_11343;
/* u1_3947 Output nets */
wire t_11344,  t_11345;
/* u2_3948 Output nets */
wire t_11346,  t_11347,  t_11348;
/* u1_3949 Output nets */
wire t_11349,  t_11350;
/* u2_3950 Output nets */
wire t_11351,  t_11352,  t_11353;
/* u0_3951 Output nets */
wire t_11354,  t_11355;
/* u2_3952 Output nets */
wire t_11356,  t_11357,  t_11358;
/* u1_3953 Output nets */
wire t_11359,  t_11360;
/* u2_3954 Output nets */
wire t_11361,  t_11362,  t_11363;
/* u0_3955 Output nets */
wire t_11364,  t_11365;
/* u2_3956 Output nets */
wire t_11366,  t_11367,  t_11368;
/* u0_3957 Output nets */
wire t_11369,  t_11370;
/* u2_3958 Output nets */
wire t_11371,  t_11372,  t_11373;
/* u0_3959 Output nets */
wire t_11374,  t_11375;
/* u2_3960 Output nets */
wire t_11376,  t_11377,  t_11378;
/* u0_3961 Output nets */
wire t_11379,  t_11380;
/* u2_3962 Output nets */
wire t_11381,  t_11382,  t_11383;
/* u0_3963 Output nets */
wire t_11384,  t_11385;
/* u2_3964 Output nets */
wire t_11386,  t_11387,  t_11388;
/* u0_3965 Output nets */
wire t_11389,  t_11390;
/* u2_3966 Output nets */
wire t_11391,  t_11392,  t_11393;
/* u0_3967 Output nets */
wire t_11394,  t_11395;
/* u2_3968 Output nets */
wire t_11396,  t_11397,  t_11398;
/* u0_3969 Output nets */
wire t_11399,  t_11400;
/* u2_3970 Output nets */
wire t_11401,  t_11402,  t_11403;
/* u2_3971 Output nets */
wire t_11404,  t_11405,  t_11406;
/* u2_3972 Output nets */
wire t_11407,  t_11408,  t_11409;
/* u2_3973 Output nets */
wire t_11410,  t_11411,  t_11412;
/* u2_3974 Output nets */
wire t_11413,  t_11414,  t_11415;
/* u2_3975 Output nets */
wire t_11416,  t_11417,  t_11418;
/* u1_3976 Output nets */
wire t_11419,  t_11420;
/* u1_3977 Output nets */
wire t_11421,  t_11422;
/* u1_3978 Output nets */
wire t_11423,  t_11424;
/* u1_3979 Output nets */
wire t_11425,  t_11426;
/* u1_3980 Output nets */
wire t_11427,  t_11428;
/* u1_3981 Output nets */
wire t_11429,  t_11430;
/* u1_3982 Output nets */
wire t_11431,  t_11432;
/* u1_3983 Output nets */
wire t_11433,  t_11434;
/* u1_3984 Output nets */
wire t_11435,  t_11436;
/* u1_3985 Output nets */
wire t_11437,  t_11438;
/* u0_3986 Output nets */
wire t_11439,  t_11440;
/* u1_3987 Output nets */
wire t_11441,  t_11442;
/* u0_3988 Output nets */
wire t_11443,  t_11444;
/* u0_3989 Output nets */
wire t_11445,  t_11446;
/* u0_3990 Output nets */
wire t_11447,  t_11448;
/* u0_3991 Output nets */
wire t_11449,  t_11450;
/* u0_3992 Output nets */
wire t_11451,  t_11452;
/* u0_3993 Output nets */
wire t_11453,  t_11454;
/* u0_3994 Output nets */
wire t_11455,  t_11456;
/* u0_3995 Output nets */
wire t_11457,  t_11458;
/* u0_3996 Output nets */
wire t_11459;

/* compress stage 3 */
half_adder u0_3362(.a(t_6442), .b(t_2), .o(t_9728), .cout(t_9729));
half_adder u0_3363(.a(t_6444), .b(t_6), .o(t_9730), .cout(t_9731));
half_adder u0_3364(.a(t_6446), .b(t_6447), .o(t_9732), .cout(t_9733));
half_adder u0_3365(.a(t_6448), .b(t_6449), .o(t_9734), .cout(t_9735));
half_adder u0_3366(.a(t_6450), .b(t_6451), .o(t_9736), .cout(t_9737));
half_adder u0_3367(.a(t_6452), .b(t_6453), .o(t_9738), .cout(t_9739));
compressor_3_2 u1_3368(.a(t_6456), .b(t_6458), .cin(t_28), .o(t_9740), .cout(t_9741));
half_adder u0_3369(.a(t_6459), .b(t_6460), .o(t_9742), .cout(t_9743));
half_adder u0_3370(.a(t_6462), .b(t_41), .o(t_9744), .cout(t_9745));
half_adder u0_3371(.a(t_6463), .b(t_6465), .o(t_9746), .cout(t_9747));
half_adder u0_3372(.a(t_6466), .b(t_6468), .o(t_9748), .cout(t_9749));
compressor_3_2 u1_3373(.a(t_6469), .b(t_6471), .cin(t_58), .o(t_9750), .cout(t_9751));
compressor_3_2 u1_3374(.a(t_6472), .b(t_6474), .cin(t_64), .o(t_9752), .cout(t_9753));
compressor_3_2 u1_3375(.a(t_6475), .b(t_6480), .cin(t_6477), .o(t_9754), .cout(t_9755));
compressor_3_2 u1_3376(.a(t_6478), .b(t_6485), .cin(t_6482), .o(t_9756), .cout(t_9757));
compressor_3_2 u1_3377(.a(t_6483), .b(t_6490), .cin(t_6487), .o(t_9758), .cout(t_9759));
compressor_4_2 u2_3378(.a(t_6488), .b(t_6495), .c(t_6492), .d(t_99), .cin(t_9759), .o(t_9760), .co(t_9761), .cout(t_9762));
compressor_3_2 u1_3379(.a(t_6500), .b(t_6497), .cin(t_9762), .o(t_9763), .cout(t_9764));
compressor_3_2 u1_3380(.a(t_6498), .b(t_6505), .cin(t_6502), .o(t_9765), .cout(t_9766));
compressor_4_2 u2_3381(.a(t_6503), .b(t_6510), .c(t_6507), .d(t_125), .cin(t_9766), .o(t_9767), .co(t_9768), .cout(t_9769));
compressor_4_2 u2_3382(.a(t_6508), .b(t_6515), .c(t_6512), .d(t_134), .cin(t_9769), .o(t_9770), .co(t_9771), .cout(t_9772));
compressor_3_2 u1_3383(.a(t_6520), .b(t_6517), .cin(t_9772), .o(t_9773), .cout(t_9774));
compressor_4_2 u2_3384(.a(t_6521), .b(t_6518), .c(t_6526), .d(t_6523), .cin(t_156), .o(t_9775), .co(t_9776), .cout(t_9777));
compressor_4_2 u2_3385(.a(t_6524), .b(t_6531), .c(t_6528), .d(t_167), .cin(t_9777), .o(t_9778), .co(t_9779), .cout(t_9780));
compressor_4_2 u2_3386(.a(t_6529), .b(t_6536), .c(t_6533), .d(t_181), .cin(t_9780), .o(t_9781), .co(t_9782), .cout(t_9783));
compressor_4_2 u2_3387(.a(t_6537), .b(t_6534), .c(t_6542), .d(t_6539), .cin(t_9783), .o(t_9784), .co(t_9785), .cout(t_9786));
compressor_4_2 u2_3388(.a(t_6543), .b(t_6540), .c(t_6548), .d(t_6545), .cin(t_9786), .o(t_9787), .co(t_9788), .cout(t_9789));
compressor_4_2 u2_3389(.a(t_6546), .b(t_6554), .c(t_6551), .d(t_216), .cin(t_9789), .o(t_9790), .co(t_9791), .cout(t_9792));
compressor_4_2 u2_3390(.a(t_6552), .b(t_6560), .c(t_6557), .d(t_228), .cin(t_9792), .o(t_9793), .co(t_9794), .cout(t_9795));
compressor_4_2 u2_3391(.a(t_6558), .b(t_6569), .c(t_6566), .d(t_6563), .cin(t_9795), .o(t_9796), .co(t_9797), .cout(t_9798));
compressor_4_2 u2_3392(.a(t_6564), .b(t_6577), .c(t_6574), .d(t_6571), .cin(t_9798), .o(t_9799), .co(t_9800), .cout(t_9801));
compressor_4_2 u2_3393(.a(t_6572), .b(t_6585), .c(t_6582), .d(t_6579), .cin(t_9801), .o(t_9802), .co(t_9803), .cout(t_9804));
compressor_4_2 u2_3394(.a(t_6593), .b(t_6590), .c(t_6587), .d(t_287), .cin(t_9804), .o(t_9805), .co(t_9806), .cout(t_9807));
half_adder u0_3395(.a(t_6583), .b(t_6580), .o(t_9808), .cout(t_9809));
compressor_4_2 u2_3396(.a(t_6601), .b(t_6598), .c(t_6595), .d(t_9807), .cin(t_9809), .o(t_9810), .co(t_9811), .cout(t_9812));
half_adder u0_3397(.a(t_6591), .b(t_6588), .o(t_9813), .cout(t_9814));
compressor_4_2 u2_3398(.a(t_6609), .b(t_6606), .c(t_6603), .d(t_9812), .cin(t_9814), .o(t_9815), .co(t_9816), .cout(t_9817));
half_adder u0_3399(.a(t_6599), .b(t_6596), .o(t_9818), .cout(t_9819));
compressor_4_2 u2_3400(.a(t_6614), .b(t_6611), .c(t_331), .d(t_9817), .cin(t_9819), .o(t_9820), .co(t_9821), .cout(t_9822));
compressor_3_2 u1_3401(.a(t_6607), .b(t_6604), .cin(t_6617), .o(t_9823), .cout(t_9824));
compressor_4_2 u2_3402(.a(t_6622), .b(t_6619), .c(t_346), .d(t_9822), .cin(t_9824), .o(t_9825), .co(t_9826), .cout(t_9827));
compressor_3_2 u1_3403(.a(t_6615), .b(t_6612), .cin(t_6625), .o(t_9828), .cout(t_9829));
compressor_4_2 u2_3404(.a(t_6633), .b(t_6630), .c(t_6627), .d(t_9827), .cin(t_9829), .o(t_9830), .co(t_9831), .cout(t_9832));
half_adder u0_3405(.a(t_6623), .b(t_6620), .o(t_9833), .cout(t_9834));
compressor_4_2 u2_3406(.a(t_6639), .b(t_6636), .c(t_380), .d(t_9832), .cin(t_9834), .o(t_9835), .co(t_9836), .cout(t_9837));
compressor_3_2 u1_3407(.a(t_6631), .b(t_6628), .cin(t_6642), .o(t_9838), .cout(t_9839));
compressor_4_2 u2_3408(.a(t_6647), .b(t_6644), .c(t_397), .d(t_9837), .cin(t_9839), .o(t_9840), .co(t_9841), .cout(t_9842));
compressor_3_2 u1_3409(.a(t_6640), .b(t_6637), .cin(t_6650), .o(t_9843), .cout(t_9844));
compressor_4_2 u2_3410(.a(t_6655), .b(t_6652), .c(t_417), .d(t_9842), .cin(t_9844), .o(t_9845), .co(t_9846), .cout(t_9847));
compressor_3_2 u1_3411(.a(t_6648), .b(t_6645), .cin(t_6658), .o(t_9848), .cout(t_9849));
compressor_4_2 u2_3412(.a(t_6667), .b(t_6664), .c(t_6661), .d(t_9847), .cin(t_9849), .o(t_9850), .co(t_9851), .cout(t_9852));
compressor_3_2 u1_3413(.a(t_6659), .b(t_6656), .cin(t_6653), .o(t_9853), .cout(t_9854));
compressor_4_2 u2_3414(.a(t_6676), .b(t_6673), .c(t_6670), .d(t_9852), .cin(t_9854), .o(t_9855), .co(t_9856), .cout(t_9857));
compressor_3_2 u1_3415(.a(t_6668), .b(t_6665), .cin(t_6662), .o(t_9858), .cout(t_9859));
compressor_4_2 u2_3416(.a(t_6682), .b(t_6679), .c(t_470), .d(t_9857), .cin(t_9859), .o(t_9860), .co(t_9861), .cout(t_9862));
compressor_3_2 u1_3417(.a(t_6674), .b(t_6671), .cin(t_6685), .o(t_9863), .cout(t_9864));
compressor_4_2 u2_3418(.a(t_6691), .b(t_6688), .c(t_488), .d(t_9862), .cin(t_9864), .o(t_9865), .co(t_9866), .cout(t_9867));
compressor_3_2 u1_3419(.a(t_6683), .b(t_6680), .cin(t_6694), .o(t_9868), .cout(t_9869));
compressor_4_2 u2_3420(.a(t_6703), .b(t_6700), .c(t_6697), .d(t_9867), .cin(t_9869), .o(t_9870), .co(t_9871), .cout(t_9872));
compressor_3_2 u1_3421(.a(t_6692), .b(t_6689), .cin(t_6706), .o(t_9873), .cout(t_9874));
compressor_4_2 u2_3422(.a(t_6714), .b(t_6711), .c(t_6708), .d(t_9872), .cin(t_9874), .o(t_9875), .co(t_9876), .cout(t_9877));
compressor_3_2 u1_3423(.a(t_6701), .b(t_6698), .cin(t_6717), .o(t_9878), .cout(t_9879));
compressor_4_2 u2_3424(.a(t_6725), .b(t_6722), .c(t_6719), .d(t_9877), .cin(t_9879), .o(t_9880), .co(t_9881), .cout(t_9882));
compressor_3_2 u1_3425(.a(t_6712), .b(t_6709), .cin(t_6728), .o(t_9883), .cout(t_9884));
compressor_4_2 u2_3426(.a(t_6733), .b(t_6730), .c(t_571), .d(t_9882), .cin(t_9884), .o(t_9885), .co(t_9886), .cout(t_9887));
compressor_4_2 u2_3427(.a(t_6726), .b(t_6723), .c(t_6720), .d(t_6739), .cin(t_6736), .o(t_9888), .co(t_9889), .cout(t_9890));
compressor_4_2 u2_3428(.a(t_6747), .b(t_6744), .c(t_6741), .d(t_9887), .cin(t_9890), .o(t_9891), .co(t_9892), .cout(t_9893));
compressor_3_2 u1_3429(.a(t_6734), .b(t_6731), .cin(t_6750), .o(t_9894), .cout(t_9895));
compressor_4_2 u2_3430(.a(t_6758), .b(t_6755), .c(t_6752), .d(t_9893), .cin(t_9895), .o(t_9896), .co(t_9897), .cout(t_9898));
compressor_3_2 u1_3431(.a(t_6745), .b(t_6742), .cin(t_6761), .o(t_9899), .cout(t_9900));
compressor_4_2 u2_3432(.a(t_6766), .b(t_6763), .c(t_633), .d(t_9898), .cin(t_9900), .o(t_9901), .co(t_9902), .cout(t_9903));
compressor_4_2 u2_3433(.a(t_6759), .b(t_6756), .c(t_6753), .d(t_6772), .cin(t_6769), .o(t_9904), .co(t_9905), .cout(t_9906));
compressor_4_2 u2_3434(.a(t_6777), .b(t_6774), .c(t_654), .d(t_9903), .cin(t_9906), .o(t_9907), .co(t_9908), .cout(t_9909));
compressor_4_2 u2_3435(.a(t_6770), .b(t_6767), .c(t_6764), .d(t_6783), .cin(t_6780), .o(t_9910), .co(t_9911), .cout(t_9912));
compressor_4_2 u2_3436(.a(t_6791), .b(t_6788), .c(t_6785), .d(t_9909), .cin(t_9912), .o(t_9913), .co(t_9914), .cout(t_9915));
compressor_3_2 u1_3437(.a(t_6778), .b(t_6775), .cin(t_6794), .o(t_9916), .cout(t_9917));
compressor_4_2 u2_3438(.a(t_6800), .b(t_6797), .c(t_700), .d(t_9915), .cin(t_9917), .o(t_9918), .co(t_9919), .cout(t_9920));
compressor_4_2 u2_3439(.a(t_6792), .b(t_6789), .c(t_6786), .d(t_6806), .cin(t_6803), .o(t_9921), .co(t_9922), .cout(t_9923));
compressor_4_2 u2_3440(.a(t_6811), .b(t_6808), .c(t_723), .d(t_9920), .cin(t_9923), .o(t_9924), .co(t_9925), .cout(t_9926));
compressor_4_2 u2_3441(.a(t_6804), .b(t_6801), .c(t_6798), .d(t_6817), .cin(t_6814), .o(t_9927), .co(t_9928), .cout(t_9929));
compressor_4_2 u2_3442(.a(t_6822), .b(t_6819), .c(t_749), .d(t_9926), .cin(t_9929), .o(t_9930), .co(t_9931), .cout(t_9932));
compressor_4_2 u2_3443(.a(t_6815), .b(t_6812), .c(t_6809), .d(t_6828), .cin(t_6825), .o(t_9933), .co(t_9934), .cout(t_9935));
compressor_4_2 u2_3444(.a(t_6837), .b(t_6834), .c(t_6831), .d(t_9932), .cin(t_9935), .o(t_9936), .co(t_9937), .cout(t_9938));
compressor_4_2 u2_3445(.a(t_6829), .b(t_6826), .c(t_6823), .d(t_6820), .cin(t_6840), .o(t_9939), .co(t_9940), .cout(t_9941));
compressor_4_2 u2_3446(.a(t_6849), .b(t_6846), .c(t_6843), .d(t_9938), .cin(t_9941), .o(t_9942), .co(t_9943), .cout(t_9944));
compressor_4_2 u2_3447(.a(t_6841), .b(t_6838), .c(t_6835), .d(t_6832), .cin(t_6852), .o(t_9945), .co(t_9946), .cout(t_9947));
compressor_4_2 u2_3448(.a(t_6858), .b(t_6855), .c(t_820), .d(t_9944), .cin(t_9947), .o(t_9948), .co(t_9949), .cout(t_9950));
compressor_4_2 u2_3449(.a(t_6850), .b(t_6847), .c(t_6844), .d(t_6864), .cin(t_6861), .o(t_9951), .co(t_9952), .cout(t_9953));
compressor_4_2 u2_3450(.a(t_6870), .b(t_6867), .c(t_844), .d(t_9950), .cin(t_9953), .o(t_9954), .co(t_9955), .cout(t_9956));
compressor_4_2 u2_3451(.a(t_6862), .b(t_6859), .c(t_6856), .d(t_6876), .cin(t_6873), .o(t_9957), .co(t_9958), .cout(t_9959));
compressor_4_2 u2_3452(.a(t_6885), .b(t_6882), .c(t_6879), .d(t_9956), .cin(t_9959), .o(t_9960), .co(t_9961), .cout(t_9962));
compressor_4_2 u2_3453(.a(t_6874), .b(t_6871), .c(t_6868), .d(t_6891), .cin(t_6888), .o(t_9963), .co(t_9964), .cout(t_9965));
compressor_4_2 u2_3454(.a(t_6899), .b(t_6896), .c(t_6893), .d(t_9962), .cin(t_9965), .o(t_9966), .co(t_9967), .cout(t_9968));
compressor_4_2 u2_3455(.a(t_6886), .b(t_6883), .c(t_6880), .d(t_6905), .cin(t_6902), .o(t_9969), .co(t_9970), .cout(t_9971));
compressor_4_2 u2_3456(.a(t_6913), .b(t_6910), .c(t_6907), .d(t_9968), .cin(t_9971), .o(t_9972), .co(t_9973), .cout(t_9974));
compressor_4_2 u2_3457(.a(t_6900), .b(t_6897), .c(t_6894), .d(t_6919), .cin(t_6916), .o(t_9975), .co(t_9976), .cout(t_9977));
compressor_4_2 u2_3458(.a(t_6924), .b(t_6921), .c(t_951), .d(t_9974), .cin(t_9977), .o(t_9978), .co(t_9979), .cout(t_9980));
compressor_4_2 u2_3459(.a(t_6911), .b(t_6908), .c(t_6933), .d(t_6930), .cin(t_6927), .o(t_9981), .co(t_9982), .cout(t_9983));
half_adder u0_3460(.a(t_6917), .b(t_6914), .o(t_9984), .cout(t_9985));
compressor_4_2 u2_3461(.a(t_6941), .b(t_6938), .c(t_6935), .d(t_9980), .cin(t_9983), .o(t_9986), .co(t_9987), .cout(t_9988));
compressor_4_2 u2_3462(.a(t_6925), .b(t_6922), .c(t_6947), .d(t_6944), .cin(t_9985), .o(t_9989), .co(t_9990), .cout(t_9991));
half_adder u0_3463(.a(t_6931), .b(t_6928), .o(t_9992), .cout(t_9993));
compressor_4_2 u2_3464(.a(t_6955), .b(t_6952), .c(t_6949), .d(t_9988), .cin(t_9991), .o(t_9994), .co(t_9995), .cout(t_9996));
compressor_4_2 u2_3465(.a(t_6939), .b(t_6936), .c(t_6961), .d(t_6958), .cin(t_9993), .o(t_9997), .co(t_9998), .cout(t_9999));
half_adder u0_3466(.a(t_6945), .b(t_6942), .o(t_10000), .cout(t_10001));
compressor_4_2 u2_3467(.a(t_6966), .b(t_6963), .c(t_1031), .d(t_9996), .cin(t_9999), .o(t_10002), .co(t_10003), .cout(t_10004));
compressor_4_2 u2_3468(.a(t_6950), .b(t_6975), .c(t_6972), .d(t_6969), .cin(t_10001), .o(t_10005), .co(t_10006), .cout(t_10007));
compressor_3_2 u1_3469(.a(t_6959), .b(t_6956), .cin(t_6953), .o(t_10008), .cout(t_10009));
compressor_4_2 u2_3470(.a(t_6980), .b(t_6977), .c(t_1058), .d(t_10004), .cin(t_10007), .o(t_10010), .co(t_10011), .cout(t_10012));
compressor_4_2 u2_3471(.a(t_6964), .b(t_6989), .c(t_6986), .d(t_6983), .cin(t_10009), .o(t_10013), .co(t_10014), .cout(t_10015));
compressor_3_2 u1_3472(.a(t_6973), .b(t_6970), .cin(t_6967), .o(t_10016), .cout(t_10017));
compressor_4_2 u2_3473(.a(t_6997), .b(t_6994), .c(t_6991), .d(t_10012), .cin(t_10015), .o(t_10018), .co(t_10019), .cout(t_10020));
compressor_4_2 u2_3474(.a(t_6981), .b(t_6978), .c(t_7003), .d(t_7000), .cin(t_10017), .o(t_10021), .co(t_10022), .cout(t_10023));
half_adder u0_3475(.a(t_6987), .b(t_6984), .o(t_10024), .cout(t_10025));
compressor_4_2 u2_3476(.a(t_7009), .b(t_7006), .c(t_1116), .d(t_10020), .cin(t_10023), .o(t_10026), .co(t_10027), .cout(t_10028));
compressor_4_2 u2_3477(.a(t_6992), .b(t_7018), .c(t_7015), .d(t_7012), .cin(t_10025), .o(t_10029), .co(t_10030), .cout(t_10031));
compressor_3_2 u1_3478(.a(t_7001), .b(t_6998), .cin(t_6995), .o(t_10032), .cout(t_10033));
compressor_4_2 u2_3479(.a(t_7023), .b(t_7020), .c(t_1145), .d(t_10028), .cin(t_10031), .o(t_10034), .co(t_10035), .cout(t_10036));
compressor_4_2 u2_3480(.a(t_7007), .b(t_7032), .c(t_7029), .d(t_7026), .cin(t_10033), .o(t_10037), .co(t_10038), .cout(t_10039));
compressor_3_2 u1_3481(.a(t_7016), .b(t_7013), .cin(t_7010), .o(t_10040), .cout(t_10041));
compressor_4_2 u2_3482(.a(t_7037), .b(t_7034), .c(t_1177), .d(t_10036), .cin(t_10039), .o(t_10042), .co(t_10043), .cout(t_10044));
compressor_4_2 u2_3483(.a(t_7021), .b(t_7046), .c(t_7043), .d(t_7040), .cin(t_10041), .o(t_10045), .co(t_10046), .cout(t_10047));
compressor_3_2 u1_3484(.a(t_7030), .b(t_7027), .cin(t_7024), .o(t_10048), .cout(t_10049));
compressor_4_2 u2_3485(.a(t_7055), .b(t_7052), .c(t_7049), .d(t_10044), .cin(t_10047), .o(t_10050), .co(t_10051), .cout(t_10052));
compressor_4_2 u2_3486(.a(t_7038), .b(t_7035), .c(t_7061), .d(t_7058), .cin(t_10049), .o(t_10053), .co(t_10054), .cout(t_10055));
compressor_3_2 u1_3487(.a(t_7047), .b(t_7044), .cin(t_7041), .o(t_10056), .cout(t_10057));
compressor_4_2 u2_3488(.a(t_7070), .b(t_7067), .c(t_7064), .d(t_10052), .cin(t_10055), .o(t_10058), .co(t_10059), .cout(t_10060));
compressor_4_2 u2_3489(.a(t_7053), .b(t_7050), .c(t_7076), .d(t_7073), .cin(t_10057), .o(t_10061), .co(t_10062), .cout(t_10063));
compressor_3_2 u1_3490(.a(t_7062), .b(t_7059), .cin(t_7056), .o(t_10064), .cout(t_10065));
compressor_4_2 u2_3491(.a(t_7082), .b(t_7079), .c(t_1266), .d(t_10060), .cin(t_10063), .o(t_10066), .co(t_10067), .cout(t_10068));
compressor_4_2 u2_3492(.a(t_7065), .b(t_7091), .c(t_7088), .d(t_7085), .cin(t_10065), .o(t_10069), .co(t_10070), .cout(t_10071));
compressor_3_2 u1_3493(.a(t_7074), .b(t_7071), .cin(t_7068), .o(t_10072), .cout(t_10073));
compressor_4_2 u2_3494(.a(t_7097), .b(t_7094), .c(t_1296), .d(t_10068), .cin(t_10071), .o(t_10074), .co(t_10075), .cout(t_10076));
compressor_4_2 u2_3495(.a(t_7080), .b(t_7106), .c(t_7103), .d(t_7100), .cin(t_10073), .o(t_10077), .co(t_10078), .cout(t_10079));
compressor_3_2 u1_3496(.a(t_7089), .b(t_7086), .cin(t_7083), .o(t_10080), .cout(t_10081));
compressor_4_2 u2_3497(.a(t_7115), .b(t_7112), .c(t_7109), .d(t_10076), .cin(t_10079), .o(t_10082), .co(t_10083), .cout(t_10084));
compressor_4_2 u2_3498(.a(t_7095), .b(t_7124), .c(t_7121), .d(t_7118), .cin(t_10081), .o(t_10085), .co(t_10086), .cout(t_10087));
compressor_3_2 u1_3499(.a(t_7104), .b(t_7101), .cin(t_7098), .o(t_10088), .cout(t_10089));
compressor_4_2 u2_3500(.a(t_7132), .b(t_7129), .c(t_7126), .d(t_10084), .cin(t_10087), .o(t_10090), .co(t_10091), .cout(t_10092));
compressor_4_2 u2_3501(.a(t_7110), .b(t_7141), .c(t_7138), .d(t_7135), .cin(t_10089), .o(t_10093), .co(t_10094), .cout(t_10095));
compressor_3_2 u1_3502(.a(t_7119), .b(t_7116), .cin(t_7113), .o(t_10096), .cout(t_10097));
compressor_4_2 u2_3503(.a(t_7149), .b(t_7146), .c(t_7143), .d(t_10092), .cin(t_10095), .o(t_10098), .co(t_10099), .cout(t_10100));
compressor_4_2 u2_3504(.a(t_7127), .b(t_7158), .c(t_7155), .d(t_7152), .cin(t_10097), .o(t_10101), .co(t_10102), .cout(t_10103));
compressor_3_2 u1_3505(.a(t_7136), .b(t_7133), .cin(t_7130), .o(t_10104), .cout(t_10105));
compressor_4_2 u2_3506(.a(t_7163), .b(t_7160), .c(t_1427), .d(t_10100), .cin(t_10103), .o(t_10106), .co(t_10107), .cout(t_10108));
compressor_4_2 u2_3507(.a(t_7175), .b(t_7172), .c(t_7169), .d(t_7166), .cin(t_10105), .o(t_10109), .co(t_10110), .cout(t_10111));
compressor_4_2 u2_3508(.a(t_7156), .b(t_7153), .c(t_7150), .d(t_7147), .cin(t_7144), .o(t_10112), .co(t_10113), .cout(t_10114));
compressor_4_2 u2_3509(.a(t_7183), .b(t_7180), .c(t_7177), .d(t_10108), .cin(t_10111), .o(t_10115), .co(t_10116), .cout(t_10117));
compressor_4_2 u2_3510(.a(t_7161), .b(t_7192), .c(t_7189), .d(t_7186), .cin(t_10114), .o(t_10118), .co(t_10119), .cout(t_10120));
compressor_3_2 u1_3511(.a(t_7170), .b(t_7167), .cin(t_7164), .o(t_10121), .cout(t_10122));
compressor_4_2 u2_3512(.a(t_7200), .b(t_7197), .c(t_7194), .d(t_10117), .cin(t_10120), .o(t_10123), .co(t_10124), .cout(t_10125));
compressor_4_2 u2_3513(.a(t_7178), .b(t_7209), .c(t_7206), .d(t_7203), .cin(t_10122), .o(t_10126), .co(t_10127), .cout(t_10128));
compressor_3_2 u1_3514(.a(t_7187), .b(t_7184), .cin(t_7181), .o(t_10129), .cout(t_10130));
compressor_4_2 u2_3515(.a(t_7214), .b(t_7211), .c(t_1525), .d(t_10125), .cin(t_10128), .o(t_10131), .co(t_10132), .cout(t_10133));
compressor_4_2 u2_3516(.a(t_7226), .b(t_7223), .c(t_7220), .d(t_7217), .cin(t_10130), .o(t_10134), .co(t_10135), .cout(t_10136));
compressor_4_2 u2_3517(.a(t_7207), .b(t_7204), .c(t_7201), .d(t_7198), .cin(t_7195), .o(t_10137), .co(t_10138), .cout(t_10139));
compressor_4_2 u2_3518(.a(t_7231), .b(t_7228), .c(t_1558), .d(t_10133), .cin(t_10136), .o(t_10140), .co(t_10141), .cout(t_10142));
compressor_4_2 u2_3519(.a(t_7243), .b(t_7240), .c(t_7237), .d(t_7234), .cin(t_10139), .o(t_10143), .co(t_10144), .cout(t_10145));
compressor_4_2 u2_3520(.a(t_7224), .b(t_7221), .c(t_7218), .d(t_7215), .cin(t_7212), .o(t_10146), .co(t_10147), .cout(t_10148));
compressor_4_2 u2_3521(.a(t_7251), .b(t_7248), .c(t_7245), .d(t_10142), .cin(t_10145), .o(t_10149), .co(t_10150), .cout(t_10151));
compressor_4_2 u2_3522(.a(t_7229), .b(t_7260), .c(t_7257), .d(t_7254), .cin(t_10148), .o(t_10152), .co(t_10153), .cout(t_10154));
compressor_3_2 u1_3523(.a(t_7238), .b(t_7235), .cin(t_7232), .o(t_10155), .cout(t_10156));
compressor_4_2 u2_3524(.a(t_7266), .b(t_7263), .c(t_1628), .d(t_10151), .cin(t_10154), .o(t_10157), .co(t_10158), .cout(t_10159));
compressor_4_2 u2_3525(.a(t_7278), .b(t_7275), .c(t_7272), .d(t_7269), .cin(t_10156), .o(t_10160), .co(t_10161), .cout(t_10162));
compressor_4_2 u2_3526(.a(t_7258), .b(t_7255), .c(t_7252), .d(t_7249), .cin(t_7246), .o(t_10163), .co(t_10164), .cout(t_10165));
compressor_4_2 u2_3527(.a(t_7283), .b(t_7280), .c(t_1663), .d(t_10159), .cin(t_10162), .o(t_10166), .co(t_10167), .cout(t_10168));
compressor_4_2 u2_3528(.a(t_7295), .b(t_7292), .c(t_7289), .d(t_7286), .cin(t_10165), .o(t_10169), .co(t_10170), .cout(t_10171));
compressor_4_2 u2_3529(.a(t_7276), .b(t_7273), .c(t_7270), .d(t_7267), .cin(t_7264), .o(t_10172), .co(t_10173), .cout(t_10174));
compressor_4_2 u2_3530(.a(t_7300), .b(t_7297), .c(t_1701), .d(t_10168), .cin(t_10171), .o(t_10175), .co(t_10176), .cout(t_10177));
compressor_4_2 u2_3531(.a(t_7312), .b(t_7309), .c(t_7306), .d(t_7303), .cin(t_10174), .o(t_10178), .co(t_10179), .cout(t_10180));
compressor_4_2 u2_3532(.a(t_7293), .b(t_7290), .c(t_7287), .d(t_7284), .cin(t_7281), .o(t_10181), .co(t_10182), .cout(t_10183));
compressor_4_2 u2_3533(.a(t_7321), .b(t_7318), .c(t_7315), .d(t_10177), .cin(t_10180), .o(t_10184), .co(t_10185), .cout(t_10186));
compressor_4_2 u2_3534(.a(t_7298), .b(t_7330), .c(t_7327), .d(t_7324), .cin(t_10183), .o(t_10187), .co(t_10188), .cout(t_10189));
compressor_4_2 u2_3535(.a(t_7313), .b(t_7310), .c(t_7307), .d(t_7304), .cin(t_7301), .o(t_10190), .co(t_10191), .cout(t_10192));
compressor_4_2 u2_3536(.a(t_7339), .b(t_7336), .c(t_7333), .d(t_10186), .cin(t_10189), .o(t_10193), .co(t_10194), .cout(t_10195));
compressor_4_2 u2_3537(.a(t_7316), .b(t_7348), .c(t_7345), .d(t_7342), .cin(t_10192), .o(t_10196), .co(t_10197), .cout(t_10198));
compressor_4_2 u2_3538(.a(t_7331), .b(t_7328), .c(t_7325), .d(t_7322), .cin(t_7319), .o(t_10199), .co(t_10200), .cout(t_10201));
compressor_4_2 u2_3539(.a(t_7354), .b(t_7351), .c(t_1808), .d(t_10195), .cin(t_10198), .o(t_10202), .co(t_10203), .cout(t_10204));
compressor_4_2 u2_3540(.a(t_7366), .b(t_7363), .c(t_7360), .d(t_7357), .cin(t_10201), .o(t_10205), .co(t_10206), .cout(t_10207));
compressor_4_2 u2_3541(.a(t_7346), .b(t_7343), .c(t_7340), .d(t_7337), .cin(t_7334), .o(t_10208), .co(t_10209), .cout(t_10210));
compressor_4_2 u2_3542(.a(t_7372), .b(t_7369), .c(t_1844), .d(t_10204), .cin(t_10207), .o(t_10211), .co(t_10212), .cout(t_10213));
compressor_4_2 u2_3543(.a(t_7384), .b(t_7381), .c(t_7378), .d(t_7375), .cin(t_10210), .o(t_10214), .co(t_10215), .cout(t_10216));
compressor_4_2 u2_3544(.a(t_7364), .b(t_7361), .c(t_7358), .d(t_7355), .cin(t_7352), .o(t_10217), .co(t_10218), .cout(t_10219));
compressor_4_2 u2_3545(.a(t_7393), .b(t_7390), .c(t_7387), .d(t_10213), .cin(t_10216), .o(t_10220), .co(t_10221), .cout(t_10222));
compressor_4_2 u2_3546(.a(t_7405), .b(t_7402), .c(t_7399), .d(t_7396), .cin(t_10219), .o(t_10223), .co(t_10224), .cout(t_10225));
compressor_4_2 u2_3547(.a(t_7382), .b(t_7379), .c(t_7376), .d(t_7373), .cin(t_7370), .o(t_10226), .co(t_10227), .cout(t_10228));
compressor_4_2 u2_3548(.a(t_7413), .b(t_7410), .c(t_7407), .d(t_10222), .cin(t_10225), .o(t_10229), .co(t_10230), .cout(t_10231));
compressor_4_2 u2_3549(.a(t_7425), .b(t_7422), .c(t_7419), .d(t_7416), .cin(t_10228), .o(t_10232), .co(t_10233), .cout(t_10234));
compressor_4_2 u2_3550(.a(t_7400), .b(t_7397), .c(t_7394), .d(t_7391), .cin(t_7388), .o(t_10235), .co(t_10236), .cout(t_10237));
compressor_4_2 u2_3551(.a(t_7433), .b(t_7430), .c(t_7427), .d(t_10231), .cin(t_10234), .o(t_10238), .co(t_10239), .cout(t_10240));
compressor_4_2 u2_3552(.a(t_7445), .b(t_7442), .c(t_7439), .d(t_7436), .cin(t_10237), .o(t_10241), .co(t_10242), .cout(t_10243));
compressor_4_2 u2_3553(.a(t_7420), .b(t_7417), .c(t_7414), .d(t_7411), .cin(t_7408), .o(t_10244), .co(t_10245), .cout(t_10246));
compressor_4_2 u2_3554(.a(t_7450), .b(t_7447), .c(t_1999), .d(t_10240), .cin(t_10243), .o(t_10247), .co(t_10248), .cout(t_10249));
compressor_4_2 u2_3555(.a(t_7462), .b(t_7459), .c(t_7456), .d(t_7453), .cin(t_10246), .o(t_10250), .co(t_10251), .cout(t_10252));
compressor_4_2 u2_3556(.a(t_7437), .b(t_7434), .c(t_7431), .d(t_7428), .cin(t_7465), .o(t_10253), .co(t_10254), .cout(t_10255));
half_adder u0_3557(.a(t_7443), .b(t_7440), .o(t_10256), .cout(t_10257));
compressor_4_2 u2_3558(.a(t_7473), .b(t_7470), .c(t_7467), .d(t_10249), .cin(t_10252), .o(t_10258), .co(t_10259), .cout(t_10260));
compressor_4_2 u2_3559(.a(t_7482), .b(t_7479), .c(t_7476), .d(t_10255), .cin(t_10257), .o(t_10261), .co(t_10262), .cout(t_10263));
compressor_4_2 u2_3560(.a(t_7457), .b(t_7454), .c(t_7451), .d(t_7448), .cin(t_7485), .o(t_10264), .co(t_10265), .cout(t_10266));
half_adder u0_3561(.a(t_7463), .b(t_7460), .o(t_10267), .cout(t_10268));
compressor_4_2 u2_3562(.a(t_7493), .b(t_7490), .c(t_7487), .d(t_10260), .cin(t_10263), .o(t_10269), .co(t_10270), .cout(t_10271));
compressor_4_2 u2_3563(.a(t_7502), .b(t_7499), .c(t_7496), .d(t_10266), .cin(t_10268), .o(t_10272), .co(t_10273), .cout(t_10274));
compressor_4_2 u2_3564(.a(t_7477), .b(t_7474), .c(t_7471), .d(t_7468), .cin(t_7505), .o(t_10275), .co(t_10276), .cout(t_10277));
half_adder u0_3565(.a(t_7483), .b(t_7480), .o(t_10278), .cout(t_10279));
compressor_4_2 u2_3566(.a(t_7510), .b(t_7507), .c(t_2115), .d(t_10271), .cin(t_10274), .o(t_10280), .co(t_10281), .cout(t_10282));
compressor_4_2 u2_3567(.a(t_7519), .b(t_7516), .c(t_7513), .d(t_10277), .cin(t_10279), .o(t_10283), .co(t_10284), .cout(t_10285));
compressor_4_2 u2_3568(.a(t_7494), .b(t_7491), .c(t_7488), .d(t_7525), .cin(t_7522), .o(t_10286), .co(t_10287), .cout(t_10288));
compressor_3_2 u1_3569(.a(t_7503), .b(t_7500), .cin(t_7497), .o(t_10289), .cout(t_10290));
compressor_4_2 u2_3570(.a(t_7530), .b(t_7527), .c(t_2154), .d(t_10282), .cin(t_10285), .o(t_10291), .co(t_10292), .cout(t_10293));
compressor_4_2 u2_3571(.a(t_7539), .b(t_7536), .c(t_7533), .d(t_10288), .cin(t_10290), .o(t_10294), .co(t_10295), .cout(t_10296));
compressor_4_2 u2_3572(.a(t_7514), .b(t_7511), .c(t_7508), .d(t_7545), .cin(t_7542), .o(t_10297), .co(t_10298), .cout(t_10299));
compressor_3_2 u1_3573(.a(t_7523), .b(t_7520), .cin(t_7517), .o(t_10300), .cout(t_10301));
compressor_4_2 u2_3574(.a(t_7553), .b(t_7550), .c(t_7547), .d(t_10293), .cin(t_10296), .o(t_10302), .co(t_10303), .cout(t_10304));
compressor_4_2 u2_3575(.a(t_7562), .b(t_7559), .c(t_7556), .d(t_10299), .cin(t_10301), .o(t_10305), .co(t_10306), .cout(t_10307));
compressor_4_2 u2_3576(.a(t_7537), .b(t_7534), .c(t_7531), .d(t_7528), .cin(t_7565), .o(t_10308), .co(t_10309), .cout(t_10310));
half_adder u0_3577(.a(t_7543), .b(t_7540), .o(t_10311), .cout(t_10312));
compressor_4_2 u2_3578(.a(t_7571), .b(t_7568), .c(t_2236), .d(t_10304), .cin(t_10307), .o(t_10313), .co(t_10314), .cout(t_10315));
compressor_4_2 u2_3579(.a(t_7580), .b(t_7577), .c(t_7574), .d(t_10310), .cin(t_10312), .o(t_10316), .co(t_10317), .cout(t_10318));
compressor_4_2 u2_3580(.a(t_7554), .b(t_7551), .c(t_7548), .d(t_7586), .cin(t_7583), .o(t_10319), .co(t_10320), .cout(t_10321));
compressor_3_2 u1_3581(.a(t_7563), .b(t_7560), .cin(t_7557), .o(t_10322), .cout(t_10323));
compressor_4_2 u2_3582(.a(t_7591), .b(t_7588), .c(t_2277), .d(t_10315), .cin(t_10318), .o(t_10324), .co(t_10325), .cout(t_10326));
compressor_4_2 u2_3583(.a(t_7600), .b(t_7597), .c(t_7594), .d(t_10321), .cin(t_10323), .o(t_10327), .co(t_10328), .cout(t_10329));
compressor_4_2 u2_3584(.a(t_7575), .b(t_7572), .c(t_7569), .d(t_7606), .cin(t_7603), .o(t_10330), .co(t_10331), .cout(t_10332));
compressor_3_2 u1_3585(.a(t_7584), .b(t_7581), .cin(t_7578), .o(t_10333), .cout(t_10334));
compressor_4_2 u2_3586(.a(t_7611), .b(t_7608), .c(t_2321), .d(t_10326), .cin(t_10329), .o(t_10335), .co(t_10336), .cout(t_10337));
compressor_4_2 u2_3587(.a(t_7620), .b(t_7617), .c(t_7614), .d(t_10332), .cin(t_10334), .o(t_10338), .co(t_10339), .cout(t_10340));
compressor_4_2 u2_3588(.a(t_7595), .b(t_7592), .c(t_7589), .d(t_7626), .cin(t_7623), .o(t_10341), .co(t_10342), .cout(t_10343));
compressor_3_2 u1_3589(.a(t_7604), .b(t_7601), .cin(t_7598), .o(t_10344), .cout(t_10345));
compressor_4_2 u2_3590(.a(t_7635), .b(t_7632), .c(t_7629), .d(t_10337), .cin(t_10340), .o(t_10346), .co(t_10347), .cout(t_10348));
compressor_4_2 u2_3591(.a(t_7644), .b(t_7641), .c(t_7638), .d(t_10343), .cin(t_10345), .o(t_10349), .co(t_10350), .cout(t_10351));
compressor_4_2 u2_3592(.a(t_7618), .b(t_7615), .c(t_7612), .d(t_7609), .cin(t_7647), .o(t_10352), .co(t_10353), .cout(t_10354));
compressor_3_2 u1_3593(.a(t_7627), .b(t_7624), .cin(t_7621), .o(t_10355), .cout(t_10356));
compressor_4_2 u2_3594(.a(t_7656), .b(t_7653), .c(t_7650), .d(t_10348), .cin(t_10351), .o(t_10357), .co(t_10358), .cout(t_10359));
compressor_4_2 u2_3595(.a(t_7665), .b(t_7662), .c(t_7659), .d(t_10354), .cin(t_10356), .o(t_10360), .co(t_10361), .cout(t_10362));
compressor_4_2 u2_3596(.a(t_7639), .b(t_7636), .c(t_7633), .d(t_7630), .cin(t_7668), .o(t_10363), .co(t_10364), .cout(t_10365));
compressor_3_2 u1_3597(.a(t_7648), .b(t_7645), .cin(t_7642), .o(t_10366), .cout(t_10367));
compressor_4_2 u2_3598(.a(t_7674), .b(t_7671), .c(t_2446), .d(t_10359), .cin(t_10362), .o(t_10368), .co(t_10369), .cout(t_10370));
compressor_4_2 u2_3599(.a(t_7683), .b(t_7680), .c(t_7677), .d(t_10365), .cin(t_10367), .o(t_10371), .co(t_10372), .cout(t_10373));
compressor_4_2 u2_3600(.a(t_7657), .b(t_7654), .c(t_7651), .d(t_7689), .cin(t_7686), .o(t_10374), .co(t_10375), .cout(t_10376));
compressor_3_2 u1_3601(.a(t_7666), .b(t_7663), .cin(t_7660), .o(t_10377), .cout(t_10378));
compressor_4_2 u2_3602(.a(t_7695), .b(t_7692), .c(t_2488), .d(t_10370), .cin(t_10373), .o(t_10379), .co(t_10380), .cout(t_10381));
compressor_4_2 u2_3603(.a(t_7704), .b(t_7701), .c(t_7698), .d(t_10376), .cin(t_10378), .o(t_10382), .co(t_10383), .cout(t_10384));
compressor_4_2 u2_3604(.a(t_7678), .b(t_7675), .c(t_7672), .d(t_7710), .cin(t_7707), .o(t_10385), .co(t_10386), .cout(t_10387));
compressor_3_2 u1_3605(.a(t_7687), .b(t_7684), .cin(t_7681), .o(t_10388), .cout(t_10389));
compressor_4_2 u2_3606(.a(t_7719), .b(t_7716), .c(t_7713), .d(t_10381), .cin(t_10384), .o(t_10390), .co(t_10391), .cout(t_10392));
compressor_4_2 u2_3607(.a(t_7728), .b(t_7725), .c(t_7722), .d(t_10387), .cin(t_10389), .o(t_10393), .co(t_10394), .cout(t_10395));
compressor_4_2 u2_3608(.a(t_7699), .b(t_7696), .c(t_7693), .d(t_7734), .cin(t_7731), .o(t_10396), .co(t_10397), .cout(t_10398));
compressor_3_2 u1_3609(.a(t_7708), .b(t_7705), .cin(t_7702), .o(t_10399), .cout(t_10400));
compressor_4_2 u2_3610(.a(t_7742), .b(t_7739), .c(t_7736), .d(t_10392), .cin(t_10395), .o(t_10401), .co(t_10402), .cout(t_10403));
compressor_4_2 u2_3611(.a(t_7751), .b(t_7748), .c(t_7745), .d(t_10398), .cin(t_10400), .o(t_10404), .co(t_10405), .cout(t_10406));
compressor_4_2 u2_3612(.a(t_7720), .b(t_7717), .c(t_7714), .d(t_7757), .cin(t_7754), .o(t_10407), .co(t_10408), .cout(t_10409));
compressor_3_2 u1_3613(.a(t_7729), .b(t_7726), .cin(t_7723), .o(t_10410), .cout(t_10411));
compressor_4_2 u2_3614(.a(t_7765), .b(t_7762), .c(t_7759), .d(t_10403), .cin(t_10406), .o(t_10412), .co(t_10413), .cout(t_10414));
compressor_4_2 u2_3615(.a(t_7774), .b(t_7771), .c(t_7768), .d(t_10409), .cin(t_10411), .o(t_10415), .co(t_10416), .cout(t_10417));
compressor_4_2 u2_3616(.a(t_7743), .b(t_7740), .c(t_7737), .d(t_7780), .cin(t_7777), .o(t_10418), .co(t_10419), .cout(t_10420));
compressor_3_2 u1_3617(.a(t_7752), .b(t_7749), .cin(t_7746), .o(t_10421), .cout(t_10422));
compressor_4_2 u2_3618(.a(t_7785), .b(t_7782), .c(t_2667), .d(t_10414), .cin(t_10417), .o(t_10423), .co(t_10424), .cout(t_10425));
compressor_4_2 u2_3619(.a(t_7794), .b(t_7791), .c(t_7788), .d(t_10420), .cin(t_10422), .o(t_10426), .co(t_10427), .cout(t_10428));
compressor_4_2 u2_3620(.a(t_7763), .b(t_7760), .c(t_7803), .d(t_7800), .cin(t_7797), .o(t_10429), .co(t_10430), .cout(t_10431));
compressor_4_2 u2_3621(.a(t_7778), .b(t_7775), .c(t_7772), .d(t_7769), .cin(t_7766), .o(t_10432), .co(t_10433), .cout(t_10434));
compressor_4_2 u2_3622(.a(t_7811), .b(t_7808), .c(t_7805), .d(t_10425), .cin(t_10428), .o(t_10435), .co(t_10436), .cout(t_10437));
compressor_4_2 u2_3623(.a(t_7820), .b(t_7817), .c(t_7814), .d(t_10431), .cin(t_10434), .o(t_10438), .co(t_10439), .cout(t_10440));
compressor_4_2 u2_3624(.a(t_7789), .b(t_7786), .c(t_7783), .d(t_7826), .cin(t_7823), .o(t_10441), .co(t_10442), .cout(t_10443));
compressor_3_2 u1_3625(.a(t_7798), .b(t_7795), .cin(t_7792), .o(t_10444), .cout(t_10445));
compressor_4_2 u2_3626(.a(t_7834), .b(t_7831), .c(t_7828), .d(t_10437), .cin(t_10440), .o(t_10446), .co(t_10447), .cout(t_10448));
compressor_4_2 u2_3627(.a(t_7843), .b(t_7840), .c(t_7837), .d(t_10443), .cin(t_10445), .o(t_10449), .co(t_10450), .cout(t_10451));
compressor_4_2 u2_3628(.a(t_7812), .b(t_7809), .c(t_7806), .d(t_7849), .cin(t_7846), .o(t_10452), .co(t_10453), .cout(t_10454));
compressor_3_2 u1_3629(.a(t_7821), .b(t_7818), .cin(t_7815), .o(t_10455), .cout(t_10456));
compressor_4_2 u2_3630(.a(t_7854), .b(t_7851), .c(t_2801), .d(t_10448), .cin(t_10451), .o(t_10457), .co(t_10458), .cout(t_10459));
compressor_4_2 u2_3631(.a(t_7863), .b(t_7860), .c(t_7857), .d(t_10454), .cin(t_10456), .o(t_10460), .co(t_10461), .cout(t_10462));
compressor_4_2 u2_3632(.a(t_7832), .b(t_7829), .c(t_7872), .d(t_7869), .cin(t_7866), .o(t_10463), .co(t_10464), .cout(t_10465));
compressor_4_2 u2_3633(.a(t_7847), .b(t_7844), .c(t_7841), .d(t_7838), .cin(t_7835), .o(t_10466), .co(t_10467), .cout(t_10468));
compressor_4_2 u2_3634(.a(t_7877), .b(t_7874), .c(t_2846), .d(t_10459), .cin(t_10462), .o(t_10469), .co(t_10470), .cout(t_10471));
compressor_4_2 u2_3635(.a(t_7886), .b(t_7883), .c(t_7880), .d(t_10465), .cin(t_10468), .o(t_10472), .co(t_10473), .cout(t_10474));
compressor_4_2 u2_3636(.a(t_7855), .b(t_7852), .c(t_7895), .d(t_7892), .cin(t_7889), .o(t_10475), .co(t_10476), .cout(t_10477));
compressor_4_2 u2_3637(.a(t_7870), .b(t_7867), .c(t_7864), .d(t_7861), .cin(t_7858), .o(t_10478), .co(t_10479), .cout(t_10480));
compressor_4_2 u2_3638(.a(t_7903), .b(t_7900), .c(t_7897), .d(t_10471), .cin(t_10474), .o(t_10481), .co(t_10482), .cout(t_10483));
compressor_4_2 u2_3639(.a(t_7912), .b(t_7909), .c(t_7906), .d(t_10477), .cin(t_10480), .o(t_10484), .co(t_10485), .cout(t_10486));
compressor_4_2 u2_3640(.a(t_7881), .b(t_7878), .c(t_7875), .d(t_7918), .cin(t_7915), .o(t_10487), .co(t_10488), .cout(t_10489));
compressor_3_2 u1_3641(.a(t_7890), .b(t_7887), .cin(t_7884), .o(t_10490), .cout(t_10491));
compressor_4_2 u2_3642(.a(t_7924), .b(t_7921), .c(t_2940), .d(t_10483), .cin(t_10486), .o(t_10492), .co(t_10493), .cout(t_10494));
compressor_4_2 u2_3643(.a(t_7933), .b(t_7930), .c(t_7927), .d(t_10489), .cin(t_10491), .o(t_10495), .co(t_10496), .cout(t_10497));
compressor_4_2 u2_3644(.a(t_7901), .b(t_7898), .c(t_7942), .d(t_7939), .cin(t_7936), .o(t_10498), .co(t_10499), .cout(t_10500));
compressor_4_2 u2_3645(.a(t_7916), .b(t_7913), .c(t_7910), .d(t_7907), .cin(t_7904), .o(t_10501), .co(t_10502), .cout(t_10503));
compressor_4_2 u2_3646(.a(t_7947), .b(t_7944), .c(t_2987), .d(t_10494), .cin(t_10497), .o(t_10504), .co(t_10505), .cout(t_10506));
compressor_4_2 u2_3647(.a(t_7956), .b(t_7953), .c(t_7950), .d(t_10500), .cin(t_10503), .o(t_10507), .co(t_10508), .cout(t_10509));
compressor_4_2 u2_3648(.a(t_7925), .b(t_7922), .c(t_7965), .d(t_7962), .cin(t_7959), .o(t_10510), .co(t_10511), .cout(t_10512));
compressor_4_2 u2_3649(.a(t_7940), .b(t_7937), .c(t_7934), .d(t_7931), .cin(t_7928), .o(t_10513), .co(t_10514), .cout(t_10515));
compressor_4_2 u2_3650(.a(t_7970), .b(t_7967), .c(t_3037), .d(t_10506), .cin(t_10509), .o(t_10516), .co(t_10517), .cout(t_10518));
compressor_4_2 u2_3651(.a(t_7979), .b(t_7976), .c(t_7973), .d(t_10512), .cin(t_10515), .o(t_10519), .co(t_10520), .cout(t_10521));
compressor_4_2 u2_3652(.a(t_7948), .b(t_7945), .c(t_7988), .d(t_7985), .cin(t_7982), .o(t_10522), .co(t_10523), .cout(t_10524));
compressor_4_2 u2_3653(.a(t_7963), .b(t_7960), .c(t_7957), .d(t_7954), .cin(t_7951), .o(t_10525), .co(t_10526), .cout(t_10527));
compressor_4_2 u2_3654(.a(t_7997), .b(t_7994), .c(t_7991), .d(t_10518), .cin(t_10521), .o(t_10528), .co(t_10529), .cout(t_10530));
compressor_4_2 u2_3655(.a(t_8006), .b(t_8003), .c(t_8000), .d(t_10524), .cin(t_10527), .o(t_10531), .co(t_10532), .cout(t_10533));
compressor_4_2 u2_3656(.a(t_7974), .b(t_7971), .c(t_7968), .d(t_8012), .cin(t_8009), .o(t_10534), .co(t_10535), .cout(t_10536));
compressor_4_2 u2_3657(.a(t_7989), .b(t_7986), .c(t_7983), .d(t_7980), .cin(t_7977), .o(t_10537), .co(t_10538), .cout(t_10539));
compressor_4_2 u2_3658(.a(t_8021), .b(t_8018), .c(t_8015), .d(t_10530), .cin(t_10533), .o(t_10540), .co(t_10541), .cout(t_10542));
compressor_4_2 u2_3659(.a(t_8030), .b(t_8027), .c(t_8024), .d(t_10536), .cin(t_10539), .o(t_10543), .co(t_10544), .cout(t_10545));
compressor_4_2 u2_3660(.a(t_7998), .b(t_7995), .c(t_7992), .d(t_8036), .cin(t_8033), .o(t_10546), .co(t_10547), .cout(t_10548));
compressor_4_2 u2_3661(.a(t_8013), .b(t_8010), .c(t_8007), .d(t_8004), .cin(t_8001), .o(t_10549), .co(t_10550), .cout(t_10551));
compressor_4_2 u2_3662(.a(t_8042), .b(t_8039), .c(t_3180), .d(t_10542), .cin(t_10545), .o(t_10552), .co(t_10553), .cout(t_10554));
compressor_4_2 u2_3663(.a(t_8051), .b(t_8048), .c(t_8045), .d(t_10548), .cin(t_10551), .o(t_10555), .co(t_10556), .cout(t_10557));
compressor_4_2 u2_3664(.a(t_8019), .b(t_8016), .c(t_8060), .d(t_8057), .cin(t_8054), .o(t_10558), .co(t_10559), .cout(t_10560));
compressor_4_2 u2_3665(.a(t_8034), .b(t_8031), .c(t_8028), .d(t_8025), .cin(t_8022), .o(t_10561), .co(t_10562), .cout(t_10563));
compressor_4_2 u2_3666(.a(t_8066), .b(t_8063), .c(t_3228), .d(t_10554), .cin(t_10557), .o(t_10564), .co(t_10565), .cout(t_10566));
compressor_4_2 u2_3667(.a(t_8075), .b(t_8072), .c(t_8069), .d(t_10560), .cin(t_10563), .o(t_10567), .co(t_10568), .cout(t_10569));
compressor_4_2 u2_3668(.a(t_8043), .b(t_8040), .c(t_8084), .d(t_8081), .cin(t_8078), .o(t_10570), .co(t_10571), .cout(t_10572));
compressor_4_2 u2_3669(.a(t_8058), .b(t_8055), .c(t_8052), .d(t_8049), .cin(t_8046), .o(t_10573), .co(t_10574), .cout(t_10575));
compressor_4_2 u2_3670(.a(t_8093), .b(t_8090), .c(t_8087), .d(t_10566), .cin(t_10569), .o(t_10576), .co(t_10577), .cout(t_10578));
compressor_4_2 u2_3671(.a(t_8102), .b(t_8099), .c(t_8096), .d(t_10572), .cin(t_10575), .o(t_10579), .co(t_10580), .cout(t_10581));
compressor_4_2 u2_3672(.a(t_8070), .b(t_8067), .c(t_8064), .d(t_8108), .cin(t_8105), .o(t_10582), .co(t_10583), .cout(t_10584));
compressor_4_2 u2_3673(.a(t_8085), .b(t_8082), .c(t_8079), .d(t_8076), .cin(t_8073), .o(t_10585), .co(t_10586), .cout(t_10587));
compressor_4_2 u2_3674(.a(t_8117), .b(t_8114), .c(t_8111), .d(t_10578), .cin(t_10581), .o(t_10588), .co(t_10589), .cout(t_10590));
compressor_4_2 u2_3675(.a(t_8126), .b(t_8123), .c(t_8120), .d(t_10584), .cin(t_10587), .o(t_10591), .co(t_10592), .cout(t_10593));
compressor_4_2 u2_3676(.a(t_8094), .b(t_8091), .c(t_8088), .d(t_8132), .cin(t_8129), .o(t_10594), .co(t_10595), .cout(t_10596));
compressor_4_2 u2_3677(.a(t_8109), .b(t_8106), .c(t_8103), .d(t_8100), .cin(t_8097), .o(t_10597), .co(t_10598), .cout(t_10599));
compressor_4_2 u2_3678(.a(t_8138), .b(t_8135), .c(t_3372), .d(t_10590), .cin(t_10593), .o(t_10600), .co(t_10601), .cout(t_10602));
compressor_4_2 u2_3679(.a(t_8147), .b(t_8144), .c(t_8141), .d(t_10596), .cin(t_10599), .o(t_10603), .co(t_10604), .cout(t_10605));
compressor_4_2 u2_3680(.a(t_8115), .b(t_8112), .c(t_8156), .d(t_8153), .cin(t_8150), .o(t_10606), .co(t_10607), .cout(t_10608));
compressor_4_2 u2_3681(.a(t_8130), .b(t_8127), .c(t_8124), .d(t_8121), .cin(t_8118), .o(t_10609), .co(t_10610), .cout(t_10611));
compressor_4_2 u2_3682(.a(t_8165), .b(t_8162), .c(t_8159), .d(t_10602), .cin(t_10605), .o(t_10612), .co(t_10613), .cout(t_10614));
compressor_4_2 u2_3683(.a(t_8174), .b(t_8171), .c(t_8168), .d(t_10608), .cin(t_10611), .o(t_10615), .co(t_10616), .cout(t_10617));
compressor_4_2 u2_3684(.a(t_8142), .b(t_8139), .c(t_8136), .d(t_8180), .cin(t_8177), .o(t_10618), .co(t_10619), .cout(t_10620));
compressor_4_2 u2_3685(.a(t_8157), .b(t_8154), .c(t_8151), .d(t_8148), .cin(t_8145), .o(t_10621), .co(t_10622), .cout(t_10623));
compressor_4_2 u2_3686(.a(t_8186), .b(t_8183), .c(t_3464), .d(t_10614), .cin(t_10617), .o(t_10624), .co(t_10625), .cout(t_10626));
compressor_4_2 u2_3687(.a(t_8195), .b(t_8192), .c(t_8189), .d(t_10620), .cin(t_10623), .o(t_10627), .co(t_10628), .cout(t_10629));
compressor_4_2 u2_3688(.a(t_8163), .b(t_8160), .c(t_8204), .d(t_8201), .cin(t_8198), .o(t_10630), .co(t_10631), .cout(t_10632));
compressor_4_2 u2_3689(.a(t_8178), .b(t_8175), .c(t_8172), .d(t_8169), .cin(t_8166), .o(t_10633), .co(t_10634), .cout(t_10635));
compressor_4_2 u2_3690(.a(t_8209), .b(t_8206), .c(t_3511), .d(t_10626), .cin(t_10629), .o(t_10636), .co(t_10637), .cout(t_10638));
compressor_4_2 u2_3691(.a(t_8218), .b(t_8215), .c(t_8212), .d(t_10632), .cin(t_10635), .o(t_10639), .co(t_10640), .cout(t_10641));
compressor_4_2 u2_3692(.a(t_8187), .b(t_8184), .c(t_8227), .d(t_8224), .cin(t_8221), .o(t_10642), .co(t_10643), .cout(t_10644));
compressor_4_2 u2_3693(.a(t_8202), .b(t_8199), .c(t_8196), .d(t_8193), .cin(t_8190), .o(t_10645), .co(t_10646), .cout(t_10647));
compressor_4_2 u2_3694(.a(t_8232), .b(t_8229), .c(t_3558), .d(t_10638), .cin(t_10641), .o(t_10648), .co(t_10649), .cout(t_10650));
compressor_4_2 u2_3695(.a(t_8241), .b(t_8238), .c(t_8235), .d(t_10644), .cin(t_10647), .o(t_10651), .co(t_10652), .cout(t_10653));
compressor_4_2 u2_3696(.a(t_8210), .b(t_8207), .c(t_8250), .d(t_8247), .cin(t_8244), .o(t_10654), .co(t_10655), .cout(t_10656));
compressor_4_2 u2_3697(.a(t_8225), .b(t_8222), .c(t_8219), .d(t_8216), .cin(t_8213), .o(t_10657), .co(t_10658), .cout(t_10659));
compressor_4_2 u2_3698(.a(t_8255), .b(t_8252), .c(t_3605), .d(t_10650), .cin(t_10653), .o(t_10660), .co(t_10661), .cout(t_10662));
compressor_4_2 u2_3699(.a(t_8264), .b(t_8261), .c(t_8258), .d(t_10656), .cin(t_10659), .o(t_10663), .co(t_10664), .cout(t_10665));
compressor_4_2 u2_3700(.a(t_8233), .b(t_8230), .c(t_8273), .d(t_8270), .cin(t_8267), .o(t_10666), .co(t_10667), .cout(t_10668));
compressor_4_2 u2_3701(.a(t_8248), .b(t_8245), .c(t_8242), .d(t_8239), .cin(t_8236), .o(t_10669), .co(t_10670), .cout(t_10671));
compressor_4_2 u2_3702(.a(t_8278), .b(t_8275), .c(t_3652), .d(t_10662), .cin(t_10665), .o(t_10672), .co(t_10673), .cout(t_10674));
compressor_4_2 u2_3703(.a(t_8287), .b(t_8284), .c(t_8281), .d(t_10668), .cin(t_10671), .o(t_10675), .co(t_10676), .cout(t_10677));
compressor_4_2 u2_3704(.a(t_8256), .b(t_8253), .c(t_8296), .d(t_8293), .cin(t_8290), .o(t_10678), .co(t_10679), .cout(t_10680));
compressor_4_2 u2_3705(.a(t_8271), .b(t_8268), .c(t_8265), .d(t_8262), .cin(t_8259), .o(t_10681), .co(t_10682), .cout(t_10683));
compressor_4_2 u2_3706(.a(t_8304), .b(t_8301), .c(t_8298), .d(t_10674), .cin(t_10677), .o(t_10684), .co(t_10685), .cout(t_10686));
compressor_4_2 u2_3707(.a(t_8313), .b(t_8310), .c(t_8307), .d(t_10680), .cin(t_10683), .o(t_10687), .co(t_10688), .cout(t_10689));
compressor_4_2 u2_3708(.a(t_8282), .b(t_8279), .c(t_8276), .d(t_8319), .cin(t_8316), .o(t_10690), .co(t_10691), .cout(t_10692));
compressor_3_2 u1_3709(.a(t_8291), .b(t_8288), .cin(t_8285), .o(t_10693), .cout(t_10694));
compressor_4_2 u2_3710(.a(t_8324), .b(t_8321), .c(t_3744), .d(t_10686), .cin(t_10689), .o(t_10695), .co(t_10696), .cout(t_10697));
compressor_4_2 u2_3711(.a(t_8333), .b(t_8330), .c(t_8327), .d(t_10692), .cin(t_10694), .o(t_10698), .co(t_10699), .cout(t_10700));
compressor_4_2 u2_3712(.a(t_8302), .b(t_8299), .c(t_8342), .d(t_8339), .cin(t_8336), .o(t_10701), .co(t_10702), .cout(t_10703));
compressor_4_2 u2_3713(.a(t_8317), .b(t_8314), .c(t_8311), .d(t_8308), .cin(t_8305), .o(t_10704), .co(t_10705), .cout(t_10706));
compressor_4_2 u2_3714(.a(t_8350), .b(t_8347), .c(t_8344), .d(t_10697), .cin(t_10700), .o(t_10707), .co(t_10708), .cout(t_10709));
compressor_4_2 u2_3715(.a(t_8359), .b(t_8356), .c(t_8353), .d(t_10703), .cin(t_10706), .o(t_10710), .co(t_10711), .cout(t_10712));
compressor_4_2 u2_3716(.a(t_8328), .b(t_8325), .c(t_8322), .d(t_8365), .cin(t_8362), .o(t_10713), .co(t_10714), .cout(t_10715));
compressor_3_2 u1_3717(.a(t_8337), .b(t_8334), .cin(t_8331), .o(t_10716), .cout(t_10717));
compressor_4_2 u2_3718(.a(t_8373), .b(t_8370), .c(t_8367), .d(t_10709), .cin(t_10712), .o(t_10718), .co(t_10719), .cout(t_10720));
compressor_4_2 u2_3719(.a(t_8382), .b(t_8379), .c(t_8376), .d(t_10715), .cin(t_10717), .o(t_10721), .co(t_10722), .cout(t_10723));
compressor_4_2 u2_3720(.a(t_8351), .b(t_8348), .c(t_8345), .d(t_8388), .cin(t_8385), .o(t_10724), .co(t_10725), .cout(t_10726));
compressor_3_2 u1_3721(.a(t_8360), .b(t_8357), .cin(t_8354), .o(t_10727), .cout(t_10728));
compressor_4_2 u2_3722(.a(t_8396), .b(t_8393), .c(t_8390), .d(t_10720), .cin(t_10723), .o(t_10729), .co(t_10730), .cout(t_10731));
compressor_4_2 u2_3723(.a(t_8405), .b(t_8402), .c(t_8399), .d(t_10726), .cin(t_10728), .o(t_10732), .co(t_10733), .cout(t_10734));
compressor_4_2 u2_3724(.a(t_8374), .b(t_8371), .c(t_8368), .d(t_8411), .cin(t_8408), .o(t_10735), .co(t_10736), .cout(t_10737));
compressor_3_2 u1_3725(.a(t_8383), .b(t_8380), .cin(t_8377), .o(t_10738), .cout(t_10739));
compressor_4_2 u2_3726(.a(t_8419), .b(t_8416), .c(t_8413), .d(t_10731), .cin(t_10734), .o(t_10740), .co(t_10741), .cout(t_10742));
compressor_4_2 u2_3727(.a(t_8428), .b(t_8425), .c(t_8422), .d(t_10737), .cin(t_10739), .o(t_10743), .co(t_10744), .cout(t_10745));
compressor_4_2 u2_3728(.a(t_8397), .b(t_8394), .c(t_8391), .d(t_8434), .cin(t_8431), .o(t_10746), .co(t_10747), .cout(t_10748));
compressor_3_2 u1_3729(.a(t_8406), .b(t_8403), .cin(t_8400), .o(t_10749), .cout(t_10750));
compressor_4_2 u2_3730(.a(t_8442), .b(t_8439), .c(t_8436), .d(t_10742), .cin(t_10745), .o(t_10751), .co(t_10752), .cout(t_10753));
compressor_4_2 u2_3731(.a(t_8451), .b(t_8448), .c(t_8445), .d(t_10748), .cin(t_10750), .o(t_10754), .co(t_10755), .cout(t_10756));
compressor_4_2 u2_3732(.a(t_8420), .b(t_8417), .c(t_8414), .d(t_8457), .cin(t_8454), .o(t_10757), .co(t_10758), .cout(t_10759));
compressor_3_2 u1_3733(.a(t_8429), .b(t_8426), .cin(t_8423), .o(t_10760), .cout(t_10761));
compressor_4_2 u2_3734(.a(t_8465), .b(t_8462), .c(t_8459), .d(t_10753), .cin(t_10756), .o(t_10762), .co(t_10763), .cout(t_10764));
compressor_4_2 u2_3735(.a(t_8474), .b(t_8471), .c(t_8468), .d(t_10759), .cin(t_10761), .o(t_10765), .co(t_10766), .cout(t_10767));
compressor_4_2 u2_3736(.a(t_8443), .b(t_8440), .c(t_8437), .d(t_8480), .cin(t_8477), .o(t_10768), .co(t_10769), .cout(t_10770));
compressor_3_2 u1_3737(.a(t_8452), .b(t_8449), .cin(t_8446), .o(t_10771), .cout(t_10772));
compressor_4_2 u2_3738(.a(t_8485), .b(t_8482), .c(t_4050), .d(t_10764), .cin(t_10767), .o(t_10773), .co(t_10774), .cout(t_10775));
compressor_4_2 u2_3739(.a(t_8494), .b(t_8491), .c(t_8488), .d(t_10770), .cin(t_10772), .o(t_10776), .co(t_10777), .cout(t_10778));
compressor_4_2 u2_3740(.a(t_8466), .b(t_8463), .c(t_8460), .d(t_8500), .cin(t_8497), .o(t_10779), .co(t_10780), .cout(t_10781));
compressor_3_2 u1_3741(.a(t_8475), .b(t_8472), .cin(t_8469), .o(t_10782), .cout(t_10783));
compressor_4_2 u2_3742(.a(t_8506), .b(t_8503), .c(t_4092), .d(t_10775), .cin(t_10778), .o(t_10784), .co(t_10785), .cout(t_10786));
compressor_4_2 u2_3743(.a(t_8515), .b(t_8512), .c(t_8509), .d(t_10781), .cin(t_10783), .o(t_10787), .co(t_10788), .cout(t_10789));
compressor_4_2 u2_3744(.a(t_8489), .b(t_8486), .c(t_8483), .d(t_8521), .cin(t_8518), .o(t_10790), .co(t_10791), .cout(t_10792));
compressor_3_2 u1_3745(.a(t_8498), .b(t_8495), .cin(t_8492), .o(t_10793), .cout(t_10794));
compressor_4_2 u2_3746(.a(t_8530), .b(t_8527), .c(t_8524), .d(t_10786), .cin(t_10789), .o(t_10795), .co(t_10796), .cout(t_10797));
compressor_4_2 u2_3747(.a(t_8539), .b(t_8536), .c(t_8533), .d(t_10792), .cin(t_10794), .o(t_10798), .co(t_10799), .cout(t_10800));
compressor_4_2 u2_3748(.a(t_8513), .b(t_8510), .c(t_8507), .d(t_8504), .cin(t_8542), .o(t_10801), .co(t_10802), .cout(t_10803));
compressor_3_2 u1_3749(.a(t_8522), .b(t_8519), .cin(t_8516), .o(t_10804), .cout(t_10805));
compressor_4_2 u2_3750(.a(t_8548), .b(t_8545), .c(t_4172), .d(t_10797), .cin(t_10800), .o(t_10806), .co(t_10807), .cout(t_10808));
compressor_4_2 u2_3751(.a(t_8557), .b(t_8554), .c(t_8551), .d(t_10803), .cin(t_10805), .o(t_10809), .co(t_10810), .cout(t_10811));
compressor_4_2 u2_3752(.a(t_8531), .b(t_8528), .c(t_8525), .d(t_8563), .cin(t_8560), .o(t_10812), .co(t_10813), .cout(t_10814));
compressor_3_2 u1_3753(.a(t_8540), .b(t_8537), .cin(t_8534), .o(t_10815), .cout(t_10816));
compressor_4_2 u2_3754(.a(t_8568), .b(t_8565), .c(t_4213), .d(t_10808), .cin(t_10811), .o(t_10817), .co(t_10818), .cout(t_10819));
compressor_4_2 u2_3755(.a(t_8577), .b(t_8574), .c(t_8571), .d(t_10814), .cin(t_10816), .o(t_10820), .co(t_10821), .cout(t_10822));
compressor_4_2 u2_3756(.a(t_8552), .b(t_8549), .c(t_8546), .d(t_8583), .cin(t_8580), .o(t_10823), .co(t_10824), .cout(t_10825));
compressor_3_2 u1_3757(.a(t_8561), .b(t_8558), .cin(t_8555), .o(t_10826), .cout(t_10827));
compressor_4_2 u2_3758(.a(t_8588), .b(t_8585), .c(t_4254), .d(t_10819), .cin(t_10822), .o(t_10828), .co(t_10829), .cout(t_10830));
compressor_4_2 u2_3759(.a(t_8597), .b(t_8594), .c(t_8591), .d(t_10825), .cin(t_10827), .o(t_10831), .co(t_10832), .cout(t_10833));
compressor_4_2 u2_3760(.a(t_8572), .b(t_8569), .c(t_8566), .d(t_8603), .cin(t_8600), .o(t_10834), .co(t_10835), .cout(t_10836));
compressor_3_2 u1_3761(.a(t_8581), .b(t_8578), .cin(t_8575), .o(t_10837), .cout(t_10838));
compressor_4_2 u2_3762(.a(t_8608), .b(t_8605), .c(t_4295), .d(t_10830), .cin(t_10833), .o(t_10839), .co(t_10840), .cout(t_10841));
compressor_4_2 u2_3763(.a(t_8617), .b(t_8614), .c(t_8611), .d(t_10836), .cin(t_10838), .o(t_10842), .co(t_10843), .cout(t_10844));
compressor_4_2 u2_3764(.a(t_8592), .b(t_8589), .c(t_8586), .d(t_8623), .cin(t_8620), .o(t_10845), .co(t_10846), .cout(t_10847));
compressor_3_2 u1_3765(.a(t_8601), .b(t_8598), .cin(t_8595), .o(t_10848), .cout(t_10849));
compressor_4_2 u2_3766(.a(t_8628), .b(t_8625), .c(t_4336), .d(t_10841), .cin(t_10844), .o(t_10850), .co(t_10851), .cout(t_10852));
compressor_4_2 u2_3767(.a(t_8637), .b(t_8634), .c(t_8631), .d(t_10847), .cin(t_10849), .o(t_10853), .co(t_10854), .cout(t_10855));
compressor_4_2 u2_3768(.a(t_8612), .b(t_8609), .c(t_8606), .d(t_8643), .cin(t_8640), .o(t_10856), .co(t_10857), .cout(t_10858));
compressor_3_2 u1_3769(.a(t_8621), .b(t_8618), .cin(t_8615), .o(t_10859), .cout(t_10860));
compressor_4_2 u2_3770(.a(t_8651), .b(t_8648), .c(t_8645), .d(t_10852), .cin(t_10855), .o(t_10861), .co(t_10862), .cout(t_10863));
compressor_4_2 u2_3771(.a(t_8660), .b(t_8657), .c(t_8654), .d(t_10858), .cin(t_10860), .o(t_10864), .co(t_10865), .cout(t_10866));
compressor_4_2 u2_3772(.a(t_8635), .b(t_8632), .c(t_8629), .d(t_8626), .cin(t_8663), .o(t_10867), .co(t_10868), .cout(t_10869));
half_adder u0_3773(.a(t_8641), .b(t_8638), .o(t_10870), .cout(t_10871));
compressor_4_2 u2_3774(.a(t_8668), .b(t_8665), .c(t_4416), .d(t_10863), .cin(t_10866), .o(t_10872), .co(t_10873), .cout(t_10874));
compressor_4_2 u2_3775(.a(t_8677), .b(t_8674), .c(t_8671), .d(t_10869), .cin(t_10871), .o(t_10875), .co(t_10876), .cout(t_10877));
compressor_4_2 u2_3776(.a(t_8652), .b(t_8649), .c(t_8646), .d(t_8683), .cin(t_8680), .o(t_10878), .co(t_10879), .cout(t_10880));
compressor_3_2 u1_3777(.a(t_8661), .b(t_8658), .cin(t_8655), .o(t_10881), .cout(t_10882));
compressor_4_2 u2_3778(.a(t_8691), .b(t_8688), .c(t_8685), .d(t_10874), .cin(t_10877), .o(t_10883), .co(t_10884), .cout(t_10885));
compressor_4_2 u2_3779(.a(t_8700), .b(t_8697), .c(t_8694), .d(t_10880), .cin(t_10882), .o(t_10886), .co(t_10887), .cout(t_10888));
compressor_4_2 u2_3780(.a(t_8675), .b(t_8672), .c(t_8669), .d(t_8666), .cin(t_8703), .o(t_10889), .co(t_10890), .cout(t_10891));
half_adder u0_3781(.a(t_8681), .b(t_8678), .o(t_10892), .cout(t_10893));
compressor_4_2 u2_3782(.a(t_8711), .b(t_8708), .c(t_8705), .d(t_10885), .cin(t_10888), .o(t_10894), .co(t_10895), .cout(t_10896));
compressor_4_2 u2_3783(.a(t_8720), .b(t_8717), .c(t_8714), .d(t_10891), .cin(t_10893), .o(t_10897), .co(t_10898), .cout(t_10899));
compressor_4_2 u2_3784(.a(t_8695), .b(t_8692), .c(t_8689), .d(t_8686), .cin(t_8723), .o(t_10900), .co(t_10901), .cout(t_10902));
half_adder u0_3785(.a(t_8701), .b(t_8698), .o(t_10903), .cout(t_10904));
compressor_4_2 u2_3786(.a(t_8731), .b(t_8728), .c(t_8725), .d(t_10896), .cin(t_10899), .o(t_10905), .co(t_10906), .cout(t_10907));
compressor_4_2 u2_3787(.a(t_8740), .b(t_8737), .c(t_8734), .d(t_10902), .cin(t_10904), .o(t_10908), .co(t_10909), .cout(t_10910));
compressor_4_2 u2_3788(.a(t_8715), .b(t_8712), .c(t_8709), .d(t_8706), .cin(t_8743), .o(t_10911), .co(t_10912), .cout(t_10913));
half_adder u0_3789(.a(t_8721), .b(t_8718), .o(t_10914), .cout(t_10915));
compressor_4_2 u2_3790(.a(t_8751), .b(t_8748), .c(t_8745), .d(t_10907), .cin(t_10910), .o(t_10916), .co(t_10917), .cout(t_10918));
compressor_4_2 u2_3791(.a(t_8760), .b(t_8757), .c(t_8754), .d(t_10913), .cin(t_10915), .o(t_10919), .co(t_10920), .cout(t_10921));
compressor_4_2 u2_3792(.a(t_8735), .b(t_8732), .c(t_8729), .d(t_8726), .cin(t_8763), .o(t_10922), .co(t_10923), .cout(t_10924));
half_adder u0_3793(.a(t_8741), .b(t_8738), .o(t_10925), .cout(t_10926));
compressor_4_2 u2_3794(.a(t_8771), .b(t_8768), .c(t_8765), .d(t_10918), .cin(t_10921), .o(t_10927), .co(t_10928), .cout(t_10929));
compressor_4_2 u2_3795(.a(t_8780), .b(t_8777), .c(t_8774), .d(t_10924), .cin(t_10926), .o(t_10930), .co(t_10931), .cout(t_10932));
compressor_4_2 u2_3796(.a(t_8755), .b(t_8752), .c(t_8749), .d(t_8746), .cin(t_8783), .o(t_10933), .co(t_10934), .cout(t_10935));
half_adder u0_3797(.a(t_8761), .b(t_8758), .o(t_10936), .cout(t_10937));
compressor_4_2 u2_3798(.a(t_8791), .b(t_8788), .c(t_8785), .d(t_10929), .cin(t_10932), .o(t_10938), .co(t_10939), .cout(t_10940));
compressor_4_2 u2_3799(.a(t_8800), .b(t_8797), .c(t_8794), .d(t_10935), .cin(t_10937), .o(t_10941), .co(t_10942), .cout(t_10943));
compressor_4_2 u2_3800(.a(t_8775), .b(t_8772), .c(t_8769), .d(t_8766), .cin(t_8803), .o(t_10944), .co(t_10945), .cout(t_10946));
half_adder u0_3801(.a(t_8781), .b(t_8778), .o(t_10947), .cout(t_10948));
compressor_4_2 u2_3802(.a(t_8808), .b(t_8805), .c(t_4680), .d(t_10940), .cin(t_10943), .o(t_10949), .co(t_10950), .cout(t_10951));
compressor_4_2 u2_3803(.a(t_8817), .b(t_8814), .c(t_8811), .d(t_10946), .cin(t_10948), .o(t_10952), .co(t_10953), .cout(t_10954));
compressor_4_2 u2_3804(.a(t_8795), .b(t_8792), .c(t_8789), .d(t_8786), .cin(t_8820), .o(t_10955), .co(t_10956), .cout(t_10957));
half_adder u0_3805(.a(t_8801), .b(t_8798), .o(t_10958), .cout(t_10959));
compressor_4_2 u2_3806(.a(t_8826), .b(t_8823), .c(t_4716), .d(t_10951), .cin(t_10954), .o(t_10960), .co(t_10961), .cout(t_10962));
compressor_4_2 u2_3807(.a(t_8835), .b(t_8832), .c(t_8829), .d(t_10957), .cin(t_10959), .o(t_10963), .co(t_10964), .cout(t_10965));
compressor_4_2 u2_3808(.a(t_8815), .b(t_8812), .c(t_8809), .d(t_8806), .cin(t_8838), .o(t_10966), .co(t_10967), .cout(t_10968));
half_adder u0_3809(.a(t_8821), .b(t_8818), .o(t_10969), .cout(t_10970));
compressor_4_2 u2_3810(.a(t_8847), .b(t_8844), .c(t_8841), .d(t_10962), .cin(t_10965), .o(t_10971), .co(t_10972), .cout(t_10973));
compressor_4_2 u2_3811(.a(t_8856), .b(t_8853), .c(t_8850), .d(t_10968), .cin(t_10970), .o(t_10974), .co(t_10975), .cout(t_10976));
compressor_4_2 u2_3812(.a(t_8836), .b(t_8833), .c(t_8830), .d(t_8827), .cin(t_8824), .o(t_10977), .co(t_10978), .cout(t_10979));
compressor_4_2 u2_3813(.a(t_8862), .b(t_8859), .c(t_4784), .d(t_10973), .cin(t_10976), .o(t_10980), .co(t_10981), .cout(t_10982));
compressor_4_2 u2_3814(.a(t_8874), .b(t_8871), .c(t_8868), .d(t_8865), .cin(t_10979), .o(t_10983), .co(t_10984), .cout(t_10985));
compressor_4_2 u2_3815(.a(t_8854), .b(t_8851), .c(t_8848), .d(t_8845), .cin(t_8842), .o(t_10986), .co(t_10987), .cout(t_10988));
compressor_4_2 u2_3816(.a(t_8879), .b(t_8876), .c(t_4819), .d(t_10982), .cin(t_10985), .o(t_10989), .co(t_10990), .cout(t_10991));
compressor_4_2 u2_3817(.a(t_8891), .b(t_8888), .c(t_8885), .d(t_8882), .cin(t_10988), .o(t_10992), .co(t_10993), .cout(t_10994));
compressor_4_2 u2_3818(.a(t_8872), .b(t_8869), .c(t_8866), .d(t_8863), .cin(t_8860), .o(t_10995), .co(t_10996), .cout(t_10997));
compressor_4_2 u2_3819(.a(t_8896), .b(t_8893), .c(t_4854), .d(t_10991), .cin(t_10994), .o(t_10998), .co(t_10999), .cout(t_11000));
compressor_4_2 u2_3820(.a(t_8908), .b(t_8905), .c(t_8902), .d(t_8899), .cin(t_10997), .o(t_11001), .co(t_11002), .cout(t_11003));
compressor_4_2 u2_3821(.a(t_8889), .b(t_8886), .c(t_8883), .d(t_8880), .cin(t_8877), .o(t_11004), .co(t_11005), .cout(t_11006));
compressor_4_2 u2_3822(.a(t_8913), .b(t_8910), .c(t_4889), .d(t_11000), .cin(t_11003), .o(t_11007), .co(t_11008), .cout(t_11009));
compressor_4_2 u2_3823(.a(t_8925), .b(t_8922), .c(t_8919), .d(t_8916), .cin(t_11006), .o(t_11010), .co(t_11011), .cout(t_11012));
compressor_4_2 u2_3824(.a(t_8906), .b(t_8903), .c(t_8900), .d(t_8897), .cin(t_8894), .o(t_11013), .co(t_11014), .cout(t_11015));
compressor_4_2 u2_3825(.a(t_8930), .b(t_8927), .c(t_4924), .d(t_11009), .cin(t_11012), .o(t_11016), .co(t_11017), .cout(t_11018));
compressor_4_2 u2_3826(.a(t_8942), .b(t_8939), .c(t_8936), .d(t_8933), .cin(t_11015), .o(t_11019), .co(t_11020), .cout(t_11021));
compressor_4_2 u2_3827(.a(t_8923), .b(t_8920), .c(t_8917), .d(t_8914), .cin(t_8911), .o(t_11022), .co(t_11023), .cout(t_11024));
compressor_4_2 u2_3828(.a(t_8950), .b(t_8947), .c(t_8944), .d(t_11018), .cin(t_11021), .o(t_11025), .co(t_11026), .cout(t_11027));
compressor_4_2 u2_3829(.a(t_8928), .b(t_8959), .c(t_8956), .d(t_8953), .cin(t_11024), .o(t_11028), .co(t_11029), .cout(t_11030));
compressor_3_2 u1_3830(.a(t_8937), .b(t_8934), .cin(t_8931), .o(t_11031), .cout(t_11032));
compressor_4_2 u2_3831(.a(t_8964), .b(t_8961), .c(t_4992), .d(t_11027), .cin(t_11030), .o(t_11033), .co(t_11034), .cout(t_11035));
compressor_4_2 u2_3832(.a(t_8976), .b(t_8973), .c(t_8970), .d(t_8967), .cin(t_11032), .o(t_11036), .co(t_11037), .cout(t_11038));
compressor_4_2 u2_3833(.a(t_8957), .b(t_8954), .c(t_8951), .d(t_8948), .cin(t_8945), .o(t_11039), .co(t_11040), .cout(t_11041));
compressor_4_2 u2_3834(.a(t_8984), .b(t_8981), .c(t_8978), .d(t_11035), .cin(t_11038), .o(t_11042), .co(t_11043), .cout(t_11044));
compressor_4_2 u2_3835(.a(t_8962), .b(t_8993), .c(t_8990), .d(t_8987), .cin(t_11041), .o(t_11045), .co(t_11046), .cout(t_11047));
compressor_3_2 u1_3836(.a(t_8971), .b(t_8968), .cin(t_8965), .o(t_11048), .cout(t_11049));
compressor_4_2 u2_3837(.a(t_9001), .b(t_8998), .c(t_8995), .d(t_11044), .cin(t_11047), .o(t_11050), .co(t_11051), .cout(t_11052));
compressor_4_2 u2_3838(.a(t_8979), .b(t_9010), .c(t_9007), .d(t_9004), .cin(t_11049), .o(t_11053), .co(t_11054), .cout(t_11055));
compressor_3_2 u1_3839(.a(t_8988), .b(t_8985), .cin(t_8982), .o(t_11056), .cout(t_11057));
compressor_4_2 u2_3840(.a(t_9018), .b(t_9015), .c(t_9012), .d(t_11052), .cin(t_11055), .o(t_11058), .co(t_11059), .cout(t_11060));
compressor_4_2 u2_3841(.a(t_8996), .b(t_9027), .c(t_9024), .d(t_9021), .cin(t_11057), .o(t_11061), .co(t_11062), .cout(t_11063));
compressor_3_2 u1_3842(.a(t_9005), .b(t_9002), .cin(t_8999), .o(t_11064), .cout(t_11065));
compressor_4_2 u2_3843(.a(t_9035), .b(t_9032), .c(t_9029), .d(t_11060), .cin(t_11063), .o(t_11066), .co(t_11067), .cout(t_11068));
compressor_4_2 u2_3844(.a(t_9013), .b(t_9044), .c(t_9041), .d(t_9038), .cin(t_11065), .o(t_11069), .co(t_11070), .cout(t_11071));
compressor_3_2 u1_3845(.a(t_9022), .b(t_9019), .cin(t_9016), .o(t_11072), .cout(t_11073));
compressor_4_2 u2_3846(.a(t_9052), .b(t_9049), .c(t_9046), .d(t_11068), .cin(t_11071), .o(t_11074), .co(t_11075), .cout(t_11076));
compressor_4_2 u2_3847(.a(t_9030), .b(t_9061), .c(t_9058), .d(t_9055), .cin(t_11073), .o(t_11077), .co(t_11078), .cout(t_11079));
compressor_3_2 u1_3848(.a(t_9039), .b(t_9036), .cin(t_9033), .o(t_11080), .cout(t_11081));
compressor_4_2 u2_3849(.a(t_9069), .b(t_9066), .c(t_9063), .d(t_11076), .cin(t_11079), .o(t_11082), .co(t_11083), .cout(t_11084));
compressor_4_2 u2_3850(.a(t_9047), .b(t_9078), .c(t_9075), .d(t_9072), .cin(t_11081), .o(t_11085), .co(t_11086), .cout(t_11087));
compressor_3_2 u1_3851(.a(t_9056), .b(t_9053), .cin(t_9050), .o(t_11088), .cout(t_11089));
compressor_4_2 u2_3852(.a(t_9083), .b(t_9080), .c(t_5214), .d(t_11084), .cin(t_11087), .o(t_11090), .co(t_11091), .cout(t_11092));
compressor_4_2 u2_3853(.a(t_9064), .b(t_9092), .c(t_9089), .d(t_9086), .cin(t_11089), .o(t_11093), .co(t_11094), .cout(t_11095));
compressor_3_2 u1_3854(.a(t_9073), .b(t_9070), .cin(t_9067), .o(t_11096), .cout(t_11097));
compressor_4_2 u2_3855(.a(t_9098), .b(t_9095), .c(t_5244), .d(t_11092), .cin(t_11095), .o(t_11098), .co(t_11099), .cout(t_11100));
compressor_4_2 u2_3856(.a(t_9081), .b(t_9107), .c(t_9104), .d(t_9101), .cin(t_11097), .o(t_11101), .co(t_11102), .cout(t_11103));
compressor_3_2 u1_3857(.a(t_9090), .b(t_9087), .cin(t_9084), .o(t_11104), .cout(t_11105));
compressor_4_2 u2_3858(.a(t_9116), .b(t_9113), .c(t_9110), .d(t_11100), .cin(t_11103), .o(t_11106), .co(t_11107), .cout(t_11108));
compressor_4_2 u2_3859(.a(t_9099), .b(t_9096), .c(t_9122), .d(t_9119), .cin(t_11105), .o(t_11109), .co(t_11110), .cout(t_11111));
compressor_3_2 u1_3860(.a(t_9108), .b(t_9105), .cin(t_9102), .o(t_11112), .cout(t_11113));
compressor_4_2 u2_3861(.a(t_9128), .b(t_9125), .c(t_5300), .d(t_11108), .cin(t_11111), .o(t_11114), .co(t_11115), .cout(t_11116));
compressor_4_2 u2_3862(.a(t_9111), .b(t_9137), .c(t_9134), .d(t_9131), .cin(t_11113), .o(t_11117), .co(t_11118), .cout(t_11119));
compressor_3_2 u1_3863(.a(t_9120), .b(t_9117), .cin(t_9114), .o(t_11120), .cout(t_11121));
compressor_4_2 u2_3864(.a(t_9142), .b(t_9139), .c(t_5329), .d(t_11116), .cin(t_11119), .o(t_11122), .co(t_11123), .cout(t_11124));
compressor_4_2 u2_3865(.a(t_9126), .b(t_9151), .c(t_9148), .d(t_9145), .cin(t_11121), .o(t_11125), .co(t_11126), .cout(t_11127));
compressor_3_2 u1_3866(.a(t_9135), .b(t_9132), .cin(t_9129), .o(t_11128), .cout(t_11129));
compressor_4_2 u2_3867(.a(t_9156), .b(t_9153), .c(t_5358), .d(t_11124), .cin(t_11127), .o(t_11130), .co(t_11131), .cout(t_11132));
compressor_4_2 u2_3868(.a(t_9140), .b(t_9165), .c(t_9162), .d(t_9159), .cin(t_11129), .o(t_11133), .co(t_11134), .cout(t_11135));
compressor_3_2 u1_3869(.a(t_9149), .b(t_9146), .cin(t_9143), .o(t_11136), .cout(t_11137));
compressor_4_2 u2_3870(.a(t_9170), .b(t_9167), .c(t_5387), .d(t_11132), .cin(t_11135), .o(t_11138), .co(t_11139), .cout(t_11140));
compressor_4_2 u2_3871(.a(t_9154), .b(t_9179), .c(t_9176), .d(t_9173), .cin(t_11137), .o(t_11141), .co(t_11142), .cout(t_11143));
compressor_3_2 u1_3872(.a(t_9163), .b(t_9160), .cin(t_9157), .o(t_11144), .cout(t_11145));
compressor_4_2 u2_3873(.a(t_9184), .b(t_9181), .c(t_5416), .d(t_11140), .cin(t_11143), .o(t_11146), .co(t_11147), .cout(t_11148));
compressor_4_2 u2_3874(.a(t_9168), .b(t_9193), .c(t_9190), .d(t_9187), .cin(t_11145), .o(t_11149), .co(t_11150), .cout(t_11151));
compressor_3_2 u1_3875(.a(t_9177), .b(t_9174), .cin(t_9171), .o(t_11152), .cout(t_11153));
compressor_4_2 u2_3876(.a(t_9201), .b(t_9198), .c(t_9195), .d(t_11148), .cin(t_11151), .o(t_11154), .co(t_11155), .cout(t_11156));
compressor_4_2 u2_3877(.a(t_9185), .b(t_9182), .c(t_9207), .d(t_9204), .cin(t_11153), .o(t_11157), .co(t_11158), .cout(t_11159));
half_adder u0_3878(.a(t_9191), .b(t_9188), .o(t_11160), .cout(t_11161));
compressor_4_2 u2_3879(.a(t_9212), .b(t_9209), .c(t_5472), .d(t_11156), .cin(t_11159), .o(t_11162), .co(t_11163), .cout(t_11164));
compressor_4_2 u2_3880(.a(t_9196), .b(t_9221), .c(t_9218), .d(t_9215), .cin(t_11161), .o(t_11165), .co(t_11166), .cout(t_11167));
compressor_3_2 u1_3881(.a(t_9205), .b(t_9202), .cin(t_9199), .o(t_11168), .cout(t_11169));
compressor_4_2 u2_3882(.a(t_9229), .b(t_9226), .c(t_9223), .d(t_11164), .cin(t_11167), .o(t_11170), .co(t_11171), .cout(t_11172));
compressor_4_2 u2_3883(.a(t_9213), .b(t_9210), .c(t_9235), .d(t_9232), .cin(t_11169), .o(t_11173), .co(t_11174), .cout(t_11175));
half_adder u0_3884(.a(t_9219), .b(t_9216), .o(t_11176), .cout(t_11177));
compressor_4_2 u2_3885(.a(t_9243), .b(t_9240), .c(t_9237), .d(t_11172), .cin(t_11175), .o(t_11178), .co(t_11179), .cout(t_11180));
compressor_4_2 u2_3886(.a(t_9227), .b(t_9224), .c(t_9249), .d(t_9246), .cin(t_11177), .o(t_11181), .co(t_11182), .cout(t_11183));
half_adder u0_3887(.a(t_9233), .b(t_9230), .o(t_11184), .cout(t_11185));
compressor_4_2 u2_3888(.a(t_9257), .b(t_9254), .c(t_9251), .d(t_11180), .cin(t_11183), .o(t_11186), .co(t_11187), .cout(t_11188));
compressor_4_2 u2_3889(.a(t_9241), .b(t_9238), .c(t_9263), .d(t_9260), .cin(t_11185), .o(t_11189), .co(t_11190), .cout(t_11191));
half_adder u0_3890(.a(t_9247), .b(t_9244), .o(t_11192), .cout(t_11193));
compressor_4_2 u2_3891(.a(t_9271), .b(t_9268), .c(t_9265), .d(t_11188), .cin(t_11191), .o(t_11194), .co(t_11195), .cout(t_11196));
compressor_4_2 u2_3892(.a(t_9255), .b(t_9252), .c(t_9277), .d(t_9274), .cin(t_11193), .o(t_11197), .co(t_11198), .cout(t_11199));
half_adder u0_3893(.a(t_9261), .b(t_9258), .o(t_11200), .cout(t_11201));
compressor_4_2 u2_3894(.a(t_9285), .b(t_9282), .c(t_9279), .d(t_11196), .cin(t_11199), .o(t_11202), .co(t_11203), .cout(t_11204));
compressor_4_2 u2_3895(.a(t_9269), .b(t_9266), .c(t_9291), .d(t_9288), .cin(t_11201), .o(t_11205), .co(t_11206), .cout(t_11207));
half_adder u0_3896(.a(t_9275), .b(t_9272), .o(t_11208), .cout(t_11209));
compressor_4_2 u2_3897(.a(t_9299), .b(t_9296), .c(t_9293), .d(t_11204), .cin(t_11207), .o(t_11210), .co(t_11211), .cout(t_11212));
compressor_4_2 u2_3898(.a(t_9283), .b(t_9280), .c(t_9305), .d(t_9302), .cin(t_11209), .o(t_11213), .co(t_11214), .cout(t_11215));
half_adder u0_3899(.a(t_9289), .b(t_9286), .o(t_11216), .cout(t_11217));
compressor_4_2 u2_3900(.a(t_9310), .b(t_9307), .c(t_5652), .d(t_11212), .cin(t_11215), .o(t_11218), .co(t_11219), .cout(t_11220));
compressor_4_2 u2_3901(.a(t_9297), .b(t_9294), .c(t_9316), .d(t_9313), .cin(t_11217), .o(t_11221), .co(t_11222), .cout(t_11223));
half_adder u0_3902(.a(t_9303), .b(t_9300), .o(t_11224), .cout(t_11225));
compressor_4_2 u2_3903(.a(t_9322), .b(t_9319), .c(t_5676), .d(t_11220), .cin(t_11223), .o(t_11226), .co(t_11227), .cout(t_11228));
compressor_4_2 u2_3904(.a(t_9311), .b(t_9308), .c(t_9328), .d(t_9325), .cin(t_11225), .o(t_11229), .co(t_11230), .cout(t_11231));
half_adder u0_3905(.a(t_9317), .b(t_9314), .o(t_11232), .cout(t_11233));
compressor_4_2 u2_3906(.a(t_9337), .b(t_9334), .c(t_9331), .d(t_11228), .cin(t_11231), .o(t_11234), .co(t_11235), .cout(t_11236));
compressor_4_2 u2_3907(.a(t_9326), .b(t_9323), .c(t_9320), .d(t_9340), .cin(t_11233), .o(t_11237), .co(t_11238), .cout(t_11239));
compressor_4_2 u2_3908(.a(t_9346), .b(t_9343), .c(t_5720), .d(t_11236), .cin(t_11239), .o(t_11240), .co(t_11241), .cout(t_11242));
compressor_4_2 u2_3909(.a(t_9338), .b(t_9335), .c(t_9332), .d(t_9352), .cin(t_9349), .o(t_11243), .co(t_11244), .cout(t_11245));
compressor_4_2 u2_3910(.a(t_9357), .b(t_9354), .c(t_5743), .d(t_11242), .cin(t_11245), .o(t_11246), .co(t_11247), .cout(t_11248));
compressor_4_2 u2_3911(.a(t_9350), .b(t_9347), .c(t_9344), .d(t_9363), .cin(t_9360), .o(t_11249), .co(t_11250), .cout(t_11251));
compressor_4_2 u2_3912(.a(t_9368), .b(t_9365), .c(t_5766), .d(t_11248), .cin(t_11251), .o(t_11252), .co(t_11253), .cout(t_11254));
compressor_4_2 u2_3913(.a(t_9361), .b(t_9358), .c(t_9355), .d(t_9374), .cin(t_9371), .o(t_11255), .co(t_11256), .cout(t_11257));
compressor_4_2 u2_3914(.a(t_9379), .b(t_9376), .c(t_5789), .d(t_11254), .cin(t_11257), .o(t_11258), .co(t_11259), .cout(t_11260));
compressor_4_2 u2_3915(.a(t_9372), .b(t_9369), .c(t_9366), .d(t_9385), .cin(t_9382), .o(t_11261), .co(t_11262), .cout(t_11263));
compressor_4_2 u2_3916(.a(t_9390), .b(t_9387), .c(t_5812), .d(t_11260), .cin(t_11263), .o(t_11264), .co(t_11265), .cout(t_11266));
compressor_4_2 u2_3917(.a(t_9383), .b(t_9380), .c(t_9377), .d(t_9396), .cin(t_9393), .o(t_11267), .co(t_11268), .cout(t_11269));
compressor_4_2 u2_3918(.a(t_9404), .b(t_9401), .c(t_9398), .d(t_11266), .cin(t_11269), .o(t_11270), .co(t_11271), .cout(t_11272));
compressor_3_2 u1_3919(.a(t_9391), .b(t_9388), .cin(t_9407), .o(t_11273), .cout(t_11274));
compressor_4_2 u2_3920(.a(t_9412), .b(t_9409), .c(t_5856), .d(t_11272), .cin(t_11274), .o(t_11275), .co(t_11276), .cout(t_11277));
compressor_4_2 u2_3921(.a(t_9405), .b(t_9402), .c(t_9399), .d(t_9418), .cin(t_9415), .o(t_11278), .co(t_11279), .cout(t_11280));
compressor_4_2 u2_3922(.a(t_9426), .b(t_9423), .c(t_9420), .d(t_11277), .cin(t_11280), .o(t_11281), .co(t_11282), .cout(t_11283));
compressor_3_2 u1_3923(.a(t_9413), .b(t_9410), .cin(t_9429), .o(t_11284), .cout(t_11285));
compressor_4_2 u2_3924(.a(t_9437), .b(t_9434), .c(t_9431), .d(t_11283), .cin(t_11285), .o(t_11286), .co(t_11287), .cout(t_11288));
compressor_3_2 u1_3925(.a(t_9424), .b(t_9421), .cin(t_9440), .o(t_11289), .cout(t_11290));
compressor_4_2 u2_3926(.a(t_9448), .b(t_9445), .c(t_9442), .d(t_11288), .cin(t_11290), .o(t_11291), .co(t_11292), .cout(t_11293));
compressor_3_2 u1_3927(.a(t_9435), .b(t_9432), .cin(t_9451), .o(t_11294), .cout(t_11295));
compressor_4_2 u2_3928(.a(t_9459), .b(t_9456), .c(t_9453), .d(t_11293), .cin(t_11295), .o(t_11296), .co(t_11297), .cout(t_11298));
compressor_3_2 u1_3929(.a(t_9446), .b(t_9443), .cin(t_9462), .o(t_11299), .cout(t_11300));
compressor_4_2 u2_3930(.a(t_9470), .b(t_9467), .c(t_9464), .d(t_11298), .cin(t_11300), .o(t_11301), .co(t_11302), .cout(t_11303));
compressor_3_2 u1_3931(.a(t_9457), .b(t_9454), .cin(t_9473), .o(t_11304), .cout(t_11305));
compressor_4_2 u2_3932(.a(t_9481), .b(t_9478), .c(t_9475), .d(t_11303), .cin(t_11305), .o(t_11306), .co(t_11307), .cout(t_11308));
compressor_3_2 u1_3933(.a(t_9468), .b(t_9465), .cin(t_9484), .o(t_11309), .cout(t_11310));
compressor_4_2 u2_3934(.a(t_9489), .b(t_9486), .c(t_5994), .d(t_11308), .cin(t_11310), .o(t_11311), .co(t_11312), .cout(t_11313));
compressor_3_2 u1_3935(.a(t_9479), .b(t_9476), .cin(t_9492), .o(t_11314), .cout(t_11315));
compressor_4_2 u2_3936(.a(t_9498), .b(t_9495), .c(t_6012), .d(t_11313), .cin(t_11315), .o(t_11316), .co(t_11317), .cout(t_11318));
compressor_3_2 u1_3937(.a(t_9490), .b(t_9487), .cin(t_9501), .o(t_11319), .cout(t_11320));
compressor_4_2 u2_3938(.a(t_9510), .b(t_9507), .c(t_9504), .d(t_11318), .cin(t_11320), .o(t_11321), .co(t_11322), .cout(t_11323));
compressor_3_2 u1_3939(.a(t_9502), .b(t_9499), .cin(t_9496), .o(t_11324), .cout(t_11325));
compressor_4_2 u2_3940(.a(t_9516), .b(t_9513), .c(t_6044), .d(t_11323), .cin(t_11325), .o(t_11326), .co(t_11327), .cout(t_11328));
compressor_3_2 u1_3941(.a(t_9508), .b(t_9505), .cin(t_9519), .o(t_11329), .cout(t_11330));
compressor_4_2 u2_3942(.a(t_9524), .b(t_9521), .c(t_6061), .d(t_11328), .cin(t_11330), .o(t_11331), .co(t_11332), .cout(t_11333));
compressor_3_2 u1_3943(.a(t_9517), .b(t_9514), .cin(t_9527), .o(t_11334), .cout(t_11335));
compressor_4_2 u2_3944(.a(t_9532), .b(t_9529), .c(t_6078), .d(t_11333), .cin(t_11335), .o(t_11336), .co(t_11337), .cout(t_11338));
compressor_3_2 u1_3945(.a(t_9525), .b(t_9522), .cin(t_9535), .o(t_11339), .cout(t_11340));
compressor_4_2 u2_3946(.a(t_9540), .b(t_9537), .c(t_6095), .d(t_11338), .cin(t_11340), .o(t_11341), .co(t_11342), .cout(t_11343));
compressor_3_2 u1_3947(.a(t_9533), .b(t_9530), .cin(t_9543), .o(t_11344), .cout(t_11345));
compressor_4_2 u2_3948(.a(t_9548), .b(t_9545), .c(t_6112), .d(t_11343), .cin(t_11345), .o(t_11346), .co(t_11347), .cout(t_11348));
compressor_3_2 u1_3949(.a(t_9541), .b(t_9538), .cin(t_9551), .o(t_11349), .cout(t_11350));
compressor_4_2 u2_3950(.a(t_9559), .b(t_9556), .c(t_9553), .d(t_11348), .cin(t_11350), .o(t_11351), .co(t_11352), .cout(t_11353));
half_adder u0_3951(.a(t_9549), .b(t_9546), .o(t_11354), .cout(t_11355));
compressor_4_2 u2_3952(.a(t_9564), .b(t_9561), .c(t_6144), .d(t_11353), .cin(t_11355), .o(t_11356), .co(t_11357), .cout(t_11358));
compressor_3_2 u1_3953(.a(t_9557), .b(t_9554), .cin(t_9567), .o(t_11359), .cout(t_11360));
compressor_4_2 u2_3954(.a(t_9575), .b(t_9572), .c(t_9569), .d(t_11358), .cin(t_11360), .o(t_11361), .co(t_11362), .cout(t_11363));
half_adder u0_3955(.a(t_9565), .b(t_9562), .o(t_11364), .cout(t_11365));
compressor_4_2 u2_3956(.a(t_9583), .b(t_9580), .c(t_9577), .d(t_11363), .cin(t_11365), .o(t_11366), .co(t_11367), .cout(t_11368));
half_adder u0_3957(.a(t_9573), .b(t_9570), .o(t_11369), .cout(t_11370));
compressor_4_2 u2_3958(.a(t_9591), .b(t_9588), .c(t_9585), .d(t_11368), .cin(t_11370), .o(t_11371), .co(t_11372), .cout(t_11373));
half_adder u0_3959(.a(t_9581), .b(t_9578), .o(t_11374), .cout(t_11375));
compressor_4_2 u2_3960(.a(t_9599), .b(t_9596), .c(t_9593), .d(t_11373), .cin(t_11375), .o(t_11376), .co(t_11377), .cout(t_11378));
half_adder u0_3961(.a(t_9589), .b(t_9586), .o(t_11379), .cout(t_11380));
compressor_4_2 u2_3962(.a(t_9607), .b(t_9604), .c(t_9601), .d(t_11378), .cin(t_11380), .o(t_11381), .co(t_11382), .cout(t_11383));
half_adder u0_3963(.a(t_9597), .b(t_9594), .o(t_11384), .cout(t_11385));
compressor_4_2 u2_3964(.a(t_9615), .b(t_9612), .c(t_9609), .d(t_11383), .cin(t_11385), .o(t_11386), .co(t_11387), .cout(t_11388));
half_adder u0_3965(.a(t_9605), .b(t_9602), .o(t_11389), .cout(t_11390));
compressor_4_2 u2_3966(.a(t_9620), .b(t_9617), .c(t_6240), .d(t_11388), .cin(t_11390), .o(t_11391), .co(t_11392), .cout(t_11393));
half_adder u0_3967(.a(t_9613), .b(t_9610), .o(t_11394), .cout(t_11395));
compressor_4_2 u2_3968(.a(t_9626), .b(t_9623), .c(t_6252), .d(t_11393), .cin(t_11395), .o(t_11396), .co(t_11397), .cout(t_11398));
half_adder u0_3969(.a(t_9621), .b(t_9618), .o(t_11399), .cout(t_11400));
compressor_4_2 u2_3970(.a(t_9624), .b(t_9632), .c(t_9629), .d(t_11398), .cin(t_11400), .o(t_11401), .co(t_11402), .cout(t_11403));
compressor_4_2 u2_3971(.a(t_9630), .b(t_9638), .c(t_9635), .d(t_6272), .cin(t_11403), .o(t_11404), .co(t_11405), .cout(t_11406));
compressor_4_2 u2_3972(.a(t_9636), .b(t_9643), .c(t_9640), .d(t_6283), .cin(t_11406), .o(t_11407), .co(t_11408), .cout(t_11409));
compressor_4_2 u2_3973(.a(t_9641), .b(t_9648), .c(t_9645), .d(t_6294), .cin(t_11409), .o(t_11410), .co(t_11411), .cout(t_11412));
compressor_4_2 u2_3974(.a(t_9646), .b(t_9653), .c(t_9650), .d(t_6305), .cin(t_11412), .o(t_11413), .co(t_11414), .cout(t_11415));
compressor_4_2 u2_3975(.a(t_9651), .b(t_9658), .c(t_9655), .d(t_6316), .cin(t_11415), .o(t_11416), .co(t_11417), .cout(t_11418));
compressor_3_2 u1_3976(.a(t_9663), .b(t_9660), .cin(t_11418), .o(t_11419), .cout(t_11420));
compressor_3_2 u1_3977(.a(t_9668), .b(t_9665), .cin(t_6336), .o(t_11421), .cout(t_11422));
compressor_3_2 u1_3978(.a(t_9666), .b(t_9673), .cin(t_9670), .o(t_11423), .cout(t_11424));
compressor_3_2 u1_3979(.a(t_9671), .b(t_9678), .cin(t_9675), .o(t_11425), .cout(t_11426));
compressor_3_2 u1_3980(.a(t_9676), .b(t_9683), .cin(t_9680), .o(t_11427), .cout(t_11428));
compressor_3_2 u1_3981(.a(t_9681), .b(t_9688), .cin(t_9685), .o(t_11429), .cout(t_11430));
compressor_3_2 u1_3982(.a(t_9686), .b(t_9693), .cin(t_9690), .o(t_11431), .cout(t_11432));
compressor_3_2 u1_3983(.a(t_9691), .b(t_9698), .cin(t_9695), .o(t_11433), .cout(t_11434));
compressor_3_2 u1_3984(.a(t_9696), .b(t_9700), .cin(t_6390), .o(t_11435), .cout(t_11436));
compressor_3_2 u1_3985(.a(t_9701), .b(t_9703), .cin(t_6396), .o(t_11437), .cout(t_11438));
half_adder u0_3986(.a(t_9704), .b(t_9706), .o(t_11439), .cout(t_11440));
compressor_3_2 u1_3987(.a(t_9707), .b(t_9709), .cin(t_6404), .o(t_11441), .cout(t_11442));
half_adder u0_3988(.a(t_9710), .b(t_9711), .o(t_11443), .cout(t_11444));
half_adder u0_3989(.a(t_9712), .b(t_9713), .o(t_11445), .cout(t_11446));
half_adder u0_3990(.a(t_9714), .b(t_9715), .o(t_11447), .cout(t_11448));
half_adder u0_3991(.a(t_9716), .b(t_9717), .o(t_11449), .cout(t_11450));
half_adder u0_3992(.a(t_9718), .b(t_9719), .o(t_11451), .cout(t_11452));
half_adder u0_3993(.a(t_9720), .b(t_9721), .o(t_11453), .cout(t_11454));
half_adder u0_3994(.a(t_9722), .b(t_9723), .o(t_11455), .cout(t_11456));
half_adder u0_3995(.a(t_9724), .b(t_9725), .o(t_11457), .cout(t_11458));
half_adder u0_3996(.a(t_9726), .b(t_9727), .o(t_11459), .cout());

/* u0_3997 Output nets */
wire t_11460,  t_11461;
/* u0_3998 Output nets */
wire t_11462,  t_11463;
/* u0_3999 Output nets */
wire t_11464,  t_11465;
/* u0_4000 Output nets */
wire t_11466,  t_11467;
/* u0_4001 Output nets */
wire t_11468,  t_11469;
/* u0_4002 Output nets */
wire t_11470,  t_11471;
/* u0_4003 Output nets */
wire t_11472,  t_11473;
/* u0_4004 Output nets */
wire t_11474,  t_11475;
/* u0_4005 Output nets */
wire t_11476,  t_11477;
/* u0_4006 Output nets */
wire t_11478,  t_11479;
/* u0_4007 Output nets */
wire t_11480,  t_11481;
/* u0_4008 Output nets */
wire t_11482,  t_11483;
/* u0_4009 Output nets */
wire t_11484,  t_11485;
/* u0_4010 Output nets */
wire t_11486,  t_11487;
/* u0_4011 Output nets */
wire t_11488,  t_11489;
/* u1_4012 Output nets */
wire t_11490,  t_11491;
/* u0_4013 Output nets */
wire t_11492,  t_11493;
/* u0_4014 Output nets */
wire t_11494,  t_11495;
/* u1_4015 Output nets */
wire t_11496,  t_11497;
/* u0_4016 Output nets */
wire t_11498,  t_11499;
/* u0_4017 Output nets */
wire t_11500,  t_11501;
/* u0_4018 Output nets */
wire t_11502,  t_11503;
/* u0_4019 Output nets */
wire t_11504,  t_11505;
/* u0_4020 Output nets */
wire t_11506,  t_11507;
/* u1_4021 Output nets */
wire t_11508,  t_11509;
/* u1_4022 Output nets */
wire t_11510,  t_11511;
/* u1_4023 Output nets */
wire t_11512,  t_11513;
/* u1_4024 Output nets */
wire t_11514,  t_11515;
/* u1_4025 Output nets */
wire t_11516,  t_11517;
/* u1_4026 Output nets */
wire t_11518,  t_11519;
/* u1_4027 Output nets */
wire t_11520,  t_11521;
/* u1_4028 Output nets */
wire t_11522,  t_11523;
/* u1_4029 Output nets */
wire t_11524,  t_11525;
/* u1_4030 Output nets */
wire t_11526,  t_11527;
/* u1_4031 Output nets */
wire t_11528,  t_11529;
/* u2_4032 Output nets */
wire t_11530,  t_11531,  t_11532;
/* u1_4033 Output nets */
wire t_11533,  t_11534;
/* u1_4034 Output nets */
wire t_11535,  t_11536;
/* u1_4035 Output nets */
wire t_11537,  t_11538;
/* u1_4036 Output nets */
wire t_11539,  t_11540;
/* u2_4037 Output nets */
wire t_11541,  t_11542,  t_11543;
/* u2_4038 Output nets */
wire t_11544,  t_11545,  t_11546;
/* u2_4039 Output nets */
wire t_11547,  t_11548,  t_11549;
/* u2_4040 Output nets */
wire t_11550,  t_11551,  t_11552;
/* u2_4041 Output nets */
wire t_11553,  t_11554,  t_11555;
/* u1_4042 Output nets */
wire t_11556,  t_11557;
/* u2_4043 Output nets */
wire t_11558,  t_11559,  t_11560;
/* u2_4044 Output nets */
wire t_11561,  t_11562,  t_11563;
/* u1_4045 Output nets */
wire t_11564,  t_11565;
/* u1_4046 Output nets */
wire t_11566,  t_11567;
/* u2_4047 Output nets */
wire t_11568,  t_11569,  t_11570;
/* u2_4048 Output nets */
wire t_11571,  t_11572,  t_11573;
/* u2_4049 Output nets */
wire t_11574,  t_11575,  t_11576;
/* u2_4050 Output nets */
wire t_11577,  t_11578,  t_11579;
/* u2_4051 Output nets */
wire t_11580,  t_11581,  t_11582;
/* u2_4052 Output nets */
wire t_11583,  t_11584,  t_11585;
/* u2_4053 Output nets */
wire t_11586,  t_11587,  t_11588;
/* u2_4054 Output nets */
wire t_11589,  t_11590,  t_11591;
/* u2_4055 Output nets */
wire t_11592,  t_11593,  t_11594;
/* u2_4056 Output nets */
wire t_11595,  t_11596,  t_11597;
/* u2_4057 Output nets */
wire t_11598,  t_11599,  t_11600;
/* u2_4058 Output nets */
wire t_11601,  t_11602,  t_11603;
/* u2_4059 Output nets */
wire t_11604,  t_11605,  t_11606;
/* u2_4060 Output nets */
wire t_11607,  t_11608,  t_11609;
/* u2_4061 Output nets */
wire t_11610,  t_11611,  t_11612;
/* u2_4062 Output nets */
wire t_11613,  t_11614,  t_11615;
/* u2_4063 Output nets */
wire t_11616,  t_11617,  t_11618;
/* u2_4064 Output nets */
wire t_11619,  t_11620,  t_11621;
/* u0_4065 Output nets */
wire t_11622,  t_11623;
/* u2_4066 Output nets */
wire t_11624,  t_11625,  t_11626;
/* u0_4067 Output nets */
wire t_11627,  t_11628;
/* u2_4068 Output nets */
wire t_11629,  t_11630,  t_11631;
/* u0_4069 Output nets */
wire t_11632,  t_11633;
/* u2_4070 Output nets */
wire t_11634,  t_11635,  t_11636;
/* u0_4071 Output nets */
wire t_11637,  t_11638;
/* u2_4072 Output nets */
wire t_11639,  t_11640,  t_11641;
/* u0_4073 Output nets */
wire t_11642,  t_11643;
/* u2_4074 Output nets */
wire t_11644,  t_11645,  t_11646;
/* u1_4075 Output nets */
wire t_11647,  t_11648;
/* u2_4076 Output nets */
wire t_11649,  t_11650,  t_11651;
/* u1_4077 Output nets */
wire t_11652,  t_11653;
/* u2_4078 Output nets */
wire t_11654,  t_11655,  t_11656;
/* u1_4079 Output nets */
wire t_11657,  t_11658;
/* u2_4080 Output nets */
wire t_11659,  t_11660,  t_11661;
/* u1_4081 Output nets */
wire t_11662,  t_11663;
/* u2_4082 Output nets */
wire t_11664,  t_11665,  t_11666;
/* u1_4083 Output nets */
wire t_11667,  t_11668;
/* u2_4084 Output nets */
wire t_11669,  t_11670,  t_11671;
/* u0_4085 Output nets */
wire t_11672,  t_11673;
/* u2_4086 Output nets */
wire t_11674,  t_11675,  t_11676;
/* u1_4087 Output nets */
wire t_11677,  t_11678;
/* u2_4088 Output nets */
wire t_11679,  t_11680,  t_11681;
/* u1_4089 Output nets */
wire t_11682,  t_11683;
/* u2_4090 Output nets */
wire t_11684,  t_11685,  t_11686;
/* u0_4091 Output nets */
wire t_11687,  t_11688;
/* u2_4092 Output nets */
wire t_11689,  t_11690,  t_11691;
/* u1_4093 Output nets */
wire t_11692,  t_11693;
/* u2_4094 Output nets */
wire t_11694,  t_11695,  t_11696;
/* u1_4095 Output nets */
wire t_11697,  t_11698;
/* u2_4096 Output nets */
wire t_11699,  t_11700,  t_11701;
/* u1_4097 Output nets */
wire t_11702,  t_11703;
/* u2_4098 Output nets */
wire t_11704,  t_11705,  t_11706;
/* u1_4099 Output nets */
wire t_11707,  t_11708;
/* u2_4100 Output nets */
wire t_11709,  t_11710,  t_11711;
/* u1_4101 Output nets */
wire t_11712,  t_11713;
/* u2_4102 Output nets */
wire t_11714,  t_11715,  t_11716;
/* u1_4103 Output nets */
wire t_11717,  t_11718;
/* u2_4104 Output nets */
wire t_11719,  t_11720,  t_11721;
/* u1_4105 Output nets */
wire t_11722,  t_11723;
/* u2_4106 Output nets */
wire t_11724,  t_11725,  t_11726;
/* u1_4107 Output nets */
wire t_11727,  t_11728;
/* u2_4108 Output nets */
wire t_11729,  t_11730,  t_11731;
/* u1_4109 Output nets */
wire t_11732,  t_11733;
/* u2_4110 Output nets */
wire t_11734,  t_11735,  t_11736;
/* u1_4111 Output nets */
wire t_11737,  t_11738;
/* u2_4112 Output nets */
wire t_11739,  t_11740,  t_11741;
/* u1_4113 Output nets */
wire t_11742,  t_11743;
/* u2_4114 Output nets */
wire t_11744,  t_11745,  t_11746;
/* u1_4115 Output nets */
wire t_11747,  t_11748;
/* u2_4116 Output nets */
wire t_11749,  t_11750,  t_11751;
/* u1_4117 Output nets */
wire t_11752,  t_11753;
/* u2_4118 Output nets */
wire t_11754,  t_11755,  t_11756;
/* u1_4119 Output nets */
wire t_11757,  t_11758;
/* u2_4120 Output nets */
wire t_11759,  t_11760,  t_11761;
/* u1_4121 Output nets */
wire t_11762,  t_11763;
/* u2_4122 Output nets */
wire t_11764,  t_11765,  t_11766;
/* u1_4123 Output nets */
wire t_11767,  t_11768;
/* u2_4124 Output nets */
wire t_11769,  t_11770,  t_11771;
/* u1_4125 Output nets */
wire t_11772,  t_11773;
/* u2_4126 Output nets */
wire t_11774,  t_11775,  t_11776;
/* u1_4127 Output nets */
wire t_11777,  t_11778;
/* u2_4128 Output nets */
wire t_11779,  t_11780,  t_11781;
/* u2_4129 Output nets */
wire t_11782,  t_11783,  t_11784;
/* u2_4130 Output nets */
wire t_11785,  t_11786,  t_11787;
/* u1_4131 Output nets */
wire t_11788,  t_11789;
/* u2_4132 Output nets */
wire t_11790,  t_11791,  t_11792;
/* u1_4133 Output nets */
wire t_11793,  t_11794;
/* u2_4134 Output nets */
wire t_11795,  t_11796,  t_11797;
/* u1_4135 Output nets */
wire t_11798,  t_11799;
/* u2_4136 Output nets */
wire t_11800,  t_11801,  t_11802;
/* u1_4137 Output nets */
wire t_11803,  t_11804;
/* u2_4138 Output nets */
wire t_11805,  t_11806,  t_11807;
/* u2_4139 Output nets */
wire t_11808,  t_11809,  t_11810;
/* u2_4140 Output nets */
wire t_11811,  t_11812,  t_11813;
/* u2_4141 Output nets */
wire t_11814,  t_11815,  t_11816;
/* u2_4142 Output nets */
wire t_11817,  t_11818,  t_11819;
/* u2_4143 Output nets */
wire t_11820,  t_11821,  t_11822;
/* u2_4144 Output nets */
wire t_11823,  t_11824,  t_11825;
/* u2_4145 Output nets */
wire t_11826,  t_11827,  t_11828;
/* u2_4146 Output nets */
wire t_11829,  t_11830,  t_11831;
/* u2_4147 Output nets */
wire t_11832,  t_11833,  t_11834;
/* u2_4148 Output nets */
wire t_11835,  t_11836,  t_11837;
/* u1_4149 Output nets */
wire t_11838,  t_11839;
/* u2_4150 Output nets */
wire t_11840,  t_11841,  t_11842;
/* u2_4151 Output nets */
wire t_11843,  t_11844,  t_11845;
/* u2_4152 Output nets */
wire t_11846,  t_11847,  t_11848;
/* u2_4153 Output nets */
wire t_11849,  t_11850,  t_11851;
/* u2_4154 Output nets */
wire t_11852,  t_11853,  t_11854;
/* u1_4155 Output nets */
wire t_11855,  t_11856;
/* u2_4156 Output nets */
wire t_11857,  t_11858,  t_11859;
/* u2_4157 Output nets */
wire t_11860,  t_11861,  t_11862;
/* u2_4158 Output nets */
wire t_11863,  t_11864,  t_11865;
/* u2_4159 Output nets */
wire t_11866,  t_11867,  t_11868;
/* u2_4160 Output nets */
wire t_11869,  t_11870,  t_11871;
/* u2_4161 Output nets */
wire t_11872,  t_11873,  t_11874;
/* u2_4162 Output nets */
wire t_11875,  t_11876,  t_11877;
/* u2_4163 Output nets */
wire t_11878,  t_11879,  t_11880;
/* u2_4164 Output nets */
wire t_11881,  t_11882,  t_11883;
/* u2_4165 Output nets */
wire t_11884,  t_11885,  t_11886;
/* u2_4166 Output nets */
wire t_11887,  t_11888,  t_11889;
/* u2_4167 Output nets */
wire t_11890,  t_11891,  t_11892;
/* u2_4168 Output nets */
wire t_11893,  t_11894,  t_11895;
/* u2_4169 Output nets */
wire t_11896,  t_11897,  t_11898;
/* u2_4170 Output nets */
wire t_11899,  t_11900,  t_11901;
/* u2_4171 Output nets */
wire t_11902,  t_11903,  t_11904;
/* u2_4172 Output nets */
wire t_11905,  t_11906,  t_11907;
/* u2_4173 Output nets */
wire t_11908,  t_11909,  t_11910;
/* u2_4174 Output nets */
wire t_11911,  t_11912,  t_11913;
/* u2_4175 Output nets */
wire t_11914,  t_11915,  t_11916;
/* u2_4176 Output nets */
wire t_11917,  t_11918,  t_11919;
/* u2_4177 Output nets */
wire t_11920,  t_11921,  t_11922;
/* u2_4178 Output nets */
wire t_11923,  t_11924,  t_11925;
/* u2_4179 Output nets */
wire t_11926,  t_11927,  t_11928;
/* u2_4180 Output nets */
wire t_11929,  t_11930,  t_11931;
/* u2_4181 Output nets */
wire t_11932,  t_11933,  t_11934;
/* u2_4182 Output nets */
wire t_11935,  t_11936,  t_11937;
/* u2_4183 Output nets */
wire t_11938,  t_11939,  t_11940;
/* u2_4184 Output nets */
wire t_11941,  t_11942,  t_11943;
/* u2_4185 Output nets */
wire t_11944,  t_11945,  t_11946;
/* u2_4186 Output nets */
wire t_11947,  t_11948,  t_11949;
/* u2_4187 Output nets */
wire t_11950,  t_11951,  t_11952;
/* u2_4188 Output nets */
wire t_11953,  t_11954,  t_11955;
/* u2_4189 Output nets */
wire t_11956,  t_11957,  t_11958;
/* u2_4190 Output nets */
wire t_11959,  t_11960,  t_11961;
/* u2_4191 Output nets */
wire t_11962,  t_11963,  t_11964;
/* u2_4192 Output nets */
wire t_11965,  t_11966,  t_11967;
/* u2_4193 Output nets */
wire t_11968,  t_11969,  t_11970;
/* u2_4194 Output nets */
wire t_11971,  t_11972,  t_11973;
/* u1_4195 Output nets */
wire t_11974,  t_11975;
/* u2_4196 Output nets */
wire t_11976,  t_11977,  t_11978;
/* u2_4197 Output nets */
wire t_11979,  t_11980,  t_11981;
/* u2_4198 Output nets */
wire t_11982,  t_11983,  t_11984;
/* u2_4199 Output nets */
wire t_11985,  t_11986,  t_11987;
/* u2_4200 Output nets */
wire t_11988,  t_11989,  t_11990;
/* u2_4201 Output nets */
wire t_11991,  t_11992,  t_11993;
/* u2_4202 Output nets */
wire t_11994,  t_11995,  t_11996;
/* u2_4203 Output nets */
wire t_11997,  t_11998,  t_11999;
/* u2_4204 Output nets */
wire t_12000,  t_12001,  t_12002;
/* u2_4205 Output nets */
wire t_12003,  t_12004,  t_12005;
/* u2_4206 Output nets */
wire t_12006,  t_12007,  t_12008;
/* u2_4207 Output nets */
wire t_12009,  t_12010,  t_12011;
/* u2_4208 Output nets */
wire t_12012,  t_12013,  t_12014;
/* u2_4209 Output nets */
wire t_12015,  t_12016,  t_12017;
/* u2_4210 Output nets */
wire t_12018,  t_12019,  t_12020;
/* u2_4211 Output nets */
wire t_12021,  t_12022,  t_12023;
/* u2_4212 Output nets */
wire t_12024,  t_12025,  t_12026;
/* u1_4213 Output nets */
wire t_12027,  t_12028;
/* u2_4214 Output nets */
wire t_12029,  t_12030,  t_12031;
/* u2_4215 Output nets */
wire t_12032,  t_12033,  t_12034;
/* u2_4216 Output nets */
wire t_12035,  t_12036,  t_12037;
/* u1_4217 Output nets */
wire t_12038,  t_12039;
/* u2_4218 Output nets */
wire t_12040,  t_12041,  t_12042;
/* u1_4219 Output nets */
wire t_12043,  t_12044;
/* u2_4220 Output nets */
wire t_12045,  t_12046,  t_12047;
/* u1_4221 Output nets */
wire t_12048,  t_12049;
/* u2_4222 Output nets */
wire t_12050,  t_12051,  t_12052;
/* u1_4223 Output nets */
wire t_12053,  t_12054;
/* u2_4224 Output nets */
wire t_12055,  t_12056,  t_12057;
/* u1_4225 Output nets */
wire t_12058,  t_12059;
/* u2_4226 Output nets */
wire t_12060,  t_12061,  t_12062;
/* u1_4227 Output nets */
wire t_12063,  t_12064;
/* u2_4228 Output nets */
wire t_12065,  t_12066,  t_12067;
/* u1_4229 Output nets */
wire t_12068,  t_12069;
/* u2_4230 Output nets */
wire t_12070,  t_12071,  t_12072;
/* u1_4231 Output nets */
wire t_12073,  t_12074;
/* u2_4232 Output nets */
wire t_12075,  t_12076,  t_12077;
/* u1_4233 Output nets */
wire t_12078,  t_12079;
/* u2_4234 Output nets */
wire t_12080,  t_12081,  t_12082;
/* u1_4235 Output nets */
wire t_12083,  t_12084;
/* u2_4236 Output nets */
wire t_12085,  t_12086,  t_12087;
/* u1_4237 Output nets */
wire t_12088,  t_12089;
/* u2_4238 Output nets */
wire t_12090,  t_12091,  t_12092;
/* u1_4239 Output nets */
wire t_12093,  t_12094;
/* u2_4240 Output nets */
wire t_12095,  t_12096,  t_12097;
/* u1_4241 Output nets */
wire t_12098,  t_12099;
/* u2_4242 Output nets */
wire t_12100,  t_12101,  t_12102;
/* u1_4243 Output nets */
wire t_12103,  t_12104;
/* u2_4244 Output nets */
wire t_12105,  t_12106,  t_12107;
/* u1_4245 Output nets */
wire t_12108,  t_12109;
/* u2_4246 Output nets */
wire t_12110,  t_12111,  t_12112;
/* u1_4247 Output nets */
wire t_12113,  t_12114;
/* u2_4248 Output nets */
wire t_12115,  t_12116,  t_12117;
/* u1_4249 Output nets */
wire t_12118,  t_12119;
/* u2_4250 Output nets */
wire t_12120,  t_12121,  t_12122;
/* u1_4251 Output nets */
wire t_12123,  t_12124;
/* u2_4252 Output nets */
wire t_12125,  t_12126,  t_12127;
/* u1_4253 Output nets */
wire t_12128,  t_12129;
/* u2_4254 Output nets */
wire t_12130,  t_12131,  t_12132;
/* u1_4255 Output nets */
wire t_12133,  t_12134;
/* u2_4256 Output nets */
wire t_12135,  t_12136,  t_12137;
/* u1_4257 Output nets */
wire t_12138,  t_12139;
/* u2_4258 Output nets */
wire t_12140,  t_12141,  t_12142;
/* u0_4259 Output nets */
wire t_12143,  t_12144;
/* u2_4260 Output nets */
wire t_12145,  t_12146,  t_12147;
/* u1_4261 Output nets */
wire t_12148,  t_12149;
/* u2_4262 Output nets */
wire t_12150,  t_12151,  t_12152;
/* u1_4263 Output nets */
wire t_12153,  t_12154;
/* u2_4264 Output nets */
wire t_12155,  t_12156,  t_12157;
/* u1_4265 Output nets */
wire t_12158,  t_12159;
/* u2_4266 Output nets */
wire t_12160,  t_12161,  t_12162;
/* u1_4267 Output nets */
wire t_12163,  t_12164;
/* u2_4268 Output nets */
wire t_12165,  t_12166,  t_12167;
/* u1_4269 Output nets */
wire t_12168,  t_12169;
/* u2_4270 Output nets */
wire t_12170,  t_12171,  t_12172;
/* u1_4271 Output nets */
wire t_12173,  t_12174;
/* u2_4272 Output nets */
wire t_12175,  t_12176,  t_12177;
/* u1_4273 Output nets */
wire t_12178,  t_12179;
/* u2_4274 Output nets */
wire t_12180,  t_12181,  t_12182;
/* u1_4275 Output nets */
wire t_12183,  t_12184;
/* u2_4276 Output nets */
wire t_12185,  t_12186,  t_12187;
/* u0_4277 Output nets */
wire t_12188,  t_12189;
/* u2_4278 Output nets */
wire t_12190,  t_12191,  t_12192;
/* u1_4279 Output nets */
wire t_12193,  t_12194;
/* u2_4280 Output nets */
wire t_12195,  t_12196,  t_12197;
/* u0_4281 Output nets */
wire t_12198,  t_12199;
/* u2_4282 Output nets */
wire t_12200,  t_12201,  t_12202;
/* u0_4283 Output nets */
wire t_12203,  t_12204;
/* u2_4284 Output nets */
wire t_12205,  t_12206,  t_12207;
/* u0_4285 Output nets */
wire t_12208,  t_12209;
/* u2_4286 Output nets */
wire t_12210,  t_12211,  t_12212;
/* u0_4287 Output nets */
wire t_12213,  t_12214;
/* u2_4288 Output nets */
wire t_12215,  t_12216,  t_12217;
/* u0_4289 Output nets */
wire t_12218,  t_12219;
/* u2_4290 Output nets */
wire t_12220,  t_12221,  t_12222;
/* u0_4291 Output nets */
wire t_12223,  t_12224;
/* u2_4292 Output nets */
wire t_12225,  t_12226,  t_12227;
/* u0_4293 Output nets */
wire t_12228,  t_12229;
/* u2_4294 Output nets */
wire t_12230,  t_12231,  t_12232;
/* u0_4295 Output nets */
wire t_12233,  t_12234;
/* u2_4296 Output nets */
wire t_12235,  t_12236,  t_12237;
/* u0_4297 Output nets */
wire t_12238,  t_12239;
/* u2_4298 Output nets */
wire t_12240,  t_12241,  t_12242;
/* u0_4299 Output nets */
wire t_12243,  t_12244;
/* u2_4300 Output nets */
wire t_12245,  t_12246,  t_12247;
/* u0_4301 Output nets */
wire t_12248,  t_12249;
/* u2_4302 Output nets */
wire t_12250,  t_12251,  t_12252;
/* u0_4303 Output nets */
wire t_12253,  t_12254;
/* u2_4304 Output nets */
wire t_12255,  t_12256,  t_12257;
/* u0_4305 Output nets */
wire t_12258,  t_12259;
/* u2_4306 Output nets */
wire t_12260,  t_12261,  t_12262;
/* u0_4307 Output nets */
wire t_12263,  t_12264;
/* u2_4308 Output nets */
wire t_12265,  t_12266,  t_12267;
/* u0_4309 Output nets */
wire t_12268,  t_12269;
/* u2_4310 Output nets */
wire t_12270,  t_12271,  t_12272;
/* u0_4311 Output nets */
wire t_12273,  t_12274;
/* u2_4312 Output nets */
wire t_12275,  t_12276,  t_12277;
/* u2_4313 Output nets */
wire t_12278,  t_12279,  t_12280;
/* u2_4314 Output nets */
wire t_12281,  t_12282,  t_12283;
/* u2_4315 Output nets */
wire t_12284,  t_12285,  t_12286;
/* u2_4316 Output nets */
wire t_12287,  t_12288,  t_12289;
/* u1_4317 Output nets */
wire t_12290,  t_12291;
/* u2_4318 Output nets */
wire t_12292,  t_12293,  t_12294;
/* u2_4319 Output nets */
wire t_12295,  t_12296,  t_12297;
/* u2_4320 Output nets */
wire t_12298,  t_12299,  t_12300;
/* u2_4321 Output nets */
wire t_12301,  t_12302,  t_12303;
/* u2_4322 Output nets */
wire t_12304,  t_12305,  t_12306;
/* u2_4323 Output nets */
wire t_12307,  t_12308,  t_12309;
/* u2_4324 Output nets */
wire t_12310,  t_12311,  t_12312;
/* u2_4325 Output nets */
wire t_12313,  t_12314,  t_12315;
/* u1_4326 Output nets */
wire t_12316,  t_12317;
/* u1_4327 Output nets */
wire t_12318,  t_12319;
/* u1_4328 Output nets */
wire t_12320,  t_12321;
/* u1_4329 Output nets */
wire t_12322,  t_12323;
/* u1_4330 Output nets */
wire t_12324,  t_12325;
/* u1_4331 Output nets */
wire t_12326,  t_12327;
/* u1_4332 Output nets */
wire t_12328,  t_12329;
/* u1_4333 Output nets */
wire t_12330,  t_12331;
/* u1_4334 Output nets */
wire t_12332,  t_12333;
/* u1_4335 Output nets */
wire t_12334,  t_12335;
/* u1_4336 Output nets */
wire t_12336,  t_12337;
/* u1_4337 Output nets */
wire t_12338,  t_12339;
/* u1_4338 Output nets */
wire t_12340,  t_12341;
/* u1_4339 Output nets */
wire t_12342,  t_12343;
/* u1_4340 Output nets */
wire t_12344,  t_12345;
/* u1_4341 Output nets */
wire t_12346,  t_12347;
/* u1_4342 Output nets */
wire t_12348,  t_12349;
/* u1_4343 Output nets */
wire t_12350,  t_12351;
/* u0_4344 Output nets */
wire t_12352,  t_12353;
/* u0_4345 Output nets */
wire t_12354,  t_12355;
/* u0_4346 Output nets */
wire t_12356,  t_12357;
/* u0_4347 Output nets */
wire t_12358,  t_12359;
/* u1_4348 Output nets */
wire t_12360,  t_12361;
/* u1_4349 Output nets */
wire t_12362,  t_12363;
/* u0_4350 Output nets */
wire t_12364,  t_12365;
/* u0_4351 Output nets */
wire t_12366,  t_12367;
/* u0_4352 Output nets */
wire t_12368,  t_12369;
/* u0_4353 Output nets */
wire t_12370,  t_12371;
/* u0_4354 Output nets */
wire t_12372,  t_12373;
/* u0_4355 Output nets */
wire t_12374,  t_12375;
/* u0_4356 Output nets */
wire t_12376,  t_12377;
/* u0_4357 Output nets */
wire t_12378,  t_12379;
/* u0_4358 Output nets */
wire t_12380,  t_12381;
/* u0_4359 Output nets */
wire t_12382,  t_12383;
/* u0_4360 Output nets */
wire t_12384,  t_12385;
/* u0_4361 Output nets */
wire t_12386,  t_12387;
/* u0_4362 Output nets */
wire t_12388,  t_12389;
/* u0_4363 Output nets */
wire t_12390,  t_12391;
/* u0_4364 Output nets */
wire t_12392,  t_12393;
/* u0_4365 Output nets */
wire t_12394,  t_12395;
/* u0_4366 Output nets */
wire t_12396,  t_12397;
/* u0_4367 Output nets */
wire t_12398,  t_12399;
/* u0_4368 Output nets */
wire t_12400;

/* compress stage 4 */
half_adder u0_3997(.a(t_9729), .b(t_6443), .o(t_11460), .cout(t_11461));
half_adder u0_3998(.a(t_9731), .b(t_6445), .o(t_11462), .cout(t_11463));
half_adder u0_3999(.a(t_9733), .b(t_9734), .o(t_11464), .cout(t_11465));
half_adder u0_4000(.a(t_9735), .b(t_9736), .o(t_11466), .cout(t_11467));
half_adder u0_4001(.a(t_9737), .b(t_9738), .o(t_11468), .cout(t_11469));
half_adder u0_4002(.a(t_9739), .b(t_6455), .o(t_11470), .cout(t_11471));
half_adder u0_4003(.a(t_9741), .b(t_9742), .o(t_11472), .cout(t_11473));
half_adder u0_4004(.a(t_9743), .b(t_9744), .o(t_11474), .cout(t_11475));
half_adder u0_4005(.a(t_9745), .b(t_9746), .o(t_11476), .cout(t_11477));
half_adder u0_4006(.a(t_9747), .b(t_9748), .o(t_11478), .cout(t_11479));
half_adder u0_4007(.a(t_9749), .b(t_9750), .o(t_11480), .cout(t_11481));
half_adder u0_4008(.a(t_9751), .b(t_9752), .o(t_11482), .cout(t_11483));
half_adder u0_4009(.a(t_9753), .b(t_9754), .o(t_11484), .cout(t_11485));
half_adder u0_4010(.a(t_9755), .b(t_9756), .o(t_11486), .cout(t_11487));
half_adder u0_4011(.a(t_9757), .b(t_9758), .o(t_11488), .cout(t_11489));
compressor_3_2 u1_4012(.a(t_9761), .b(t_9763), .cin(t_6493), .o(t_11490), .cout(t_11491));
half_adder u0_4013(.a(t_9764), .b(t_9765), .o(t_11492), .cout(t_11493));
half_adder u0_4014(.a(t_9768), .b(t_9770), .o(t_11494), .cout(t_11495));
compressor_3_2 u1_4015(.a(t_9771), .b(t_9773), .cin(t_6513), .o(t_11496), .cout(t_11497));
half_adder u0_4016(.a(t_9774), .b(t_9775), .o(t_11498), .cout(t_11499));
half_adder u0_4017(.a(t_9776), .b(t_9778), .o(t_11500), .cout(t_11501));
half_adder u0_4018(.a(t_9779), .b(t_9781), .o(t_11502), .cout(t_11503));
half_adder u0_4019(.a(t_9782), .b(t_9784), .o(t_11504), .cout(t_11505));
half_adder u0_4020(.a(t_9785), .b(t_9787), .o(t_11506), .cout(t_11507));
compressor_3_2 u1_4021(.a(t_9788), .b(t_9790), .cin(t_6549), .o(t_11508), .cout(t_11509));
compressor_3_2 u1_4022(.a(t_9791), .b(t_9793), .cin(t_6555), .o(t_11510), .cout(t_11511));
compressor_3_2 u1_4023(.a(t_9794), .b(t_9796), .cin(t_6561), .o(t_11512), .cout(t_11513));
compressor_3_2 u1_4024(.a(t_9797), .b(t_9799), .cin(t_6567), .o(t_11514), .cout(t_11515));
compressor_3_2 u1_4025(.a(t_9800), .b(t_9802), .cin(t_6575), .o(t_11516), .cout(t_11517));
compressor_3_2 u1_4026(.a(t_9803), .b(t_9808), .cin(t_9805), .o(t_11518), .cout(t_11519));
compressor_3_2 u1_4027(.a(t_9806), .b(t_9813), .cin(t_9810), .o(t_11520), .cout(t_11521));
compressor_3_2 u1_4028(.a(t_9811), .b(t_9818), .cin(t_9815), .o(t_11522), .cout(t_11523));
compressor_3_2 u1_4029(.a(t_9816), .b(t_9823), .cin(t_9820), .o(t_11524), .cout(t_11525));
compressor_3_2 u1_4030(.a(t_9821), .b(t_9828), .cin(t_9825), .o(t_11526), .cout(t_11527));
compressor_3_2 u1_4031(.a(t_9826), .b(t_9833), .cin(t_9830), .o(t_11528), .cout(t_11529));
compressor_4_2 u2_4032(.a(t_9831), .b(t_9838), .c(t_9835), .d(t_6634), .cin(t_11529), .o(t_11530), .co(t_11531), .cout(t_11532));
compressor_3_2 u1_4033(.a(t_9843), .b(t_9840), .cin(t_11532), .o(t_11533), .cout(t_11534));
compressor_3_2 u1_4034(.a(t_9841), .b(t_9848), .cin(t_9845), .o(t_11535), .cout(t_11536));
compressor_3_2 u1_4035(.a(t_9846), .b(t_9853), .cin(t_9850), .o(t_11537), .cout(t_11538));
compressor_3_2 u1_4036(.a(t_9851), .b(t_9858), .cin(t_9855), .o(t_11539), .cout(t_11540));
compressor_4_2 u2_4037(.a(t_9856), .b(t_9863), .c(t_9860), .d(t_6677), .cin(t_11540), .o(t_11541), .co(t_11542), .cout(t_11543));
compressor_4_2 u2_4038(.a(t_9861), .b(t_9868), .c(t_9865), .d(t_6686), .cin(t_11543), .o(t_11544), .co(t_11545), .cout(t_11546));
compressor_4_2 u2_4039(.a(t_9866), .b(t_9873), .c(t_9870), .d(t_6695), .cin(t_11546), .o(t_11547), .co(t_11548), .cout(t_11549));
compressor_4_2 u2_4040(.a(t_9871), .b(t_9878), .c(t_9875), .d(t_6704), .cin(t_11549), .o(t_11550), .co(t_11551), .cout(t_11552));
compressor_4_2 u2_4041(.a(t_9876), .b(t_9883), .c(t_9880), .d(t_6715), .cin(t_11552), .o(t_11553), .co(t_11554), .cout(t_11555));
compressor_3_2 u1_4042(.a(t_9888), .b(t_9885), .cin(t_11555), .o(t_11556), .cout(t_11557));
compressor_4_2 u2_4043(.a(t_9889), .b(t_9886), .c(t_9894), .d(t_9891), .cin(t_6737), .o(t_11558), .co(t_11559), .cout(t_11560));
compressor_4_2 u2_4044(.a(t_9892), .b(t_9899), .c(t_9896), .d(t_6748), .cin(t_11560), .o(t_11561), .co(t_11562), .cout(t_11563));
compressor_3_2 u1_4045(.a(t_9904), .b(t_9901), .cin(t_11563), .o(t_11564), .cout(t_11565));
compressor_3_2 u1_4046(.a(t_9902), .b(t_9910), .cin(t_9907), .o(t_11566), .cout(t_11567));
compressor_4_2 u2_4047(.a(t_9908), .b(t_9916), .c(t_9913), .d(t_6781), .cin(t_11567), .o(t_11568), .co(t_11569), .cout(t_11570));
compressor_4_2 u2_4048(.a(t_9914), .b(t_9921), .c(t_9918), .d(t_6795), .cin(t_11570), .o(t_11571), .co(t_11572), .cout(t_11573));
compressor_4_2 u2_4049(.a(t_9922), .b(t_9919), .c(t_9927), .d(t_9924), .cin(t_11573), .o(t_11574), .co(t_11575), .cout(t_11576));
compressor_4_2 u2_4050(.a(t_9928), .b(t_9925), .c(t_9933), .d(t_9930), .cin(t_11576), .o(t_11577), .co(t_11578), .cout(t_11579));
compressor_4_2 u2_4051(.a(t_9934), .b(t_9931), .c(t_9939), .d(t_9936), .cin(t_11579), .o(t_11580), .co(t_11581), .cout(t_11582));
compressor_4_2 u2_4052(.a(t_9940), .b(t_9937), .c(t_9945), .d(t_9942), .cin(t_11582), .o(t_11583), .co(t_11584), .cout(t_11585));
compressor_4_2 u2_4053(.a(t_9943), .b(t_9951), .c(t_9948), .d(t_6853), .cin(t_11585), .o(t_11586), .co(t_11587), .cout(t_11588));
compressor_4_2 u2_4054(.a(t_9949), .b(t_9957), .c(t_9954), .d(t_6865), .cin(t_11588), .o(t_11589), .co(t_11590), .cout(t_11591));
compressor_4_2 u2_4055(.a(t_9955), .b(t_9963), .c(t_9960), .d(t_6877), .cin(t_11591), .o(t_11592), .co(t_11593), .cout(t_11594));
compressor_4_2 u2_4056(.a(t_9961), .b(t_9969), .c(t_9966), .d(t_6889), .cin(t_11594), .o(t_11595), .co(t_11596), .cout(t_11597));
compressor_4_2 u2_4057(.a(t_9967), .b(t_9975), .c(t_9972), .d(t_6903), .cin(t_11597), .o(t_11598), .co(t_11599), .cout(t_11600));
compressor_4_2 u2_4058(.a(t_9973), .b(t_9984), .c(t_9981), .d(t_9978), .cin(t_11600), .o(t_11601), .co(t_11602), .cout(t_11603));
compressor_4_2 u2_4059(.a(t_9979), .b(t_9992), .c(t_9989), .d(t_9986), .cin(t_11603), .o(t_11604), .co(t_11605), .cout(t_11606));
compressor_4_2 u2_4060(.a(t_9987), .b(t_10000), .c(t_9997), .d(t_9994), .cin(t_11606), .o(t_11607), .co(t_11608), .cout(t_11609));
compressor_4_2 u2_4061(.a(t_9995), .b(t_10008), .c(t_10005), .d(t_10002), .cin(t_11609), .o(t_11610), .co(t_11611), .cout(t_11612));
compressor_4_2 u2_4062(.a(t_10003), .b(t_10016), .c(t_10013), .d(t_10010), .cin(t_11612), .o(t_11613), .co(t_11614), .cout(t_11615));
compressor_4_2 u2_4063(.a(t_10011), .b(t_10024), .c(t_10021), .d(t_10018), .cin(t_11615), .o(t_11616), .co(t_11617), .cout(t_11618));
compressor_4_2 u2_4064(.a(t_10032), .b(t_10029), .c(t_10026), .d(t_7004), .cin(t_11618), .o(t_11619), .co(t_11620), .cout(t_11621));
half_adder u0_4065(.a(t_10022), .b(t_10019), .o(t_11622), .cout(t_11623));
compressor_4_2 u2_4066(.a(t_10040), .b(t_10037), .c(t_10034), .d(t_11621), .cin(t_11623), .o(t_11624), .co(t_11625), .cout(t_11626));
half_adder u0_4067(.a(t_10030), .b(t_10027), .o(t_11627), .cout(t_11628));
compressor_4_2 u2_4068(.a(t_10048), .b(t_10045), .c(t_10042), .d(t_11626), .cin(t_11628), .o(t_11629), .co(t_11630), .cout(t_11631));
half_adder u0_4069(.a(t_10038), .b(t_10035), .o(t_11632), .cout(t_11633));
compressor_4_2 u2_4070(.a(t_10056), .b(t_10053), .c(t_10050), .d(t_11631), .cin(t_11633), .o(t_11634), .co(t_11635), .cout(t_11636));
half_adder u0_4071(.a(t_10046), .b(t_10043), .o(t_11637), .cout(t_11638));
compressor_4_2 u2_4072(.a(t_10064), .b(t_10061), .c(t_10058), .d(t_11636), .cin(t_11638), .o(t_11639), .co(t_11640), .cout(t_11641));
half_adder u0_4073(.a(t_10054), .b(t_10051), .o(t_11642), .cout(t_11643));
compressor_4_2 u2_4074(.a(t_10069), .b(t_10066), .c(t_7077), .d(t_11641), .cin(t_11643), .o(t_11644), .co(t_11645), .cout(t_11646));
compressor_3_2 u1_4075(.a(t_10062), .b(t_10059), .cin(t_10072), .o(t_11647), .cout(t_11648));
compressor_4_2 u2_4076(.a(t_10077), .b(t_10074), .c(t_7092), .d(t_11646), .cin(t_11648), .o(t_11649), .co(t_11650), .cout(t_11651));
compressor_3_2 u1_4077(.a(t_10070), .b(t_10067), .cin(t_10080), .o(t_11652), .cout(t_11653));
compressor_4_2 u2_4078(.a(t_10085), .b(t_10082), .c(t_7107), .d(t_11651), .cin(t_11653), .o(t_11654), .co(t_11655), .cout(t_11656));
compressor_3_2 u1_4079(.a(t_10078), .b(t_10075), .cin(t_10088), .o(t_11657), .cout(t_11658));
compressor_4_2 u2_4080(.a(t_10093), .b(t_10090), .c(t_7122), .d(t_11656), .cin(t_11658), .o(t_11659), .co(t_11660), .cout(t_11661));
compressor_3_2 u1_4081(.a(t_10086), .b(t_10083), .cin(t_10096), .o(t_11662), .cout(t_11663));
compressor_4_2 u2_4082(.a(t_10101), .b(t_10098), .c(t_7139), .d(t_11661), .cin(t_11663), .o(t_11664), .co(t_11665), .cout(t_11666));
compressor_3_2 u1_4083(.a(t_10094), .b(t_10091), .cin(t_10104), .o(t_11667), .cout(t_11668));
compressor_4_2 u2_4084(.a(t_10112), .b(t_10109), .c(t_10106), .d(t_11666), .cin(t_11668), .o(t_11669), .co(t_11670), .cout(t_11671));
half_adder u0_4085(.a(t_10102), .b(t_10099), .o(t_11672), .cout(t_11673));
compressor_4_2 u2_4086(.a(t_10118), .b(t_10115), .c(t_7173), .d(t_11671), .cin(t_11673), .o(t_11674), .co(t_11675), .cout(t_11676));
compressor_3_2 u1_4087(.a(t_10110), .b(t_10107), .cin(t_10121), .o(t_11677), .cout(t_11678));
compressor_4_2 u2_4088(.a(t_10126), .b(t_10123), .c(t_7190), .d(t_11676), .cin(t_11678), .o(t_11679), .co(t_11680), .cout(t_11681));
compressor_3_2 u1_4089(.a(t_10119), .b(t_10116), .cin(t_10129), .o(t_11682), .cout(t_11683));
compressor_4_2 u2_4090(.a(t_10137), .b(t_10134), .c(t_10131), .d(t_11681), .cin(t_11683), .o(t_11684), .co(t_11685), .cout(t_11686));
half_adder u0_4091(.a(t_10127), .b(t_10124), .o(t_11687), .cout(t_11688));
compressor_4_2 u2_4092(.a(t_10146), .b(t_10143), .c(t_10140), .d(t_11686), .cin(t_11688), .o(t_11689), .co(t_11690), .cout(t_11691));
compressor_3_2 u1_4093(.a(t_10138), .b(t_10135), .cin(t_10132), .o(t_11692), .cout(t_11693));
compressor_4_2 u2_4094(.a(t_10152), .b(t_10149), .c(t_7241), .d(t_11691), .cin(t_11693), .o(t_11694), .co(t_11695), .cout(t_11696));
compressor_3_2 u1_4095(.a(t_10144), .b(t_10141), .cin(t_10155), .o(t_11697), .cout(t_11698));
compressor_4_2 u2_4096(.a(t_10160), .b(t_10157), .c(t_7261), .d(t_11696), .cin(t_11698), .o(t_11699), .co(t_11700), .cout(t_11701));
compressor_3_2 u1_4097(.a(t_10153), .b(t_10150), .cin(t_10163), .o(t_11702), .cout(t_11703));
compressor_4_2 u2_4098(.a(t_10172), .b(t_10169), .c(t_10166), .d(t_11701), .cin(t_11703), .o(t_11704), .co(t_11705), .cout(t_11706));
compressor_3_2 u1_4099(.a(t_10164), .b(t_10161), .cin(t_10158), .o(t_11707), .cout(t_11708));
compressor_4_2 u2_4100(.a(t_10181), .b(t_10178), .c(t_10175), .d(t_11706), .cin(t_11708), .o(t_11709), .co(t_11710), .cout(t_11711));
compressor_3_2 u1_4101(.a(t_10173), .b(t_10170), .cin(t_10167), .o(t_11712), .cout(t_11713));
compressor_4_2 u2_4102(.a(t_10190), .b(t_10187), .c(t_10184), .d(t_11711), .cin(t_11713), .o(t_11714), .co(t_11715), .cout(t_11716));
compressor_3_2 u1_4103(.a(t_10182), .b(t_10179), .cin(t_10176), .o(t_11717), .cout(t_11718));
compressor_4_2 u2_4104(.a(t_10199), .b(t_10196), .c(t_10193), .d(t_11716), .cin(t_11718), .o(t_11719), .co(t_11720), .cout(t_11721));
compressor_3_2 u1_4105(.a(t_10191), .b(t_10188), .cin(t_10185), .o(t_11722), .cout(t_11723));
compressor_4_2 u2_4106(.a(t_10205), .b(t_10202), .c(t_7349), .d(t_11721), .cin(t_11723), .o(t_11724), .co(t_11725), .cout(t_11726));
compressor_3_2 u1_4107(.a(t_10197), .b(t_10194), .cin(t_10208), .o(t_11727), .cout(t_11728));
compressor_4_2 u2_4108(.a(t_10214), .b(t_10211), .c(t_7367), .d(t_11726), .cin(t_11728), .o(t_11729), .co(t_11730), .cout(t_11731));
compressor_3_2 u1_4109(.a(t_10206), .b(t_10203), .cin(t_10217), .o(t_11732), .cout(t_11733));
compressor_4_2 u2_4110(.a(t_10223), .b(t_10220), .c(t_7385), .d(t_11731), .cin(t_11733), .o(t_11734), .co(t_11735), .cout(t_11736));
compressor_3_2 u1_4111(.a(t_10215), .b(t_10212), .cin(t_10226), .o(t_11737), .cout(t_11738));
compressor_4_2 u2_4112(.a(t_10232), .b(t_10229), .c(t_7403), .d(t_11736), .cin(t_11738), .o(t_11739), .co(t_11740), .cout(t_11741));
compressor_3_2 u1_4113(.a(t_10224), .b(t_10221), .cin(t_10235), .o(t_11742), .cout(t_11743));
compressor_4_2 u2_4114(.a(t_10241), .b(t_10238), .c(t_7423), .d(t_11741), .cin(t_11743), .o(t_11744), .co(t_11745), .cout(t_11746));
compressor_3_2 u1_4115(.a(t_10233), .b(t_10230), .cin(t_10244), .o(t_11747), .cout(t_11748));
compressor_4_2 u2_4116(.a(t_10253), .b(t_10250), .c(t_10247), .d(t_11746), .cin(t_11748), .o(t_11749), .co(t_11750), .cout(t_11751));
compressor_3_2 u1_4117(.a(t_10242), .b(t_10239), .cin(t_10256), .o(t_11752), .cout(t_11753));
compressor_4_2 u2_4118(.a(t_10264), .b(t_10261), .c(t_10258), .d(t_11751), .cin(t_11753), .o(t_11754), .co(t_11755), .cout(t_11756));
compressor_3_2 u1_4119(.a(t_10251), .b(t_10248), .cin(t_10267), .o(t_11757), .cout(t_11758));
compressor_4_2 u2_4120(.a(t_10275), .b(t_10272), .c(t_10269), .d(t_11756), .cin(t_11758), .o(t_11759), .co(t_11760), .cout(t_11761));
compressor_3_2 u1_4121(.a(t_10262), .b(t_10259), .cin(t_10278), .o(t_11762), .cout(t_11763));
compressor_4_2 u2_4122(.a(t_10286), .b(t_10283), .c(t_10280), .d(t_11761), .cin(t_11763), .o(t_11764), .co(t_11765), .cout(t_11766));
compressor_3_2 u1_4123(.a(t_10273), .b(t_10270), .cin(t_10289), .o(t_11767), .cout(t_11768));
compressor_4_2 u2_4124(.a(t_10297), .b(t_10294), .c(t_10291), .d(t_11766), .cin(t_11768), .o(t_11769), .co(t_11770), .cout(t_11771));
compressor_3_2 u1_4125(.a(t_10284), .b(t_10281), .cin(t_10300), .o(t_11772), .cout(t_11773));
compressor_4_2 u2_4126(.a(t_10308), .b(t_10305), .c(t_10302), .d(t_11771), .cin(t_11773), .o(t_11774), .co(t_11775), .cout(t_11776));
compressor_3_2 u1_4127(.a(t_10295), .b(t_10292), .cin(t_10311), .o(t_11777), .cout(t_11778));
compressor_4_2 u2_4128(.a(t_10316), .b(t_10313), .c(t_7566), .d(t_11776), .cin(t_11778), .o(t_11779), .co(t_11780), .cout(t_11781));
compressor_4_2 u2_4129(.a(t_10309), .b(t_10306), .c(t_10303), .d(t_10322), .cin(t_10319), .o(t_11782), .co(t_11783), .cout(t_11784));
compressor_4_2 u2_4130(.a(t_10330), .b(t_10327), .c(t_10324), .d(t_11781), .cin(t_11784), .o(t_11785), .co(t_11786), .cout(t_11787));
compressor_3_2 u1_4131(.a(t_10317), .b(t_10314), .cin(t_10333), .o(t_11788), .cout(t_11789));
compressor_4_2 u2_4132(.a(t_10341), .b(t_10338), .c(t_10335), .d(t_11787), .cin(t_11789), .o(t_11790), .co(t_11791), .cout(t_11792));
compressor_3_2 u1_4133(.a(t_10328), .b(t_10325), .cin(t_10344), .o(t_11793), .cout(t_11794));
compressor_4_2 u2_4134(.a(t_10352), .b(t_10349), .c(t_10346), .d(t_11792), .cin(t_11794), .o(t_11795), .co(t_11796), .cout(t_11797));
compressor_3_2 u1_4135(.a(t_10339), .b(t_10336), .cin(t_10355), .o(t_11798), .cout(t_11799));
compressor_4_2 u2_4136(.a(t_10363), .b(t_10360), .c(t_10357), .d(t_11797), .cin(t_11799), .o(t_11800), .co(t_11801), .cout(t_11802));
compressor_3_2 u1_4137(.a(t_10350), .b(t_10347), .cin(t_10366), .o(t_11803), .cout(t_11804));
compressor_4_2 u2_4138(.a(t_10371), .b(t_10368), .c(t_7669), .d(t_11802), .cin(t_11804), .o(t_11805), .co(t_11806), .cout(t_11807));
compressor_4_2 u2_4139(.a(t_10364), .b(t_10361), .c(t_10358), .d(t_10377), .cin(t_10374), .o(t_11808), .co(t_11809), .cout(t_11810));
compressor_4_2 u2_4140(.a(t_10382), .b(t_10379), .c(t_7690), .d(t_11807), .cin(t_11810), .o(t_11811), .co(t_11812), .cout(t_11813));
compressor_4_2 u2_4141(.a(t_10375), .b(t_10372), .c(t_10369), .d(t_10388), .cin(t_10385), .o(t_11814), .co(t_11815), .cout(t_11816));
compressor_4_2 u2_4142(.a(t_10393), .b(t_10390), .c(t_7711), .d(t_11813), .cin(t_11816), .o(t_11817), .co(t_11818), .cout(t_11819));
compressor_4_2 u2_4143(.a(t_10386), .b(t_10383), .c(t_10380), .d(t_10399), .cin(t_10396), .o(t_11820), .co(t_11821), .cout(t_11822));
compressor_4_2 u2_4144(.a(t_10404), .b(t_10401), .c(t_7732), .d(t_11819), .cin(t_11822), .o(t_11823), .co(t_11824), .cout(t_11825));
compressor_4_2 u2_4145(.a(t_10397), .b(t_10394), .c(t_10391), .d(t_10410), .cin(t_10407), .o(t_11826), .co(t_11827), .cout(t_11828));
compressor_4_2 u2_4146(.a(t_10415), .b(t_10412), .c(t_7755), .d(t_11825), .cin(t_11828), .o(t_11829), .co(t_11830), .cout(t_11831));
compressor_4_2 u2_4147(.a(t_10408), .b(t_10405), .c(t_10402), .d(t_10421), .cin(t_10418), .o(t_11832), .co(t_11833), .cout(t_11834));
compressor_4_2 u2_4148(.a(t_10429), .b(t_10426), .c(t_10423), .d(t_11831), .cin(t_11834), .o(t_11835), .co(t_11836), .cout(t_11837));
compressor_3_2 u1_4149(.a(t_10416), .b(t_10413), .cin(t_10432), .o(t_11838), .cout(t_11839));
compressor_4_2 u2_4150(.a(t_10438), .b(t_10435), .c(t_7801), .d(t_11837), .cin(t_11839), .o(t_11840), .co(t_11841), .cout(t_11842));
compressor_4_2 u2_4151(.a(t_10430), .b(t_10427), .c(t_10424), .d(t_10444), .cin(t_10441), .o(t_11843), .co(t_11844), .cout(t_11845));
compressor_4_2 u2_4152(.a(t_10449), .b(t_10446), .c(t_7824), .d(t_11842), .cin(t_11845), .o(t_11846), .co(t_11847), .cout(t_11848));
compressor_4_2 u2_4153(.a(t_10442), .b(t_10439), .c(t_10436), .d(t_10455), .cin(t_10452), .o(t_11849), .co(t_11850), .cout(t_11851));
compressor_4_2 u2_4154(.a(t_10463), .b(t_10460), .c(t_10457), .d(t_11848), .cin(t_11851), .o(t_11852), .co(t_11853), .cout(t_11854));
compressor_3_2 u1_4155(.a(t_10450), .b(t_10447), .cin(t_10466), .o(t_11855), .cout(t_11856));
compressor_4_2 u2_4156(.a(t_10475), .b(t_10472), .c(t_10469), .d(t_11854), .cin(t_11856), .o(t_11857), .co(t_11858), .cout(t_11859));
compressor_4_2 u2_4157(.a(t_10467), .b(t_10464), .c(t_10461), .d(t_10458), .cin(t_10478), .o(t_11860), .co(t_11861), .cout(t_11862));
compressor_4_2 u2_4158(.a(t_10484), .b(t_10481), .c(t_7893), .d(t_11859), .cin(t_11862), .o(t_11863), .co(t_11864), .cout(t_11865));
compressor_4_2 u2_4159(.a(t_10476), .b(t_10473), .c(t_10470), .d(t_10490), .cin(t_10487), .o(t_11866), .co(t_11867), .cout(t_11868));
compressor_4_2 u2_4160(.a(t_10495), .b(t_10492), .c(t_7919), .d(t_11865), .cin(t_11868), .o(t_11869), .co(t_11870), .cout(t_11871));
compressor_4_2 u2_4161(.a(t_10488), .b(t_10485), .c(t_10482), .d(t_10501), .cin(t_10498), .o(t_11872), .co(t_11873), .cout(t_11874));
compressor_4_2 u2_4162(.a(t_10510), .b(t_10507), .c(t_10504), .d(t_11871), .cin(t_11874), .o(t_11875), .co(t_11876), .cout(t_11877));
compressor_4_2 u2_4163(.a(t_10502), .b(t_10499), .c(t_10496), .d(t_10493), .cin(t_10513), .o(t_11878), .co(t_11879), .cout(t_11880));
compressor_4_2 u2_4164(.a(t_10522), .b(t_10519), .c(t_10516), .d(t_11877), .cin(t_11880), .o(t_11881), .co(t_11882), .cout(t_11883));
compressor_4_2 u2_4165(.a(t_10514), .b(t_10511), .c(t_10508), .d(t_10505), .cin(t_10525), .o(t_11884), .co(t_11885), .cout(t_11886));
compressor_4_2 u2_4166(.a(t_10534), .b(t_10531), .c(t_10528), .d(t_11883), .cin(t_11886), .o(t_11887), .co(t_11888), .cout(t_11889));
compressor_4_2 u2_4167(.a(t_10526), .b(t_10523), .c(t_10520), .d(t_10517), .cin(t_10537), .o(t_11890), .co(t_11891), .cout(t_11892));
compressor_4_2 u2_4168(.a(t_10546), .b(t_10543), .c(t_10540), .d(t_11889), .cin(t_11892), .o(t_11893), .co(t_11894), .cout(t_11895));
compressor_4_2 u2_4169(.a(t_10538), .b(t_10535), .c(t_10532), .d(t_10529), .cin(t_10549), .o(t_11896), .co(t_11897), .cout(t_11898));
compressor_4_2 u2_4170(.a(t_10555), .b(t_10552), .c(t_8037), .d(t_11895), .cin(t_11898), .o(t_11899), .co(t_11900), .cout(t_11901));
compressor_4_2 u2_4171(.a(t_10547), .b(t_10544), .c(t_10541), .d(t_10561), .cin(t_10558), .o(t_11902), .co(t_11903), .cout(t_11904));
compressor_4_2 u2_4172(.a(t_10567), .b(t_10564), .c(t_8061), .d(t_11901), .cin(t_11904), .o(t_11905), .co(t_11906), .cout(t_11907));
compressor_4_2 u2_4173(.a(t_10559), .b(t_10556), .c(t_10553), .d(t_10573), .cin(t_10570), .o(t_11908), .co(t_11909), .cout(t_11910));
compressor_4_2 u2_4174(.a(t_10582), .b(t_10579), .c(t_10576), .d(t_11907), .cin(t_11910), .o(t_11911), .co(t_11912), .cout(t_11913));
compressor_4_2 u2_4175(.a(t_10574), .b(t_10571), .c(t_10568), .d(t_10565), .cin(t_10585), .o(t_11914), .co(t_11915), .cout(t_11916));
compressor_4_2 u2_4176(.a(t_10594), .b(t_10591), .c(t_10588), .d(t_11913), .cin(t_11916), .o(t_11917), .co(t_11918), .cout(t_11919));
compressor_4_2 u2_4177(.a(t_10586), .b(t_10583), .c(t_10580), .d(t_10577), .cin(t_10597), .o(t_11920), .co(t_11921), .cout(t_11922));
compressor_4_2 u2_4178(.a(t_10603), .b(t_10600), .c(t_8133), .d(t_11919), .cin(t_11922), .o(t_11923), .co(t_11924), .cout(t_11925));
compressor_4_2 u2_4179(.a(t_10595), .b(t_10592), .c(t_10589), .d(t_10609), .cin(t_10606), .o(t_11926), .co(t_11927), .cout(t_11928));
compressor_4_2 u2_4180(.a(t_10618), .b(t_10615), .c(t_10612), .d(t_11925), .cin(t_11928), .o(t_11929), .co(t_11930), .cout(t_11931));
compressor_4_2 u2_4181(.a(t_10610), .b(t_10607), .c(t_10604), .d(t_10601), .cin(t_10621), .o(t_11932), .co(t_11933), .cout(t_11934));
compressor_4_2 u2_4182(.a(t_10627), .b(t_10624), .c(t_8181), .d(t_11931), .cin(t_11934), .o(t_11935), .co(t_11936), .cout(t_11937));
compressor_4_2 u2_4183(.a(t_10619), .b(t_10616), .c(t_10613), .d(t_10633), .cin(t_10630), .o(t_11938), .co(t_11939), .cout(t_11940));
compressor_4_2 u2_4184(.a(t_10642), .b(t_10639), .c(t_10636), .d(t_11937), .cin(t_11940), .o(t_11941), .co(t_11942), .cout(t_11943));
compressor_4_2 u2_4185(.a(t_10634), .b(t_10631), .c(t_10628), .d(t_10625), .cin(t_10645), .o(t_11944), .co(t_11945), .cout(t_11946));
compressor_4_2 u2_4186(.a(t_10654), .b(t_10651), .c(t_10648), .d(t_11943), .cin(t_11946), .o(t_11947), .co(t_11948), .cout(t_11949));
compressor_4_2 u2_4187(.a(t_10646), .b(t_10643), .c(t_10640), .d(t_10637), .cin(t_10657), .o(t_11950), .co(t_11951), .cout(t_11952));
compressor_4_2 u2_4188(.a(t_10666), .b(t_10663), .c(t_10660), .d(t_11949), .cin(t_11952), .o(t_11953), .co(t_11954), .cout(t_11955));
compressor_4_2 u2_4189(.a(t_10658), .b(t_10655), .c(t_10652), .d(t_10649), .cin(t_10669), .o(t_11956), .co(t_11957), .cout(t_11958));
compressor_4_2 u2_4190(.a(t_10678), .b(t_10675), .c(t_10672), .d(t_11955), .cin(t_11958), .o(t_11959), .co(t_11960), .cout(t_11961));
compressor_4_2 u2_4191(.a(t_10670), .b(t_10667), .c(t_10664), .d(t_10661), .cin(t_10681), .o(t_11962), .co(t_11963), .cout(t_11964));
compressor_4_2 u2_4192(.a(t_10687), .b(t_10684), .c(t_8294), .d(t_11961), .cin(t_11964), .o(t_11965), .co(t_11966), .cout(t_11967));
compressor_4_2 u2_4193(.a(t_10679), .b(t_10676), .c(t_10673), .d(t_10693), .cin(t_10690), .o(t_11968), .co(t_11969), .cout(t_11970));
compressor_4_2 u2_4194(.a(t_10701), .b(t_10698), .c(t_10695), .d(t_11967), .cin(t_11970), .o(t_11971), .co(t_11972), .cout(t_11973));
compressor_3_2 u1_4195(.a(t_10688), .b(t_10685), .cin(t_10704), .o(t_11974), .cout(t_11975));
compressor_4_2 u2_4196(.a(t_10710), .b(t_10707), .c(t_8340), .d(t_11973), .cin(t_11975), .o(t_11976), .co(t_11977), .cout(t_11978));
compressor_4_2 u2_4197(.a(t_10702), .b(t_10699), .c(t_10696), .d(t_10716), .cin(t_10713), .o(t_11979), .co(t_11980), .cout(t_11981));
compressor_4_2 u2_4198(.a(t_10721), .b(t_10718), .c(t_8363), .d(t_11978), .cin(t_11981), .o(t_11982), .co(t_11983), .cout(t_11984));
compressor_4_2 u2_4199(.a(t_10714), .b(t_10711), .c(t_10708), .d(t_10727), .cin(t_10724), .o(t_11985), .co(t_11986), .cout(t_11987));
compressor_4_2 u2_4200(.a(t_10732), .b(t_10729), .c(t_8386), .d(t_11984), .cin(t_11987), .o(t_11988), .co(t_11989), .cout(t_11990));
compressor_4_2 u2_4201(.a(t_10725), .b(t_10722), .c(t_10719), .d(t_10738), .cin(t_10735), .o(t_11991), .co(t_11992), .cout(t_11993));
compressor_4_2 u2_4202(.a(t_10743), .b(t_10740), .c(t_8409), .d(t_11990), .cin(t_11993), .o(t_11994), .co(t_11995), .cout(t_11996));
compressor_4_2 u2_4203(.a(t_10736), .b(t_10733), .c(t_10730), .d(t_10749), .cin(t_10746), .o(t_11997), .co(t_11998), .cout(t_11999));
compressor_4_2 u2_4204(.a(t_10754), .b(t_10751), .c(t_8432), .d(t_11996), .cin(t_11999), .o(t_12000), .co(t_12001), .cout(t_12002));
compressor_4_2 u2_4205(.a(t_10747), .b(t_10744), .c(t_10741), .d(t_10760), .cin(t_10757), .o(t_12003), .co(t_12004), .cout(t_12005));
compressor_4_2 u2_4206(.a(t_10765), .b(t_10762), .c(t_8455), .d(t_12002), .cin(t_12005), .o(t_12006), .co(t_12007), .cout(t_12008));
compressor_4_2 u2_4207(.a(t_10758), .b(t_10755), .c(t_10752), .d(t_10771), .cin(t_10768), .o(t_12009), .co(t_12010), .cout(t_12011));
compressor_4_2 u2_4208(.a(t_10776), .b(t_10773), .c(t_8478), .d(t_12008), .cin(t_12011), .o(t_12012), .co(t_12013), .cout(t_12014));
compressor_4_2 u2_4209(.a(t_10769), .b(t_10766), .c(t_10763), .d(t_10782), .cin(t_10779), .o(t_12015), .co(t_12016), .cout(t_12017));
compressor_4_2 u2_4210(.a(t_10787), .b(t_10784), .c(t_8501), .d(t_12014), .cin(t_12017), .o(t_12018), .co(t_12019), .cout(t_12020));
compressor_4_2 u2_4211(.a(t_10780), .b(t_10777), .c(t_10774), .d(t_10793), .cin(t_10790), .o(t_12021), .co(t_12022), .cout(t_12023));
compressor_4_2 u2_4212(.a(t_10801), .b(t_10798), .c(t_10795), .d(t_12020), .cin(t_12023), .o(t_12024), .co(t_12025), .cout(t_12026));
compressor_3_2 u1_4213(.a(t_10788), .b(t_10785), .cin(t_10804), .o(t_12027), .cout(t_12028));
compressor_4_2 u2_4214(.a(t_10809), .b(t_10806), .c(t_8543), .d(t_12026), .cin(t_12028), .o(t_12029), .co(t_12030), .cout(t_12031));
compressor_4_2 u2_4215(.a(t_10802), .b(t_10799), .c(t_10796), .d(t_10815), .cin(t_10812), .o(t_12032), .co(t_12033), .cout(t_12034));
compressor_4_2 u2_4216(.a(t_10823), .b(t_10820), .c(t_10817), .d(t_12031), .cin(t_12034), .o(t_12035), .co(t_12036), .cout(t_12037));
compressor_3_2 u1_4217(.a(t_10810), .b(t_10807), .cin(t_10826), .o(t_12038), .cout(t_12039));
compressor_4_2 u2_4218(.a(t_10834), .b(t_10831), .c(t_10828), .d(t_12037), .cin(t_12039), .o(t_12040), .co(t_12041), .cout(t_12042));
compressor_3_2 u1_4219(.a(t_10821), .b(t_10818), .cin(t_10837), .o(t_12043), .cout(t_12044));
compressor_4_2 u2_4220(.a(t_10845), .b(t_10842), .c(t_10839), .d(t_12042), .cin(t_12044), .o(t_12045), .co(t_12046), .cout(t_12047));
compressor_3_2 u1_4221(.a(t_10832), .b(t_10829), .cin(t_10848), .o(t_12048), .cout(t_12049));
compressor_4_2 u2_4222(.a(t_10856), .b(t_10853), .c(t_10850), .d(t_12047), .cin(t_12049), .o(t_12050), .co(t_12051), .cout(t_12052));
compressor_3_2 u1_4223(.a(t_10843), .b(t_10840), .cin(t_10859), .o(t_12053), .cout(t_12054));
compressor_4_2 u2_4224(.a(t_10867), .b(t_10864), .c(t_10861), .d(t_12052), .cin(t_12054), .o(t_12055), .co(t_12056), .cout(t_12057));
compressor_3_2 u1_4225(.a(t_10854), .b(t_10851), .cin(t_10870), .o(t_12058), .cout(t_12059));
compressor_4_2 u2_4226(.a(t_10878), .b(t_10875), .c(t_10872), .d(t_12057), .cin(t_12059), .o(t_12060), .co(t_12061), .cout(t_12062));
compressor_3_2 u1_4227(.a(t_10865), .b(t_10862), .cin(t_10881), .o(t_12063), .cout(t_12064));
compressor_4_2 u2_4228(.a(t_10889), .b(t_10886), .c(t_10883), .d(t_12062), .cin(t_12064), .o(t_12065), .co(t_12066), .cout(t_12067));
compressor_3_2 u1_4229(.a(t_10876), .b(t_10873), .cin(t_10892), .o(t_12068), .cout(t_12069));
compressor_4_2 u2_4230(.a(t_10900), .b(t_10897), .c(t_10894), .d(t_12067), .cin(t_12069), .o(t_12070), .co(t_12071), .cout(t_12072));
compressor_3_2 u1_4231(.a(t_10887), .b(t_10884), .cin(t_10903), .o(t_12073), .cout(t_12074));
compressor_4_2 u2_4232(.a(t_10911), .b(t_10908), .c(t_10905), .d(t_12072), .cin(t_12074), .o(t_12075), .co(t_12076), .cout(t_12077));
compressor_3_2 u1_4233(.a(t_10898), .b(t_10895), .cin(t_10914), .o(t_12078), .cout(t_12079));
compressor_4_2 u2_4234(.a(t_10922), .b(t_10919), .c(t_10916), .d(t_12077), .cin(t_12079), .o(t_12080), .co(t_12081), .cout(t_12082));
compressor_3_2 u1_4235(.a(t_10909), .b(t_10906), .cin(t_10925), .o(t_12083), .cout(t_12084));
compressor_4_2 u2_4236(.a(t_10933), .b(t_10930), .c(t_10927), .d(t_12082), .cin(t_12084), .o(t_12085), .co(t_12086), .cout(t_12087));
compressor_3_2 u1_4237(.a(t_10920), .b(t_10917), .cin(t_10936), .o(t_12088), .cout(t_12089));
compressor_4_2 u2_4238(.a(t_10944), .b(t_10941), .c(t_10938), .d(t_12087), .cin(t_12089), .o(t_12090), .co(t_12091), .cout(t_12092));
compressor_3_2 u1_4239(.a(t_10931), .b(t_10928), .cin(t_10947), .o(t_12093), .cout(t_12094));
compressor_4_2 u2_4240(.a(t_10955), .b(t_10952), .c(t_10949), .d(t_12092), .cin(t_12094), .o(t_12095), .co(t_12096), .cout(t_12097));
compressor_3_2 u1_4241(.a(t_10942), .b(t_10939), .cin(t_10958), .o(t_12098), .cout(t_12099));
compressor_4_2 u2_4242(.a(t_10966), .b(t_10963), .c(t_10960), .d(t_12097), .cin(t_12099), .o(t_12100), .co(t_12101), .cout(t_12102));
compressor_3_2 u1_4243(.a(t_10953), .b(t_10950), .cin(t_10969), .o(t_12103), .cout(t_12104));
compressor_4_2 u2_4244(.a(t_10974), .b(t_10971), .c(t_8839), .d(t_12102), .cin(t_12104), .o(t_12105), .co(t_12106), .cout(t_12107));
compressor_3_2 u1_4245(.a(t_10964), .b(t_10961), .cin(t_10977), .o(t_12108), .cout(t_12109));
compressor_4_2 u2_4246(.a(t_10983), .b(t_10980), .c(t_8857), .d(t_12107), .cin(t_12109), .o(t_12110), .co(t_12111), .cout(t_12112));
compressor_3_2 u1_4247(.a(t_10975), .b(t_10972), .cin(t_10986), .o(t_12113), .cout(t_12114));
compressor_4_2 u2_4248(.a(t_10995), .b(t_10992), .c(t_10989), .d(t_12112), .cin(t_12114), .o(t_12115), .co(t_12116), .cout(t_12117));
compressor_3_2 u1_4249(.a(t_10987), .b(t_10984), .cin(t_10981), .o(t_12118), .cout(t_12119));
compressor_4_2 u2_4250(.a(t_11004), .b(t_11001), .c(t_10998), .d(t_12117), .cin(t_12119), .o(t_12120), .co(t_12121), .cout(t_12122));
compressor_3_2 u1_4251(.a(t_10996), .b(t_10993), .cin(t_10990), .o(t_12123), .cout(t_12124));
compressor_4_2 u2_4252(.a(t_11013), .b(t_11010), .c(t_11007), .d(t_12122), .cin(t_12124), .o(t_12125), .co(t_12126), .cout(t_12127));
compressor_3_2 u1_4253(.a(t_11005), .b(t_11002), .cin(t_10999), .o(t_12128), .cout(t_12129));
compressor_4_2 u2_4254(.a(t_11022), .b(t_11019), .c(t_11016), .d(t_12127), .cin(t_12129), .o(t_12130), .co(t_12131), .cout(t_12132));
compressor_3_2 u1_4255(.a(t_11014), .b(t_11011), .cin(t_11008), .o(t_12133), .cout(t_12134));
compressor_4_2 u2_4256(.a(t_11028), .b(t_11025), .c(t_8940), .d(t_12132), .cin(t_12134), .o(t_12135), .co(t_12136), .cout(t_12137));
compressor_3_2 u1_4257(.a(t_11020), .b(t_11017), .cin(t_11031), .o(t_12138), .cout(t_12139));
compressor_4_2 u2_4258(.a(t_11039), .b(t_11036), .c(t_11033), .d(t_12137), .cin(t_12139), .o(t_12140), .co(t_12141), .cout(t_12142));
half_adder u0_4259(.a(t_11029), .b(t_11026), .o(t_12143), .cout(t_12144));
compressor_4_2 u2_4260(.a(t_11045), .b(t_11042), .c(t_8974), .d(t_12142), .cin(t_12144), .o(t_12145), .co(t_12146), .cout(t_12147));
compressor_3_2 u1_4261(.a(t_11037), .b(t_11034), .cin(t_11048), .o(t_12148), .cout(t_12149));
compressor_4_2 u2_4262(.a(t_11053), .b(t_11050), .c(t_8991), .d(t_12147), .cin(t_12149), .o(t_12150), .co(t_12151), .cout(t_12152));
compressor_3_2 u1_4263(.a(t_11046), .b(t_11043), .cin(t_11056), .o(t_12153), .cout(t_12154));
compressor_4_2 u2_4264(.a(t_11061), .b(t_11058), .c(t_9008), .d(t_12152), .cin(t_12154), .o(t_12155), .co(t_12156), .cout(t_12157));
compressor_3_2 u1_4265(.a(t_11054), .b(t_11051), .cin(t_11064), .o(t_12158), .cout(t_12159));
compressor_4_2 u2_4266(.a(t_11069), .b(t_11066), .c(t_9025), .d(t_12157), .cin(t_12159), .o(t_12160), .co(t_12161), .cout(t_12162));
compressor_3_2 u1_4267(.a(t_11062), .b(t_11059), .cin(t_11072), .o(t_12163), .cout(t_12164));
compressor_4_2 u2_4268(.a(t_11077), .b(t_11074), .c(t_9042), .d(t_12162), .cin(t_12164), .o(t_12165), .co(t_12166), .cout(t_12167));
compressor_3_2 u1_4269(.a(t_11070), .b(t_11067), .cin(t_11080), .o(t_12168), .cout(t_12169));
compressor_4_2 u2_4270(.a(t_11085), .b(t_11082), .c(t_9059), .d(t_12167), .cin(t_12169), .o(t_12170), .co(t_12171), .cout(t_12172));
compressor_3_2 u1_4271(.a(t_11078), .b(t_11075), .cin(t_11088), .o(t_12173), .cout(t_12174));
compressor_4_2 u2_4272(.a(t_11093), .b(t_11090), .c(t_9076), .d(t_12172), .cin(t_12174), .o(t_12175), .co(t_12176), .cout(t_12177));
compressor_3_2 u1_4273(.a(t_11086), .b(t_11083), .cin(t_11096), .o(t_12178), .cout(t_12179));
compressor_4_2 u2_4274(.a(t_11101), .b(t_11098), .c(t_9093), .d(t_12177), .cin(t_12179), .o(t_12180), .co(t_12181), .cout(t_12182));
compressor_3_2 u1_4275(.a(t_11094), .b(t_11091), .cin(t_11104), .o(t_12183), .cout(t_12184));
compressor_4_2 u2_4276(.a(t_11112), .b(t_11109), .c(t_11106), .d(t_12182), .cin(t_12184), .o(t_12185), .co(t_12186), .cout(t_12187));
half_adder u0_4277(.a(t_11102), .b(t_11099), .o(t_12188), .cout(t_12189));
compressor_4_2 u2_4278(.a(t_11117), .b(t_11114), .c(t_9123), .d(t_12187), .cin(t_12189), .o(t_12190), .co(t_12191), .cout(t_12192));
compressor_3_2 u1_4279(.a(t_11110), .b(t_11107), .cin(t_11120), .o(t_12193), .cout(t_12194));
compressor_4_2 u2_4280(.a(t_11128), .b(t_11125), .c(t_11122), .d(t_12192), .cin(t_12194), .o(t_12195), .co(t_12196), .cout(t_12197));
half_adder u0_4281(.a(t_11118), .b(t_11115), .o(t_12198), .cout(t_12199));
compressor_4_2 u2_4282(.a(t_11136), .b(t_11133), .c(t_11130), .d(t_12197), .cin(t_12199), .o(t_12200), .co(t_12201), .cout(t_12202));
half_adder u0_4283(.a(t_11126), .b(t_11123), .o(t_12203), .cout(t_12204));
compressor_4_2 u2_4284(.a(t_11144), .b(t_11141), .c(t_11138), .d(t_12202), .cin(t_12204), .o(t_12205), .co(t_12206), .cout(t_12207));
half_adder u0_4285(.a(t_11134), .b(t_11131), .o(t_12208), .cout(t_12209));
compressor_4_2 u2_4286(.a(t_11152), .b(t_11149), .c(t_11146), .d(t_12207), .cin(t_12209), .o(t_12210), .co(t_12211), .cout(t_12212));
half_adder u0_4287(.a(t_11142), .b(t_11139), .o(t_12213), .cout(t_12214));
compressor_4_2 u2_4288(.a(t_11160), .b(t_11157), .c(t_11154), .d(t_12212), .cin(t_12214), .o(t_12215), .co(t_12216), .cout(t_12217));
half_adder u0_4289(.a(t_11150), .b(t_11147), .o(t_12218), .cout(t_12219));
compressor_4_2 u2_4290(.a(t_11168), .b(t_11165), .c(t_11162), .d(t_12217), .cin(t_12219), .o(t_12220), .co(t_12221), .cout(t_12222));
half_adder u0_4291(.a(t_11158), .b(t_11155), .o(t_12223), .cout(t_12224));
compressor_4_2 u2_4292(.a(t_11176), .b(t_11173), .c(t_11170), .d(t_12222), .cin(t_12224), .o(t_12225), .co(t_12226), .cout(t_12227));
half_adder u0_4293(.a(t_11166), .b(t_11163), .o(t_12228), .cout(t_12229));
compressor_4_2 u2_4294(.a(t_11184), .b(t_11181), .c(t_11178), .d(t_12227), .cin(t_12229), .o(t_12230), .co(t_12231), .cout(t_12232));
half_adder u0_4295(.a(t_11174), .b(t_11171), .o(t_12233), .cout(t_12234));
compressor_4_2 u2_4296(.a(t_11192), .b(t_11189), .c(t_11186), .d(t_12232), .cin(t_12234), .o(t_12235), .co(t_12236), .cout(t_12237));
half_adder u0_4297(.a(t_11182), .b(t_11179), .o(t_12238), .cout(t_12239));
compressor_4_2 u2_4298(.a(t_11200), .b(t_11197), .c(t_11194), .d(t_12237), .cin(t_12239), .o(t_12240), .co(t_12241), .cout(t_12242));
half_adder u0_4299(.a(t_11190), .b(t_11187), .o(t_12243), .cout(t_12244));
compressor_4_2 u2_4300(.a(t_11208), .b(t_11205), .c(t_11202), .d(t_12242), .cin(t_12244), .o(t_12245), .co(t_12246), .cout(t_12247));
half_adder u0_4301(.a(t_11198), .b(t_11195), .o(t_12248), .cout(t_12249));
compressor_4_2 u2_4302(.a(t_11216), .b(t_11213), .c(t_11210), .d(t_12247), .cin(t_12249), .o(t_12250), .co(t_12251), .cout(t_12252));
half_adder u0_4303(.a(t_11206), .b(t_11203), .o(t_12253), .cout(t_12254));
compressor_4_2 u2_4304(.a(t_11224), .b(t_11221), .c(t_11218), .d(t_12252), .cin(t_12254), .o(t_12255), .co(t_12256), .cout(t_12257));
half_adder u0_4305(.a(t_11214), .b(t_11211), .o(t_12258), .cout(t_12259));
compressor_4_2 u2_4306(.a(t_11232), .b(t_11229), .c(t_11226), .d(t_12257), .cin(t_12259), .o(t_12260), .co(t_12261), .cout(t_12262));
half_adder u0_4307(.a(t_11222), .b(t_11219), .o(t_12263), .cout(t_12264));
compressor_4_2 u2_4308(.a(t_11237), .b(t_11234), .c(t_9329), .d(t_12262), .cin(t_12264), .o(t_12265), .co(t_12266), .cout(t_12267));
half_adder u0_4309(.a(t_11230), .b(t_11227), .o(t_12268), .cout(t_12269));
compressor_4_2 u2_4310(.a(t_11243), .b(t_11240), .c(t_9341), .d(t_12267), .cin(t_12269), .o(t_12270), .co(t_12271), .cout(t_12272));
half_adder u0_4311(.a(t_11238), .b(t_11235), .o(t_12273), .cout(t_12274));
compressor_4_2 u2_4312(.a(t_11241), .b(t_11249), .c(t_11246), .d(t_12272), .cin(t_12274), .o(t_12275), .co(t_12276), .cout(t_12277));
compressor_4_2 u2_4313(.a(t_11250), .b(t_11247), .c(t_11255), .d(t_11252), .cin(t_12277), .o(t_12278), .co(t_12279), .cout(t_12280));
compressor_4_2 u2_4314(.a(t_11256), .b(t_11253), .c(t_11261), .d(t_11258), .cin(t_12280), .o(t_12281), .co(t_12282), .cout(t_12283));
compressor_4_2 u2_4315(.a(t_11262), .b(t_11259), .c(t_11267), .d(t_11264), .cin(t_12283), .o(t_12284), .co(t_12285), .cout(t_12286));
compressor_4_2 u2_4316(.a(t_11265), .b(t_11273), .c(t_11270), .d(t_9394), .cin(t_12286), .o(t_12287), .co(t_12288), .cout(t_12289));
compressor_3_2 u1_4317(.a(t_11278), .b(t_11275), .cin(t_12289), .o(t_12290), .cout(t_12291));
compressor_4_2 u2_4318(.a(t_11279), .b(t_11276), .c(t_11284), .d(t_11281), .cin(t_9416), .o(t_12292), .co(t_12293), .cout(t_12294));
compressor_4_2 u2_4319(.a(t_11282), .b(t_11289), .c(t_11286), .d(t_9427), .cin(t_12294), .o(t_12295), .co(t_12296), .cout(t_12297));
compressor_4_2 u2_4320(.a(t_11287), .b(t_11294), .c(t_11291), .d(t_9438), .cin(t_12297), .o(t_12298), .co(t_12299), .cout(t_12300));
compressor_4_2 u2_4321(.a(t_11292), .b(t_11299), .c(t_11296), .d(t_9449), .cin(t_12300), .o(t_12301), .co(t_12302), .cout(t_12303));
compressor_4_2 u2_4322(.a(t_11297), .b(t_11304), .c(t_11301), .d(t_9460), .cin(t_12303), .o(t_12304), .co(t_12305), .cout(t_12306));
compressor_4_2 u2_4323(.a(t_11302), .b(t_11309), .c(t_11306), .d(t_9471), .cin(t_12306), .o(t_12307), .co(t_12308), .cout(t_12309));
compressor_4_2 u2_4324(.a(t_11307), .b(t_11314), .c(t_11311), .d(t_9482), .cin(t_12309), .o(t_12310), .co(t_12311), .cout(t_12312));
compressor_4_2 u2_4325(.a(t_11312), .b(t_11319), .c(t_11316), .d(t_9493), .cin(t_12312), .o(t_12313), .co(t_12314), .cout(t_12315));
compressor_3_2 u1_4326(.a(t_11324), .b(t_11321), .cin(t_12315), .o(t_12316), .cout(t_12317));
compressor_3_2 u1_4327(.a(t_11329), .b(t_11326), .cin(t_9511), .o(t_12318), .cout(t_12319));
compressor_3_2 u1_4328(.a(t_11327), .b(t_11334), .cin(t_11331), .o(t_12320), .cout(t_12321));
compressor_3_2 u1_4329(.a(t_11332), .b(t_11339), .cin(t_11336), .o(t_12322), .cout(t_12323));
compressor_3_2 u1_4330(.a(t_11337), .b(t_11344), .cin(t_11341), .o(t_12324), .cout(t_12325));
compressor_3_2 u1_4331(.a(t_11342), .b(t_11349), .cin(t_11346), .o(t_12326), .cout(t_12327));
compressor_3_2 u1_4332(.a(t_11347), .b(t_11354), .cin(t_11351), .o(t_12328), .cout(t_12329));
compressor_3_2 u1_4333(.a(t_11352), .b(t_11359), .cin(t_11356), .o(t_12330), .cout(t_12331));
compressor_3_2 u1_4334(.a(t_11357), .b(t_11364), .cin(t_11361), .o(t_12332), .cout(t_12333));
compressor_3_2 u1_4335(.a(t_11362), .b(t_11369), .cin(t_11366), .o(t_12334), .cout(t_12335));
compressor_3_2 u1_4336(.a(t_11367), .b(t_11374), .cin(t_11371), .o(t_12336), .cout(t_12337));
compressor_3_2 u1_4337(.a(t_11372), .b(t_11379), .cin(t_11376), .o(t_12338), .cout(t_12339));
compressor_3_2 u1_4338(.a(t_11377), .b(t_11384), .cin(t_11381), .o(t_12340), .cout(t_12341));
compressor_3_2 u1_4339(.a(t_11382), .b(t_11389), .cin(t_11386), .o(t_12342), .cout(t_12343));
compressor_3_2 u1_4340(.a(t_11387), .b(t_11394), .cin(t_11391), .o(t_12344), .cout(t_12345));
compressor_3_2 u1_4341(.a(t_11392), .b(t_11399), .cin(t_11396), .o(t_12346), .cout(t_12347));
compressor_3_2 u1_4342(.a(t_11397), .b(t_11401), .cin(t_9627), .o(t_12348), .cout(t_12349));
compressor_3_2 u1_4343(.a(t_11402), .b(t_11404), .cin(t_9633), .o(t_12350), .cout(t_12351));
half_adder u0_4344(.a(t_11405), .b(t_11407), .o(t_12352), .cout(t_12353));
half_adder u0_4345(.a(t_11408), .b(t_11410), .o(t_12354), .cout(t_12355));
half_adder u0_4346(.a(t_11411), .b(t_11413), .o(t_12356), .cout(t_12357));
half_adder u0_4347(.a(t_11414), .b(t_11416), .o(t_12358), .cout(t_12359));
compressor_3_2 u1_4348(.a(t_11417), .b(t_11419), .cin(t_9656), .o(t_12360), .cout(t_12361));
compressor_3_2 u1_4349(.a(t_11420), .b(t_11421), .cin(t_9661), .o(t_12362), .cout(t_12363));
half_adder u0_4350(.a(t_11422), .b(t_11423), .o(t_12364), .cout(t_12365));
half_adder u0_4351(.a(t_11424), .b(t_11425), .o(t_12366), .cout(t_12367));
half_adder u0_4352(.a(t_11426), .b(t_11427), .o(t_12368), .cout(t_12369));
half_adder u0_4353(.a(t_11428), .b(t_11429), .o(t_12370), .cout(t_12371));
half_adder u0_4354(.a(t_11430), .b(t_11431), .o(t_12372), .cout(t_12373));
half_adder u0_4355(.a(t_11432), .b(t_11433), .o(t_12374), .cout(t_12375));
half_adder u0_4356(.a(t_11434), .b(t_11435), .o(t_12376), .cout(t_12377));
half_adder u0_4357(.a(t_11436), .b(t_11437), .o(t_12378), .cout(t_12379));
half_adder u0_4358(.a(t_11438), .b(t_11439), .o(t_12380), .cout(t_12381));
half_adder u0_4359(.a(t_11440), .b(t_11441), .o(t_12382), .cout(t_12383));
half_adder u0_4360(.a(t_11442), .b(t_11443), .o(t_12384), .cout(t_12385));
half_adder u0_4361(.a(t_11444), .b(t_11445), .o(t_12386), .cout(t_12387));
half_adder u0_4362(.a(t_11446), .b(t_11447), .o(t_12388), .cout(t_12389));
half_adder u0_4363(.a(t_11448), .b(t_11449), .o(t_12390), .cout(t_12391));
half_adder u0_4364(.a(t_11450), .b(t_11451), .o(t_12392), .cout(t_12393));
half_adder u0_4365(.a(t_11452), .b(t_11453), .o(t_12394), .cout(t_12395));
half_adder u0_4366(.a(t_11454), .b(t_11455), .o(t_12396), .cout(t_12397));
half_adder u0_4367(.a(t_11456), .b(t_11457), .o(t_12398), .cout(t_12399));
half_adder u0_4368(.a(t_11458), .b(t_11459), .o(t_12400), .cout());

/* u0_4369 Output nets */
wire t_12401,  t_12402;
/* u0_4370 Output nets */
wire t_12403,  t_12404;
/* u0_4371 Output nets */
wire t_12405,  t_12406;
/* u0_4372 Output nets */
wire t_12407,  t_12408;
/* u0_4373 Output nets */
wire t_12409,  t_12410;
/* u0_4374 Output nets */
wire t_12411,  t_12412;
/* u0_4375 Output nets */
wire t_12413,  t_12414;
/* u0_4376 Output nets */
wire t_12415,  t_12416;
/* u0_4377 Output nets */
wire t_12417,  t_12418;
/* u0_4378 Output nets */
wire t_12419,  t_12420;
/* u0_4379 Output nets */
wire t_12421,  t_12422;
/* u0_4380 Output nets */
wire t_12423,  t_12424;
/* u0_4381 Output nets */
wire t_12425,  t_12426;
/* u0_4382 Output nets */
wire t_12427,  t_12428;
/* u0_4383 Output nets */
wire t_12429,  t_12430;
/* u0_4384 Output nets */
wire t_12431,  t_12432;
/* u0_4385 Output nets */
wire t_12433,  t_12434;
/* u0_4386 Output nets */
wire t_12435,  t_12436;
/* u0_4387 Output nets */
wire t_12437,  t_12438;
/* u0_4388 Output nets */
wire t_12439,  t_12440;
/* u0_4389 Output nets */
wire t_12441,  t_12442;
/* u0_4390 Output nets */
wire t_12443,  t_12444;
/* u0_4391 Output nets */
wire t_12445,  t_12446;
/* u0_4392 Output nets */
wire t_12447,  t_12448;
/* u0_4393 Output nets */
wire t_12449,  t_12450;
/* u0_4394 Output nets */
wire t_12451,  t_12452;
/* u0_4395 Output nets */
wire t_12453,  t_12454;
/* u0_4396 Output nets */
wire t_12455,  t_12456;
/* u0_4397 Output nets */
wire t_12457,  t_12458;
/* u0_4398 Output nets */
wire t_12459,  t_12460;
/* u0_4399 Output nets */
wire t_12461,  t_12462;
/* u0_4400 Output nets */
wire t_12463,  t_12464;
/* u0_4401 Output nets */
wire t_12465,  t_12466;
/* u0_4402 Output nets */
wire t_12467,  t_12468;
/* u1_4403 Output nets */
wire t_12469,  t_12470;
/* u0_4404 Output nets */
wire t_12471,  t_12472;
/* u0_4405 Output nets */
wire t_12473,  t_12474;
/* u0_4406 Output nets */
wire t_12475,  t_12476;
/* u0_4407 Output nets */
wire t_12477,  t_12478;
/* u0_4408 Output nets */
wire t_12479,  t_12480;
/* u0_4409 Output nets */
wire t_12481,  t_12482;
/* u0_4410 Output nets */
wire t_12483,  t_12484;
/* u1_4411 Output nets */
wire t_12485,  t_12486;
/* u0_4412 Output nets */
wire t_12487,  t_12488;
/* u0_4413 Output nets */
wire t_12489,  t_12490;
/* u1_4414 Output nets */
wire t_12491,  t_12492;
/* u1_4415 Output nets */
wire t_12493,  t_12494;
/* u0_4416 Output nets */
wire t_12495,  t_12496;
/* u0_4417 Output nets */
wire t_12497,  t_12498;
/* u0_4418 Output nets */
wire t_12499,  t_12500;
/* u0_4419 Output nets */
wire t_12501,  t_12502;
/* u0_4420 Output nets */
wire t_12503,  t_12504;
/* u0_4421 Output nets */
wire t_12505,  t_12506;
/* u1_4422 Output nets */
wire t_12507,  t_12508;
/* u1_4423 Output nets */
wire t_12509,  t_12510;
/* u1_4424 Output nets */
wire t_12511,  t_12512;
/* u1_4425 Output nets */
wire t_12513,  t_12514;
/* u1_4426 Output nets */
wire t_12515,  t_12516;
/* u1_4427 Output nets */
wire t_12517,  t_12518;
/* u1_4428 Output nets */
wire t_12519,  t_12520;
/* u1_4429 Output nets */
wire t_12521,  t_12522;
/* u1_4430 Output nets */
wire t_12523,  t_12524;
/* u1_4431 Output nets */
wire t_12525,  t_12526;
/* u1_4432 Output nets */
wire t_12527,  t_12528;
/* u1_4433 Output nets */
wire t_12529,  t_12530;
/* u1_4434 Output nets */
wire t_12531,  t_12532;
/* u1_4435 Output nets */
wire t_12533,  t_12534;
/* u1_4436 Output nets */
wire t_12535,  t_12536;
/* u1_4437 Output nets */
wire t_12537,  t_12538;
/* u1_4438 Output nets */
wire t_12539,  t_12540;
/* u1_4439 Output nets */
wire t_12541,  t_12542;
/* u1_4440 Output nets */
wire t_12543,  t_12544;
/* u1_4441 Output nets */
wire t_12545,  t_12546;
/* u1_4442 Output nets */
wire t_12547,  t_12548;
/* u1_4443 Output nets */
wire t_12549,  t_12550;
/* u2_4444 Output nets */
wire t_12551,  t_12552,  t_12553;
/* u1_4445 Output nets */
wire t_12554,  t_12555;
/* u1_4446 Output nets */
wire t_12556,  t_12557;
/* u1_4447 Output nets */
wire t_12558,  t_12559;
/* u2_4448 Output nets */
wire t_12560,  t_12561,  t_12562;
/* u1_4449 Output nets */
wire t_12563,  t_12564;
/* u1_4450 Output nets */
wire t_12565,  t_12566;
/* u1_4451 Output nets */
wire t_12567,  t_12568;
/* u1_4452 Output nets */
wire t_12569,  t_12570;
/* u1_4453 Output nets */
wire t_12571,  t_12572;
/* u2_4454 Output nets */
wire t_12573,  t_12574,  t_12575;
/* u2_4455 Output nets */
wire t_12576,  t_12577,  t_12578;
/* u2_4456 Output nets */
wire t_12579,  t_12580,  t_12581;
/* u2_4457 Output nets */
wire t_12582,  t_12583,  t_12584;
/* u2_4458 Output nets */
wire t_12585,  t_12586,  t_12587;
/* u2_4459 Output nets */
wire t_12588,  t_12589,  t_12590;
/* u2_4460 Output nets */
wire t_12591,  t_12592,  t_12593;
/* u2_4461 Output nets */
wire t_12594,  t_12595,  t_12596;
/* u2_4462 Output nets */
wire t_12597,  t_12598,  t_12599;
/* u2_4463 Output nets */
wire t_12600,  t_12601,  t_12602;
/* u2_4464 Output nets */
wire t_12603,  t_12604,  t_12605;
/* u1_4465 Output nets */
wire t_12606,  t_12607;
/* u2_4466 Output nets */
wire t_12608,  t_12609,  t_12610;
/* u2_4467 Output nets */
wire t_12611,  t_12612,  t_12613;
/* u2_4468 Output nets */
wire t_12614,  t_12615,  t_12616;
/* u2_4469 Output nets */
wire t_12617,  t_12618,  t_12619;
/* u1_4470 Output nets */
wire t_12620,  t_12621;
/* u1_4471 Output nets */
wire t_12622,  t_12623;
/* u2_4472 Output nets */
wire t_12624,  t_12625,  t_12626;
/* u2_4473 Output nets */
wire t_12627,  t_12628,  t_12629;
/* u2_4474 Output nets */
wire t_12630,  t_12631,  t_12632;
/* u2_4475 Output nets */
wire t_12633,  t_12634,  t_12635;
/* u2_4476 Output nets */
wire t_12636,  t_12637,  t_12638;
/* u2_4477 Output nets */
wire t_12639,  t_12640,  t_12641;
/* u2_4478 Output nets */
wire t_12642,  t_12643,  t_12644;
/* u1_4479 Output nets */
wire t_12645,  t_12646;
/* u2_4480 Output nets */
wire t_12647,  t_12648,  t_12649;
/* u2_4481 Output nets */
wire t_12650,  t_12651,  t_12652;
/* u2_4482 Output nets */
wire t_12653,  t_12654,  t_12655;
/* u2_4483 Output nets */
wire t_12656,  t_12657,  t_12658;
/* u2_4484 Output nets */
wire t_12659,  t_12660,  t_12661;
/* u2_4485 Output nets */
wire t_12662,  t_12663,  t_12664;
/* u2_4486 Output nets */
wire t_12665,  t_12666,  t_12667;
/* u2_4487 Output nets */
wire t_12668,  t_12669,  t_12670;
/* u2_4488 Output nets */
wire t_12671,  t_12672,  t_12673;
/* u2_4489 Output nets */
wire t_12674,  t_12675,  t_12676;
/* u2_4490 Output nets */
wire t_12677,  t_12678,  t_12679;
/* u2_4491 Output nets */
wire t_12680,  t_12681,  t_12682;
/* u2_4492 Output nets */
wire t_12683,  t_12684,  t_12685;
/* u2_4493 Output nets */
wire t_12686,  t_12687,  t_12688;
/* u2_4494 Output nets */
wire t_12689,  t_12690,  t_12691;
/* u2_4495 Output nets */
wire t_12692,  t_12693,  t_12694;
/* u2_4496 Output nets */
wire t_12695,  t_12696,  t_12697;
/* u2_4497 Output nets */
wire t_12698,  t_12699,  t_12700;
/* u2_4498 Output nets */
wire t_12701,  t_12702,  t_12703;
/* u2_4499 Output nets */
wire t_12704,  t_12705,  t_12706;
/* u2_4500 Output nets */
wire t_12707,  t_12708,  t_12709;
/* u2_4501 Output nets */
wire t_12710,  t_12711,  t_12712;
/* u2_4502 Output nets */
wire t_12713,  t_12714,  t_12715;
/* u2_4503 Output nets */
wire t_12716,  t_12717,  t_12718;
/* u2_4504 Output nets */
wire t_12719,  t_12720,  t_12721;
/* u2_4505 Output nets */
wire t_12722,  t_12723,  t_12724;
/* u2_4506 Output nets */
wire t_12725,  t_12726,  t_12727;
/* u2_4507 Output nets */
wire t_12728,  t_12729,  t_12730;
/* u1_4508 Output nets */
wire t_12731,  t_12732;
/* u2_4509 Output nets */
wire t_12733,  t_12734,  t_12735;
/* u2_4510 Output nets */
wire t_12736,  t_12737,  t_12738;
/* u2_4511 Output nets */
wire t_12739,  t_12740,  t_12741;
/* u2_4512 Output nets */
wire t_12742,  t_12743,  t_12744;
/* u2_4513 Output nets */
wire t_12745,  t_12746,  t_12747;
/* u2_4514 Output nets */
wire t_12748,  t_12749,  t_12750;
/* u2_4515 Output nets */
wire t_12751,  t_12752,  t_12753;
/* u2_4516 Output nets */
wire t_12754,  t_12755,  t_12756;
/* u2_4517 Output nets */
wire t_12757,  t_12758,  t_12759;
/* u2_4518 Output nets */
wire t_12760,  t_12761,  t_12762;
/* u2_4519 Output nets */
wire t_12763,  t_12764,  t_12765;
/* u2_4520 Output nets */
wire t_12766,  t_12767,  t_12768;
/* u2_4521 Output nets */
wire t_12769,  t_12770,  t_12771;
/* u2_4522 Output nets */
wire t_12772,  t_12773,  t_12774;
/* u2_4523 Output nets */
wire t_12775,  t_12776,  t_12777;
/* u2_4524 Output nets */
wire t_12778,  t_12779,  t_12780;
/* u1_4525 Output nets */
wire t_12781,  t_12782;
/* u1_4526 Output nets */
wire t_12783,  t_12784;
/* u1_4527 Output nets */
wire t_12785,  t_12786;
/* u1_4528 Output nets */
wire t_12787,  t_12788;
/* u2_4529 Output nets */
wire t_12789,  t_12790,  t_12791;
/* u1_4530 Output nets */
wire t_12792,  t_12793;
/* u1_4531 Output nets */
wire t_12794,  t_12795;
/* u1_4532 Output nets */
wire t_12796,  t_12797;
/* u1_4533 Output nets */
wire t_12798,  t_12799;
/* u1_4534 Output nets */
wire t_12800,  t_12801;
/* u1_4535 Output nets */
wire t_12802,  t_12803;
/* u1_4536 Output nets */
wire t_12804,  t_12805;
/* u1_4537 Output nets */
wire t_12806,  t_12807;
/* u1_4538 Output nets */
wire t_12808,  t_12809;
/* u1_4539 Output nets */
wire t_12810,  t_12811;
/* u1_4540 Output nets */
wire t_12812,  t_12813;
/* u1_4541 Output nets */
wire t_12814,  t_12815;
/* u1_4542 Output nets */
wire t_12816,  t_12817;
/* u1_4543 Output nets */
wire t_12818,  t_12819;
/* u1_4544 Output nets */
wire t_12820,  t_12821;
/* u1_4545 Output nets */
wire t_12822,  t_12823;
/* u1_4546 Output nets */
wire t_12824,  t_12825;
/* u1_4547 Output nets */
wire t_12826,  t_12827;
/* u1_4548 Output nets */
wire t_12828,  t_12829;
/* u1_4549 Output nets */
wire t_12830,  t_12831;
/* u1_4550 Output nets */
wire t_12832,  t_12833;
/* u1_4551 Output nets */
wire t_12834,  t_12835;
/* u1_4552 Output nets */
wire t_12836,  t_12837;
/* u1_4553 Output nets */
wire t_12838,  t_12839;
/* u1_4554 Output nets */
wire t_12840,  t_12841;
/* u1_4555 Output nets */
wire t_12842,  t_12843;
/* u1_4556 Output nets */
wire t_12844,  t_12845;
/* u1_4557 Output nets */
wire t_12846,  t_12847;
/* u0_4558 Output nets */
wire t_12848,  t_12849;
/* u0_4559 Output nets */
wire t_12850,  t_12851;
/* u0_4560 Output nets */
wire t_12852,  t_12853;
/* u1_4561 Output nets */
wire t_12854,  t_12855;
/* u1_4562 Output nets */
wire t_12856,  t_12857;
/* u0_4563 Output nets */
wire t_12858,  t_12859;
/* u0_4564 Output nets */
wire t_12860,  t_12861;
/* u0_4565 Output nets */
wire t_12862,  t_12863;
/* u0_4566 Output nets */
wire t_12864,  t_12865;
/* u0_4567 Output nets */
wire t_12866,  t_12867;
/* u0_4568 Output nets */
wire t_12868,  t_12869;
/* u0_4569 Output nets */
wire t_12870,  t_12871;
/* u0_4570 Output nets */
wire t_12872,  t_12873;
/* u1_4571 Output nets */
wire t_12874,  t_12875;
/* u1_4572 Output nets */
wire t_12876,  t_12877;
/* u0_4573 Output nets */
wire t_12878,  t_12879;
/* u0_4574 Output nets */
wire t_12880,  t_12881;
/* u0_4575 Output nets */
wire t_12882,  t_12883;
/* u0_4576 Output nets */
wire t_12884,  t_12885;
/* u0_4577 Output nets */
wire t_12886,  t_12887;
/* u0_4578 Output nets */
wire t_12888,  t_12889;
/* u0_4579 Output nets */
wire t_12890,  t_12891;
/* u0_4580 Output nets */
wire t_12892,  t_12893;
/* u0_4581 Output nets */
wire t_12894,  t_12895;
/* u0_4582 Output nets */
wire t_12896,  t_12897;
/* u0_4583 Output nets */
wire t_12898,  t_12899;
/* u0_4584 Output nets */
wire t_12900,  t_12901;
/* u0_4585 Output nets */
wire t_12902,  t_12903;
/* u0_4586 Output nets */
wire t_12904,  t_12905;
/* u0_4587 Output nets */
wire t_12906,  t_12907;
/* u0_4588 Output nets */
wire t_12908,  t_12909;
/* u0_4589 Output nets */
wire t_12910,  t_12911;
/* u0_4590 Output nets */
wire t_12912,  t_12913;
/* u0_4591 Output nets */
wire t_12914,  t_12915;
/* u0_4592 Output nets */
wire t_12916,  t_12917;
/* u0_4593 Output nets */
wire t_12918,  t_12919;
/* u0_4594 Output nets */
wire t_12920,  t_12921;
/* u0_4595 Output nets */
wire t_12922,  t_12923;
/* u0_4596 Output nets */
wire t_12924,  t_12925;
/* u0_4597 Output nets */
wire t_12926,  t_12927;
/* u0_4598 Output nets */
wire t_12928,  t_12929;
/* u0_4599 Output nets */
wire t_12930,  t_12931;
/* u0_4600 Output nets */
wire t_12932,  t_12933;
/* u0_4601 Output nets */
wire t_12934,  t_12935;
/* u0_4602 Output nets */
wire t_12936,  t_12937;
/* u0_4603 Output nets */
wire t_12938,  t_12939;
/* u0_4604 Output nets */
wire t_12940,  t_12941;
/* u0_4605 Output nets */
wire t_12942,  t_12943;
/* u0_4606 Output nets */
wire t_12944,  t_12945;
/* u0_4607 Output nets */
wire t_12946,  t_12947;
/* u0_4608 Output nets */
wire t_12948,  t_12949;
/* u0_4609 Output nets */
wire t_12950,  t_12951;
/* u0_4610 Output nets */
wire t_12952,  t_12953;
/* u0_4611 Output nets */
wire t_12954,  t_12955;
/* u0_4612 Output nets */
wire t_12956,  t_12957;
/* u0_4613 Output nets */
wire t_12958;

/* compress stage 5 */
half_adder u0_4369(.a(t_11461), .b(t_9730), .o(t_12401), .cout(t_12402));
half_adder u0_4370(.a(t_11463), .b(t_9732), .o(t_12403), .cout(t_12404));
half_adder u0_4371(.a(t_11465), .b(t_11466), .o(t_12405), .cout(t_12406));
half_adder u0_4372(.a(t_11467), .b(t_11468), .o(t_12407), .cout(t_12408));
half_adder u0_4373(.a(t_11469), .b(t_11470), .o(t_12409), .cout(t_12410));
half_adder u0_4374(.a(t_11471), .b(t_9740), .o(t_12411), .cout(t_12412));
half_adder u0_4375(.a(t_11473), .b(t_11474), .o(t_12413), .cout(t_12414));
half_adder u0_4376(.a(t_11475), .b(t_11476), .o(t_12415), .cout(t_12416));
half_adder u0_4377(.a(t_11477), .b(t_11478), .o(t_12417), .cout(t_12418));
half_adder u0_4378(.a(t_11479), .b(t_11480), .o(t_12419), .cout(t_12420));
half_adder u0_4379(.a(t_11481), .b(t_11482), .o(t_12421), .cout(t_12422));
half_adder u0_4380(.a(t_11483), .b(t_11484), .o(t_12423), .cout(t_12424));
half_adder u0_4381(.a(t_11485), .b(t_11486), .o(t_12425), .cout(t_12426));
half_adder u0_4382(.a(t_11487), .b(t_11488), .o(t_12427), .cout(t_12428));
half_adder u0_4383(.a(t_11489), .b(t_9760), .o(t_12429), .cout(t_12430));
half_adder u0_4384(.a(t_11491), .b(t_11492), .o(t_12431), .cout(t_12432));
half_adder u0_4385(.a(t_11493), .b(t_9767), .o(t_12433), .cout(t_12434));
half_adder u0_4386(.a(t_11495), .b(t_11496), .o(t_12435), .cout(t_12436));
half_adder u0_4387(.a(t_11497), .b(t_11498), .o(t_12437), .cout(t_12438));
half_adder u0_4388(.a(t_11499), .b(t_11500), .o(t_12439), .cout(t_12440));
half_adder u0_4389(.a(t_11501), .b(t_11502), .o(t_12441), .cout(t_12442));
half_adder u0_4390(.a(t_11503), .b(t_11504), .o(t_12443), .cout(t_12444));
half_adder u0_4391(.a(t_11505), .b(t_11506), .o(t_12445), .cout(t_12446));
half_adder u0_4392(.a(t_11507), .b(t_11508), .o(t_12447), .cout(t_12448));
half_adder u0_4393(.a(t_11509), .b(t_11510), .o(t_12449), .cout(t_12450));
half_adder u0_4394(.a(t_11511), .b(t_11512), .o(t_12451), .cout(t_12452));
half_adder u0_4395(.a(t_11513), .b(t_11514), .o(t_12453), .cout(t_12454));
half_adder u0_4396(.a(t_11515), .b(t_11516), .o(t_12455), .cout(t_12456));
half_adder u0_4397(.a(t_11517), .b(t_11518), .o(t_12457), .cout(t_12458));
half_adder u0_4398(.a(t_11519), .b(t_11520), .o(t_12459), .cout(t_12460));
half_adder u0_4399(.a(t_11521), .b(t_11522), .o(t_12461), .cout(t_12462));
half_adder u0_4400(.a(t_11523), .b(t_11524), .o(t_12463), .cout(t_12464));
half_adder u0_4401(.a(t_11525), .b(t_11526), .o(t_12465), .cout(t_12466));
half_adder u0_4402(.a(t_11527), .b(t_11528), .o(t_12467), .cout(t_12468));
compressor_3_2 u1_4403(.a(t_11531), .b(t_11533), .cin(t_9836), .o(t_12469), .cout(t_12470));
half_adder u0_4404(.a(t_11534), .b(t_11535), .o(t_12471), .cout(t_12472));
half_adder u0_4405(.a(t_11536), .b(t_11537), .o(t_12473), .cout(t_12474));
half_adder u0_4406(.a(t_11538), .b(t_11539), .o(t_12475), .cout(t_12476));
half_adder u0_4407(.a(t_11542), .b(t_11544), .o(t_12477), .cout(t_12478));
half_adder u0_4408(.a(t_11545), .b(t_11547), .o(t_12479), .cout(t_12480));
half_adder u0_4409(.a(t_11548), .b(t_11550), .o(t_12481), .cout(t_12482));
half_adder u0_4410(.a(t_11551), .b(t_11553), .o(t_12483), .cout(t_12484));
compressor_3_2 u1_4411(.a(t_11554), .b(t_11556), .cin(t_9881), .o(t_12485), .cout(t_12486));
half_adder u0_4412(.a(t_11557), .b(t_11558), .o(t_12487), .cout(t_12488));
half_adder u0_4413(.a(t_11559), .b(t_11561), .o(t_12489), .cout(t_12490));
compressor_3_2 u1_4414(.a(t_11562), .b(t_11564), .cin(t_9897), .o(t_12491), .cout(t_12492));
compressor_3_2 u1_4415(.a(t_11565), .b(t_11566), .cin(t_9905), .o(t_12493), .cout(t_12494));
half_adder u0_4416(.a(t_11568), .b(t_9911), .o(t_12495), .cout(t_12496));
half_adder u0_4417(.a(t_11569), .b(t_11571), .o(t_12497), .cout(t_12498));
half_adder u0_4418(.a(t_11572), .b(t_11574), .o(t_12499), .cout(t_12500));
half_adder u0_4419(.a(t_11575), .b(t_11577), .o(t_12501), .cout(t_12502));
half_adder u0_4420(.a(t_11578), .b(t_11580), .o(t_12503), .cout(t_12504));
half_adder u0_4421(.a(t_11581), .b(t_11583), .o(t_12505), .cout(t_12506));
compressor_3_2 u1_4422(.a(t_11584), .b(t_11586), .cin(t_9946), .o(t_12507), .cout(t_12508));
compressor_3_2 u1_4423(.a(t_11587), .b(t_11589), .cin(t_9952), .o(t_12509), .cout(t_12510));
compressor_3_2 u1_4424(.a(t_11590), .b(t_11592), .cin(t_9958), .o(t_12511), .cout(t_12512));
compressor_3_2 u1_4425(.a(t_11593), .b(t_11595), .cin(t_9964), .o(t_12513), .cout(t_12514));
compressor_3_2 u1_4426(.a(t_11596), .b(t_11598), .cin(t_9970), .o(t_12515), .cout(t_12516));
compressor_3_2 u1_4427(.a(t_11599), .b(t_11601), .cin(t_9976), .o(t_12517), .cout(t_12518));
compressor_3_2 u1_4428(.a(t_11602), .b(t_11604), .cin(t_9982), .o(t_12519), .cout(t_12520));
compressor_3_2 u1_4429(.a(t_11605), .b(t_11607), .cin(t_9990), .o(t_12521), .cout(t_12522));
compressor_3_2 u1_4430(.a(t_11608), .b(t_11610), .cin(t_9998), .o(t_12523), .cout(t_12524));
compressor_3_2 u1_4431(.a(t_11611), .b(t_11613), .cin(t_10006), .o(t_12525), .cout(t_12526));
compressor_3_2 u1_4432(.a(t_11614), .b(t_11616), .cin(t_10014), .o(t_12527), .cout(t_12528));
compressor_3_2 u1_4433(.a(t_11617), .b(t_11622), .cin(t_11619), .o(t_12529), .cout(t_12530));
compressor_3_2 u1_4434(.a(t_11620), .b(t_11627), .cin(t_11624), .o(t_12531), .cout(t_12532));
compressor_3_2 u1_4435(.a(t_11625), .b(t_11632), .cin(t_11629), .o(t_12533), .cout(t_12534));
compressor_3_2 u1_4436(.a(t_11630), .b(t_11637), .cin(t_11634), .o(t_12535), .cout(t_12536));
compressor_3_2 u1_4437(.a(t_11635), .b(t_11642), .cin(t_11639), .o(t_12537), .cout(t_12538));
compressor_3_2 u1_4438(.a(t_11640), .b(t_11647), .cin(t_11644), .o(t_12539), .cout(t_12540));
compressor_3_2 u1_4439(.a(t_11645), .b(t_11652), .cin(t_11649), .o(t_12541), .cout(t_12542));
compressor_3_2 u1_4440(.a(t_11650), .b(t_11657), .cin(t_11654), .o(t_12543), .cout(t_12544));
compressor_3_2 u1_4441(.a(t_11655), .b(t_11662), .cin(t_11659), .o(t_12545), .cout(t_12546));
compressor_3_2 u1_4442(.a(t_11660), .b(t_11667), .cin(t_11664), .o(t_12547), .cout(t_12548));
compressor_3_2 u1_4443(.a(t_11665), .b(t_11672), .cin(t_11669), .o(t_12549), .cout(t_12550));
compressor_4_2 u2_4444(.a(t_11670), .b(t_11677), .c(t_11674), .d(t_10113), .cin(t_12550), .o(t_12551), .co(t_12552), .cout(t_12553));
compressor_3_2 u1_4445(.a(t_11682), .b(t_11679), .cin(t_12553), .o(t_12554), .cout(t_12555));
compressor_3_2 u1_4446(.a(t_11680), .b(t_11687), .cin(t_11684), .o(t_12556), .cout(t_12557));
compressor_3_2 u1_4447(.a(t_11685), .b(t_11692), .cin(t_11689), .o(t_12558), .cout(t_12559));
compressor_4_2 u2_4448(.a(t_11690), .b(t_11697), .c(t_11694), .d(t_10147), .cin(t_12559), .o(t_12560), .co(t_12561), .cout(t_12562));
compressor_3_2 u1_4449(.a(t_11702), .b(t_11699), .cin(t_12562), .o(t_12563), .cout(t_12564));
compressor_3_2 u1_4450(.a(t_11700), .b(t_11707), .cin(t_11704), .o(t_12565), .cout(t_12566));
compressor_3_2 u1_4451(.a(t_11705), .b(t_11712), .cin(t_11709), .o(t_12567), .cout(t_12568));
compressor_3_2 u1_4452(.a(t_11710), .b(t_11717), .cin(t_11714), .o(t_12569), .cout(t_12570));
compressor_3_2 u1_4453(.a(t_11715), .b(t_11722), .cin(t_11719), .o(t_12571), .cout(t_12572));
compressor_4_2 u2_4454(.a(t_11720), .b(t_11727), .c(t_11724), .d(t_10200), .cin(t_12572), .o(t_12573), .co(t_12574), .cout(t_12575));
compressor_4_2 u2_4455(.a(t_11725), .b(t_11732), .c(t_11729), .d(t_10209), .cin(t_12575), .o(t_12576), .co(t_12577), .cout(t_12578));
compressor_4_2 u2_4456(.a(t_11730), .b(t_11737), .c(t_11734), .d(t_10218), .cin(t_12578), .o(t_12579), .co(t_12580), .cout(t_12581));
compressor_4_2 u2_4457(.a(t_11735), .b(t_11742), .c(t_11739), .d(t_10227), .cin(t_12581), .o(t_12582), .co(t_12583), .cout(t_12584));
compressor_4_2 u2_4458(.a(t_11740), .b(t_11747), .c(t_11744), .d(t_10236), .cin(t_12584), .o(t_12585), .co(t_12586), .cout(t_12587));
compressor_4_2 u2_4459(.a(t_11745), .b(t_11752), .c(t_11749), .d(t_10245), .cin(t_12587), .o(t_12588), .co(t_12589), .cout(t_12590));
compressor_4_2 u2_4460(.a(t_11750), .b(t_11757), .c(t_11754), .d(t_10254), .cin(t_12590), .o(t_12591), .co(t_12592), .cout(t_12593));
compressor_4_2 u2_4461(.a(t_11755), .b(t_11762), .c(t_11759), .d(t_10265), .cin(t_12593), .o(t_12594), .co(t_12595), .cout(t_12596));
compressor_4_2 u2_4462(.a(t_11760), .b(t_11767), .c(t_11764), .d(t_10276), .cin(t_12596), .o(t_12597), .co(t_12598), .cout(t_12599));
compressor_4_2 u2_4463(.a(t_11765), .b(t_11772), .c(t_11769), .d(t_10287), .cin(t_12599), .o(t_12600), .co(t_12601), .cout(t_12602));
compressor_4_2 u2_4464(.a(t_11770), .b(t_11777), .c(t_11774), .d(t_10298), .cin(t_12602), .o(t_12603), .co(t_12604), .cout(t_12605));
compressor_3_2 u1_4465(.a(t_11782), .b(t_11779), .cin(t_12605), .o(t_12606), .cout(t_12607));
compressor_4_2 u2_4466(.a(t_11783), .b(t_11780), .c(t_11788), .d(t_11785), .cin(t_10320), .o(t_12608), .co(t_12609), .cout(t_12610));
compressor_4_2 u2_4467(.a(t_11786), .b(t_11793), .c(t_11790), .d(t_10331), .cin(t_12610), .o(t_12611), .co(t_12612), .cout(t_12613));
compressor_4_2 u2_4468(.a(t_11791), .b(t_11798), .c(t_11795), .d(t_10342), .cin(t_12613), .o(t_12614), .co(t_12615), .cout(t_12616));
compressor_4_2 u2_4469(.a(t_11796), .b(t_11803), .c(t_11800), .d(t_10353), .cin(t_12616), .o(t_12617), .co(t_12618), .cout(t_12619));
compressor_3_2 u1_4470(.a(t_11808), .b(t_11805), .cin(t_12619), .o(t_12620), .cout(t_12621));
compressor_3_2 u1_4471(.a(t_11806), .b(t_11814), .cin(t_11811), .o(t_12622), .cout(t_12623));
compressor_4_2 u2_4472(.a(t_11815), .b(t_11812), .c(t_11820), .d(t_11817), .cin(t_12623), .o(t_12624), .co(t_12625), .cout(t_12626));
compressor_4_2 u2_4473(.a(t_11821), .b(t_11818), .c(t_11826), .d(t_11823), .cin(t_12626), .o(t_12627), .co(t_12628), .cout(t_12629));
compressor_4_2 u2_4474(.a(t_11827), .b(t_11824), .c(t_11832), .d(t_11829), .cin(t_12629), .o(t_12630), .co(t_12631), .cout(t_12632));
compressor_4_2 u2_4475(.a(t_11830), .b(t_11838), .c(t_11835), .d(t_10419), .cin(t_12632), .o(t_12633), .co(t_12634), .cout(t_12635));
compressor_4_2 u2_4476(.a(t_11836), .b(t_11843), .c(t_11840), .d(t_10433), .cin(t_12635), .o(t_12636), .co(t_12637), .cout(t_12638));
compressor_4_2 u2_4477(.a(t_11844), .b(t_11841), .c(t_11849), .d(t_11846), .cin(t_12638), .o(t_12639), .co(t_12640), .cout(t_12641));
compressor_4_2 u2_4478(.a(t_11847), .b(t_11855), .c(t_11852), .d(t_10453), .cin(t_12641), .o(t_12642), .co(t_12643), .cout(t_12644));
compressor_3_2 u1_4479(.a(t_11860), .b(t_11857), .cin(t_12644), .o(t_12645), .cout(t_12646));
compressor_4_2 u2_4480(.a(t_11861), .b(t_11858), .c(t_11866), .d(t_11863), .cin(t_10479), .o(t_12647), .co(t_12648), .cout(t_12649));
compressor_4_2 u2_4481(.a(t_11867), .b(t_11864), .c(t_11872), .d(t_11869), .cin(t_12649), .o(t_12650), .co(t_12651), .cout(t_12652));
compressor_4_2 u2_4482(.a(t_11873), .b(t_11870), .c(t_11878), .d(t_11875), .cin(t_12652), .o(t_12653), .co(t_12654), .cout(t_12655));
compressor_4_2 u2_4483(.a(t_11879), .b(t_11876), .c(t_11884), .d(t_11881), .cin(t_12655), .o(t_12656), .co(t_12657), .cout(t_12658));
compressor_4_2 u2_4484(.a(t_11885), .b(t_11882), .c(t_11890), .d(t_11887), .cin(t_12658), .o(t_12659), .co(t_12660), .cout(t_12661));
compressor_4_2 u2_4485(.a(t_11891), .b(t_11888), .c(t_11896), .d(t_11893), .cin(t_12661), .o(t_12662), .co(t_12663), .cout(t_12664));
compressor_4_2 u2_4486(.a(t_11894), .b(t_11902), .c(t_11899), .d(t_10550), .cin(t_12664), .o(t_12665), .co(t_12666), .cout(t_12667));
compressor_4_2 u2_4487(.a(t_11900), .b(t_11908), .c(t_11905), .d(t_10562), .cin(t_12667), .o(t_12668), .co(t_12669), .cout(t_12670));
compressor_4_2 u2_4488(.a(t_11909), .b(t_11906), .c(t_11914), .d(t_11911), .cin(t_12670), .o(t_12671), .co(t_12672), .cout(t_12673));
compressor_4_2 u2_4489(.a(t_11915), .b(t_11912), .c(t_11920), .d(t_11917), .cin(t_12673), .o(t_12674), .co(t_12675), .cout(t_12676));
compressor_4_2 u2_4490(.a(t_11918), .b(t_11926), .c(t_11923), .d(t_10598), .cin(t_12676), .o(t_12677), .co(t_12678), .cout(t_12679));
compressor_4_2 u2_4491(.a(t_11927), .b(t_11924), .c(t_11932), .d(t_11929), .cin(t_12679), .o(t_12680), .co(t_12681), .cout(t_12682));
compressor_4_2 u2_4492(.a(t_11930), .b(t_11938), .c(t_11935), .d(t_10622), .cin(t_12682), .o(t_12683), .co(t_12684), .cout(t_12685));
compressor_4_2 u2_4493(.a(t_11939), .b(t_11936), .c(t_11944), .d(t_11941), .cin(t_12685), .o(t_12686), .co(t_12687), .cout(t_12688));
compressor_4_2 u2_4494(.a(t_11945), .b(t_11942), .c(t_11950), .d(t_11947), .cin(t_12688), .o(t_12689), .co(t_12690), .cout(t_12691));
compressor_4_2 u2_4495(.a(t_11951), .b(t_11948), .c(t_11956), .d(t_11953), .cin(t_12691), .o(t_12692), .co(t_12693), .cout(t_12694));
compressor_4_2 u2_4496(.a(t_11957), .b(t_11954), .c(t_11962), .d(t_11959), .cin(t_12694), .o(t_12695), .co(t_12696), .cout(t_12697));
compressor_4_2 u2_4497(.a(t_11960), .b(t_11968), .c(t_11965), .d(t_10682), .cin(t_12697), .o(t_12698), .co(t_12699), .cout(t_12700));
compressor_4_2 u2_4498(.a(t_11966), .b(t_11974), .c(t_11971), .d(t_10691), .cin(t_12700), .o(t_12701), .co(t_12702), .cout(t_12703));
compressor_4_2 u2_4499(.a(t_11972), .b(t_11979), .c(t_11976), .d(t_10705), .cin(t_12703), .o(t_12704), .co(t_12705), .cout(t_12706));
compressor_4_2 u2_4500(.a(t_11980), .b(t_11977), .c(t_11985), .d(t_11982), .cin(t_12706), .o(t_12707), .co(t_12708), .cout(t_12709));
compressor_4_2 u2_4501(.a(t_11986), .b(t_11983), .c(t_11991), .d(t_11988), .cin(t_12709), .o(t_12710), .co(t_12711), .cout(t_12712));
compressor_4_2 u2_4502(.a(t_11992), .b(t_11989), .c(t_11997), .d(t_11994), .cin(t_12712), .o(t_12713), .co(t_12714), .cout(t_12715));
compressor_4_2 u2_4503(.a(t_11998), .b(t_11995), .c(t_12003), .d(t_12000), .cin(t_12715), .o(t_12716), .co(t_12717), .cout(t_12718));
compressor_4_2 u2_4504(.a(t_12004), .b(t_12001), .c(t_12009), .d(t_12006), .cin(t_12718), .o(t_12719), .co(t_12720), .cout(t_12721));
compressor_4_2 u2_4505(.a(t_12010), .b(t_12007), .c(t_12015), .d(t_12012), .cin(t_12721), .o(t_12722), .co(t_12723), .cout(t_12724));
compressor_4_2 u2_4506(.a(t_12016), .b(t_12013), .c(t_12021), .d(t_12018), .cin(t_12724), .o(t_12725), .co(t_12726), .cout(t_12727));
compressor_4_2 u2_4507(.a(t_12019), .b(t_12027), .c(t_12024), .d(t_10791), .cin(t_12727), .o(t_12728), .co(t_12729), .cout(t_12730));
compressor_3_2 u1_4508(.a(t_12032), .b(t_12029), .cin(t_12730), .o(t_12731), .cout(t_12732));
compressor_4_2 u2_4509(.a(t_12033), .b(t_12030), .c(t_12038), .d(t_12035), .cin(t_10813), .o(t_12733), .co(t_12734), .cout(t_12735));
compressor_4_2 u2_4510(.a(t_12036), .b(t_12043), .c(t_12040), .d(t_10824), .cin(t_12735), .o(t_12736), .co(t_12737), .cout(t_12738));
compressor_4_2 u2_4511(.a(t_12041), .b(t_12048), .c(t_12045), .d(t_10835), .cin(t_12738), .o(t_12739), .co(t_12740), .cout(t_12741));
compressor_4_2 u2_4512(.a(t_12046), .b(t_12053), .c(t_12050), .d(t_10846), .cin(t_12741), .o(t_12742), .co(t_12743), .cout(t_12744));
compressor_4_2 u2_4513(.a(t_12051), .b(t_12058), .c(t_12055), .d(t_10857), .cin(t_12744), .o(t_12745), .co(t_12746), .cout(t_12747));
compressor_4_2 u2_4514(.a(t_12056), .b(t_12063), .c(t_12060), .d(t_10868), .cin(t_12747), .o(t_12748), .co(t_12749), .cout(t_12750));
compressor_4_2 u2_4515(.a(t_12061), .b(t_12068), .c(t_12065), .d(t_10879), .cin(t_12750), .o(t_12751), .co(t_12752), .cout(t_12753));
compressor_4_2 u2_4516(.a(t_12066), .b(t_12073), .c(t_12070), .d(t_10890), .cin(t_12753), .o(t_12754), .co(t_12755), .cout(t_12756));
compressor_4_2 u2_4517(.a(t_12071), .b(t_12078), .c(t_12075), .d(t_10901), .cin(t_12756), .o(t_12757), .co(t_12758), .cout(t_12759));
compressor_4_2 u2_4518(.a(t_12076), .b(t_12083), .c(t_12080), .d(t_10912), .cin(t_12759), .o(t_12760), .co(t_12761), .cout(t_12762));
compressor_4_2 u2_4519(.a(t_12081), .b(t_12088), .c(t_12085), .d(t_10923), .cin(t_12762), .o(t_12763), .co(t_12764), .cout(t_12765));
compressor_4_2 u2_4520(.a(t_12086), .b(t_12093), .c(t_12090), .d(t_10934), .cin(t_12765), .o(t_12766), .co(t_12767), .cout(t_12768));
compressor_4_2 u2_4521(.a(t_12091), .b(t_12098), .c(t_12095), .d(t_10945), .cin(t_12768), .o(t_12769), .co(t_12770), .cout(t_12771));
compressor_4_2 u2_4522(.a(t_12096), .b(t_12103), .c(t_12100), .d(t_10956), .cin(t_12771), .o(t_12772), .co(t_12773), .cout(t_12774));
compressor_4_2 u2_4523(.a(t_12101), .b(t_12108), .c(t_12105), .d(t_10967), .cin(t_12774), .o(t_12775), .co(t_12776), .cout(t_12777));
compressor_4_2 u2_4524(.a(t_12106), .b(t_12113), .c(t_12110), .d(t_10978), .cin(t_12777), .o(t_12778), .co(t_12779), .cout(t_12780));
compressor_3_2 u1_4525(.a(t_12118), .b(t_12115), .cin(t_12780), .o(t_12781), .cout(t_12782));
compressor_3_2 u1_4526(.a(t_12116), .b(t_12123), .cin(t_12120), .o(t_12783), .cout(t_12784));
compressor_3_2 u1_4527(.a(t_12121), .b(t_12128), .cin(t_12125), .o(t_12785), .cout(t_12786));
compressor_3_2 u1_4528(.a(t_12126), .b(t_12133), .cin(t_12130), .o(t_12787), .cout(t_12788));
compressor_4_2 u2_4529(.a(t_12131), .b(t_12138), .c(t_12135), .d(t_11023), .cin(t_12788), .o(t_12789), .co(t_12790), .cout(t_12791));
compressor_3_2 u1_4530(.a(t_12143), .b(t_12140), .cin(t_12791), .o(t_12792), .cout(t_12793));
compressor_3_2 u1_4531(.a(t_12148), .b(t_12145), .cin(t_11040), .o(t_12794), .cout(t_12795));
compressor_3_2 u1_4532(.a(t_12146), .b(t_12153), .cin(t_12150), .o(t_12796), .cout(t_12797));
compressor_3_2 u1_4533(.a(t_12151), .b(t_12158), .cin(t_12155), .o(t_12798), .cout(t_12799));
compressor_3_2 u1_4534(.a(t_12156), .b(t_12163), .cin(t_12160), .o(t_12800), .cout(t_12801));
compressor_3_2 u1_4535(.a(t_12161), .b(t_12168), .cin(t_12165), .o(t_12802), .cout(t_12803));
compressor_3_2 u1_4536(.a(t_12166), .b(t_12173), .cin(t_12170), .o(t_12804), .cout(t_12805));
compressor_3_2 u1_4537(.a(t_12171), .b(t_12178), .cin(t_12175), .o(t_12806), .cout(t_12807));
compressor_3_2 u1_4538(.a(t_12176), .b(t_12183), .cin(t_12180), .o(t_12808), .cout(t_12809));
compressor_3_2 u1_4539(.a(t_12181), .b(t_12188), .cin(t_12185), .o(t_12810), .cout(t_12811));
compressor_3_2 u1_4540(.a(t_12186), .b(t_12193), .cin(t_12190), .o(t_12812), .cout(t_12813));
compressor_3_2 u1_4541(.a(t_12191), .b(t_12198), .cin(t_12195), .o(t_12814), .cout(t_12815));
compressor_3_2 u1_4542(.a(t_12196), .b(t_12203), .cin(t_12200), .o(t_12816), .cout(t_12817));
compressor_3_2 u1_4543(.a(t_12201), .b(t_12208), .cin(t_12205), .o(t_12818), .cout(t_12819));
compressor_3_2 u1_4544(.a(t_12206), .b(t_12213), .cin(t_12210), .o(t_12820), .cout(t_12821));
compressor_3_2 u1_4545(.a(t_12211), .b(t_12218), .cin(t_12215), .o(t_12822), .cout(t_12823));
compressor_3_2 u1_4546(.a(t_12216), .b(t_12223), .cin(t_12220), .o(t_12824), .cout(t_12825));
compressor_3_2 u1_4547(.a(t_12221), .b(t_12228), .cin(t_12225), .o(t_12826), .cout(t_12827));
compressor_3_2 u1_4548(.a(t_12226), .b(t_12233), .cin(t_12230), .o(t_12828), .cout(t_12829));
compressor_3_2 u1_4549(.a(t_12231), .b(t_12238), .cin(t_12235), .o(t_12830), .cout(t_12831));
compressor_3_2 u1_4550(.a(t_12236), .b(t_12243), .cin(t_12240), .o(t_12832), .cout(t_12833));
compressor_3_2 u1_4551(.a(t_12241), .b(t_12248), .cin(t_12245), .o(t_12834), .cout(t_12835));
compressor_3_2 u1_4552(.a(t_12246), .b(t_12253), .cin(t_12250), .o(t_12836), .cout(t_12837));
compressor_3_2 u1_4553(.a(t_12251), .b(t_12258), .cin(t_12255), .o(t_12838), .cout(t_12839));
compressor_3_2 u1_4554(.a(t_12256), .b(t_12263), .cin(t_12260), .o(t_12840), .cout(t_12841));
compressor_3_2 u1_4555(.a(t_12261), .b(t_12268), .cin(t_12265), .o(t_12842), .cout(t_12843));
compressor_3_2 u1_4556(.a(t_12266), .b(t_12273), .cin(t_12270), .o(t_12844), .cout(t_12845));
compressor_3_2 u1_4557(.a(t_12271), .b(t_12275), .cin(t_11244), .o(t_12846), .cout(t_12847));
half_adder u0_4558(.a(t_12276), .b(t_12278), .o(t_12848), .cout(t_12849));
half_adder u0_4559(.a(t_12279), .b(t_12281), .o(t_12850), .cout(t_12851));
half_adder u0_4560(.a(t_12282), .b(t_12284), .o(t_12852), .cout(t_12853));
compressor_3_2 u1_4561(.a(t_12285), .b(t_12287), .cin(t_11268), .o(t_12854), .cout(t_12855));
compressor_3_2 u1_4562(.a(t_12288), .b(t_12290), .cin(t_11271), .o(t_12856), .cout(t_12857));
half_adder u0_4563(.a(t_12291), .b(t_12292), .o(t_12858), .cout(t_12859));
half_adder u0_4564(.a(t_12293), .b(t_12295), .o(t_12860), .cout(t_12861));
half_adder u0_4565(.a(t_12296), .b(t_12298), .o(t_12862), .cout(t_12863));
half_adder u0_4566(.a(t_12299), .b(t_12301), .o(t_12864), .cout(t_12865));
half_adder u0_4567(.a(t_12302), .b(t_12304), .o(t_12866), .cout(t_12867));
half_adder u0_4568(.a(t_12305), .b(t_12307), .o(t_12868), .cout(t_12869));
half_adder u0_4569(.a(t_12308), .b(t_12310), .o(t_12870), .cout(t_12871));
half_adder u0_4570(.a(t_12311), .b(t_12313), .o(t_12872), .cout(t_12873));
compressor_3_2 u1_4571(.a(t_12314), .b(t_12316), .cin(t_11317), .o(t_12874), .cout(t_12875));
compressor_3_2 u1_4572(.a(t_12317), .b(t_12318), .cin(t_11322), .o(t_12876), .cout(t_12877));
half_adder u0_4573(.a(t_12319), .b(t_12320), .o(t_12878), .cout(t_12879));
half_adder u0_4574(.a(t_12321), .b(t_12322), .o(t_12880), .cout(t_12881));
half_adder u0_4575(.a(t_12323), .b(t_12324), .o(t_12882), .cout(t_12883));
half_adder u0_4576(.a(t_12325), .b(t_12326), .o(t_12884), .cout(t_12885));
half_adder u0_4577(.a(t_12327), .b(t_12328), .o(t_12886), .cout(t_12887));
half_adder u0_4578(.a(t_12329), .b(t_12330), .o(t_12888), .cout(t_12889));
half_adder u0_4579(.a(t_12331), .b(t_12332), .o(t_12890), .cout(t_12891));
half_adder u0_4580(.a(t_12333), .b(t_12334), .o(t_12892), .cout(t_12893));
half_adder u0_4581(.a(t_12335), .b(t_12336), .o(t_12894), .cout(t_12895));
half_adder u0_4582(.a(t_12337), .b(t_12338), .o(t_12896), .cout(t_12897));
half_adder u0_4583(.a(t_12339), .b(t_12340), .o(t_12898), .cout(t_12899));
half_adder u0_4584(.a(t_12341), .b(t_12342), .o(t_12900), .cout(t_12901));
half_adder u0_4585(.a(t_12343), .b(t_12344), .o(t_12902), .cout(t_12903));
half_adder u0_4586(.a(t_12345), .b(t_12346), .o(t_12904), .cout(t_12905));
half_adder u0_4587(.a(t_12347), .b(t_12348), .o(t_12906), .cout(t_12907));
half_adder u0_4588(.a(t_12349), .b(t_12350), .o(t_12908), .cout(t_12909));
half_adder u0_4589(.a(t_12351), .b(t_12352), .o(t_12910), .cout(t_12911));
half_adder u0_4590(.a(t_12353), .b(t_12354), .o(t_12912), .cout(t_12913));
half_adder u0_4591(.a(t_12355), .b(t_12356), .o(t_12914), .cout(t_12915));
half_adder u0_4592(.a(t_12357), .b(t_12358), .o(t_12916), .cout(t_12917));
half_adder u0_4593(.a(t_12359), .b(t_12360), .o(t_12918), .cout(t_12919));
half_adder u0_4594(.a(t_12361), .b(t_12362), .o(t_12920), .cout(t_12921));
half_adder u0_4595(.a(t_12363), .b(t_12364), .o(t_12922), .cout(t_12923));
half_adder u0_4596(.a(t_12365), .b(t_12366), .o(t_12924), .cout(t_12925));
half_adder u0_4597(.a(t_12367), .b(t_12368), .o(t_12926), .cout(t_12927));
half_adder u0_4598(.a(t_12369), .b(t_12370), .o(t_12928), .cout(t_12929));
half_adder u0_4599(.a(t_12371), .b(t_12372), .o(t_12930), .cout(t_12931));
half_adder u0_4600(.a(t_12373), .b(t_12374), .o(t_12932), .cout(t_12933));
half_adder u0_4601(.a(t_12375), .b(t_12376), .o(t_12934), .cout(t_12935));
half_adder u0_4602(.a(t_12377), .b(t_12378), .o(t_12936), .cout(t_12937));
half_adder u0_4603(.a(t_12379), .b(t_12380), .o(t_12938), .cout(t_12939));
half_adder u0_4604(.a(t_12381), .b(t_12382), .o(t_12940), .cout(t_12941));
half_adder u0_4605(.a(t_12383), .b(t_12384), .o(t_12942), .cout(t_12943));
half_adder u0_4606(.a(t_12385), .b(t_12386), .o(t_12944), .cout(t_12945));
half_adder u0_4607(.a(t_12387), .b(t_12388), .o(t_12946), .cout(t_12947));
half_adder u0_4608(.a(t_12389), .b(t_12390), .o(t_12948), .cout(t_12949));
half_adder u0_4609(.a(t_12391), .b(t_12392), .o(t_12950), .cout(t_12951));
half_adder u0_4610(.a(t_12393), .b(t_12394), .o(t_12952), .cout(t_12953));
half_adder u0_4611(.a(t_12395), .b(t_12396), .o(t_12954), .cout(t_12955));
half_adder u0_4612(.a(t_12397), .b(t_12398), .o(t_12956), .cout(t_12957));
half_adder u0_4613(.a(t_12399), .b(t_12400), .o(t_12958), .cout());

/* u0_4614 Output nets */
wire t_12959,  t_12960;
/* u0_4615 Output nets */
wire t_12961,  t_12962;
/* u0_4616 Output nets */
wire t_12963,  t_12964;
/* u0_4617 Output nets */
wire t_12965,  t_12966;
/* u0_4618 Output nets */
wire t_12967,  t_12968;
/* u0_4619 Output nets */
wire t_12969,  t_12970;
/* u0_4620 Output nets */
wire t_12971,  t_12972;
/* u0_4621 Output nets */
wire t_12973,  t_12974;
/* u0_4622 Output nets */
wire t_12975,  t_12976;
/* u0_4623 Output nets */
wire t_12977,  t_12978;
/* u0_4624 Output nets */
wire t_12979,  t_12980;
/* u0_4625 Output nets */
wire t_12981,  t_12982;
/* u0_4626 Output nets */
wire t_12983,  t_12984;
/* u0_4627 Output nets */
wire t_12985,  t_12986;
/* u0_4628 Output nets */
wire t_12987,  t_12988;
/* u0_4629 Output nets */
wire t_12989,  t_12990;
/* u0_4630 Output nets */
wire t_12991,  t_12992;
/* u0_4631 Output nets */
wire t_12993,  t_12994;
/* u0_4632 Output nets */
wire t_12995,  t_12996;
/* u0_4633 Output nets */
wire t_12997,  t_12998;
/* u0_4634 Output nets */
wire t_12999,  t_13000;
/* u0_4635 Output nets */
wire t_13001,  t_13002;
/* u0_4636 Output nets */
wire t_13003,  t_13004;
/* u0_4637 Output nets */
wire t_13005,  t_13006;
/* u0_4638 Output nets */
wire t_13007,  t_13008;
/* u0_4639 Output nets */
wire t_13009,  t_13010;
/* u0_4640 Output nets */
wire t_13011,  t_13012;
/* u0_4641 Output nets */
wire t_13013,  t_13014;
/* u0_4642 Output nets */
wire t_13015,  t_13016;
/* u0_4643 Output nets */
wire t_13017,  t_13018;
/* u0_4644 Output nets */
wire t_13019,  t_13020;
/* u0_4645 Output nets */
wire t_13021,  t_13022;
/* u0_4646 Output nets */
wire t_13023,  t_13024;
/* u0_4647 Output nets */
wire t_13025,  t_13026;
/* u0_4648 Output nets */
wire t_13027,  t_13028;
/* u0_4649 Output nets */
wire t_13029,  t_13030;
/* u0_4650 Output nets */
wire t_13031,  t_13032;
/* u0_4651 Output nets */
wire t_13033,  t_13034;
/* u0_4652 Output nets */
wire t_13035,  t_13036;
/* u0_4653 Output nets */
wire t_13037,  t_13038;
/* u0_4654 Output nets */
wire t_13039,  t_13040;
/* u0_4655 Output nets */
wire t_13041,  t_13042;
/* u0_4656 Output nets */
wire t_13043,  t_13044;
/* u0_4657 Output nets */
wire t_13045,  t_13046;
/* u0_4658 Output nets */
wire t_13047,  t_13048;
/* u0_4659 Output nets */
wire t_13049,  t_13050;
/* u0_4660 Output nets */
wire t_13051,  t_13052;
/* u0_4661 Output nets */
wire t_13053,  t_13054;
/* u0_4662 Output nets */
wire t_13055,  t_13056;
/* u0_4663 Output nets */
wire t_13057,  t_13058;
/* u0_4664 Output nets */
wire t_13059,  t_13060;
/* u0_4665 Output nets */
wire t_13061,  t_13062;
/* u0_4666 Output nets */
wire t_13063,  t_13064;
/* u0_4667 Output nets */
wire t_13065,  t_13066;
/* u0_4668 Output nets */
wire t_13067,  t_13068;
/* u0_4669 Output nets */
wire t_13069,  t_13070;
/* u0_4670 Output nets */
wire t_13071,  t_13072;
/* u0_4671 Output nets */
wire t_13073,  t_13074;
/* u0_4672 Output nets */
wire t_13075,  t_13076;
/* u0_4673 Output nets */
wire t_13077,  t_13078;
/* u0_4674 Output nets */
wire t_13079,  t_13080;
/* u0_4675 Output nets */
wire t_13081,  t_13082;
/* u0_4676 Output nets */
wire t_13083,  t_13084;
/* u0_4677 Output nets */
wire t_13085,  t_13086;
/* u0_4678 Output nets */
wire t_13087,  t_13088;
/* u0_4679 Output nets */
wire t_13089,  t_13090;
/* u0_4680 Output nets */
wire t_13091,  t_13092;
/* u0_4681 Output nets */
wire t_13093,  t_13094;
/* u0_4682 Output nets */
wire t_13095,  t_13096;
/* u0_4683 Output nets */
wire t_13097,  t_13098;
/* u0_4684 Output nets */
wire t_13099,  t_13100;
/* u0_4685 Output nets */
wire t_13101,  t_13102;
/* u0_4686 Output nets */
wire t_13103,  t_13104;
/* u0_4687 Output nets */
wire t_13105,  t_13106;
/* u1_4688 Output nets */
wire t_13107,  t_13108;
/* u0_4689 Output nets */
wire t_13109,  t_13110;
/* u0_4690 Output nets */
wire t_13111,  t_13112;
/* u1_4691 Output nets */
wire t_13113,  t_13114;
/* u0_4692 Output nets */
wire t_13115,  t_13116;
/* u0_4693 Output nets */
wire t_13117,  t_13118;
/* u0_4694 Output nets */
wire t_13119,  t_13120;
/* u0_4695 Output nets */
wire t_13121,  t_13122;
/* u0_4696 Output nets */
wire t_13123,  t_13124;
/* u0_4697 Output nets */
wire t_13125,  t_13126;
/* u0_4698 Output nets */
wire t_13127,  t_13128;
/* u0_4699 Output nets */
wire t_13129,  t_13130;
/* u0_4700 Output nets */
wire t_13131,  t_13132;
/* u0_4701 Output nets */
wire t_13133,  t_13134;
/* u0_4702 Output nets */
wire t_13135,  t_13136;
/* u0_4703 Output nets */
wire t_13137,  t_13138;
/* u0_4704 Output nets */
wire t_13139,  t_13140;
/* u0_4705 Output nets */
wire t_13141,  t_13142;
/* u1_4706 Output nets */
wire t_13143,  t_13144;
/* u0_4707 Output nets */
wire t_13145,  t_13146;
/* u0_4708 Output nets */
wire t_13147,  t_13148;
/* u0_4709 Output nets */
wire t_13149,  t_13150;
/* u0_4710 Output nets */
wire t_13151,  t_13152;
/* u1_4711 Output nets */
wire t_13153,  t_13154;
/* u1_4712 Output nets */
wire t_13155,  t_13156;
/* u0_4713 Output nets */
wire t_13157,  t_13158;
/* u0_4714 Output nets */
wire t_13159,  t_13160;
/* u1_4715 Output nets */
wire t_13161,  t_13162;
/* u0_4716 Output nets */
wire t_13163,  t_13164;
/* u0_4717 Output nets */
wire t_13165,  t_13166;
/* u1_4718 Output nets */
wire t_13167,  t_13168;
/* u1_4719 Output nets */
wire t_13169,  t_13170;
/* u0_4720 Output nets */
wire t_13171,  t_13172;
/* u0_4721 Output nets */
wire t_13173,  t_13174;
/* u0_4722 Output nets */
wire t_13175,  t_13176;
/* u0_4723 Output nets */
wire t_13177,  t_13178;
/* u0_4724 Output nets */
wire t_13179,  t_13180;
/* u0_4725 Output nets */
wire t_13181,  t_13182;
/* u1_4726 Output nets */
wire t_13183,  t_13184;
/* u1_4727 Output nets */
wire t_13185,  t_13186;
/* u0_4728 Output nets */
wire t_13187,  t_13188;
/* u0_4729 Output nets */
wire t_13189,  t_13190;
/* u1_4730 Output nets */
wire t_13191,  t_13192;
/* u0_4731 Output nets */
wire t_13193,  t_13194;
/* u1_4732 Output nets */
wire t_13195,  t_13196;
/* u0_4733 Output nets */
wire t_13197,  t_13198;
/* u0_4734 Output nets */
wire t_13199,  t_13200;
/* u0_4735 Output nets */
wire t_13201,  t_13202;
/* u0_4736 Output nets */
wire t_13203,  t_13204;
/* u1_4737 Output nets */
wire t_13205,  t_13206;
/* u1_4738 Output nets */
wire t_13207,  t_13208;
/* u0_4739 Output nets */
wire t_13209,  t_13210;
/* u0_4740 Output nets */
wire t_13211,  t_13212;
/* u0_4741 Output nets */
wire t_13213,  t_13214;
/* u0_4742 Output nets */
wire t_13215,  t_13216;
/* u0_4743 Output nets */
wire t_13217,  t_13218;
/* u0_4744 Output nets */
wire t_13219,  t_13220;
/* u0_4745 Output nets */
wire t_13221,  t_13222;
/* u0_4746 Output nets */
wire t_13223,  t_13224;
/* u1_4747 Output nets */
wire t_13225,  t_13226;
/* u1_4748 Output nets */
wire t_13227,  t_13228;
/* u0_4749 Output nets */
wire t_13229,  t_13230;
/* u0_4750 Output nets */
wire t_13231,  t_13232;
/* u0_4751 Output nets */
wire t_13233,  t_13234;
/* u0_4752 Output nets */
wire t_13235,  t_13236;
/* u0_4753 Output nets */
wire t_13237,  t_13238;
/* u0_4754 Output nets */
wire t_13239,  t_13240;
/* u0_4755 Output nets */
wire t_13241,  t_13242;
/* u0_4756 Output nets */
wire t_13243,  t_13244;
/* u0_4757 Output nets */
wire t_13245,  t_13246;
/* u0_4758 Output nets */
wire t_13247,  t_13248;
/* u0_4759 Output nets */
wire t_13249,  t_13250;
/* u0_4760 Output nets */
wire t_13251,  t_13252;
/* u0_4761 Output nets */
wire t_13253,  t_13254;
/* u0_4762 Output nets */
wire t_13255,  t_13256;
/* u0_4763 Output nets */
wire t_13257,  t_13258;
/* u0_4764 Output nets */
wire t_13259,  t_13260;
/* u1_4765 Output nets */
wire t_13261,  t_13262;
/* u0_4766 Output nets */
wire t_13263,  t_13264;
/* u0_4767 Output nets */
wire t_13265,  t_13266;
/* u0_4768 Output nets */
wire t_13267,  t_13268;
/* u1_4769 Output nets */
wire t_13269,  t_13270;
/* u1_4770 Output nets */
wire t_13271,  t_13272;
/* u0_4771 Output nets */
wire t_13273,  t_13274;
/* u0_4772 Output nets */
wire t_13275,  t_13276;
/* u0_4773 Output nets */
wire t_13277,  t_13278;
/* u0_4774 Output nets */
wire t_13279,  t_13280;
/* u0_4775 Output nets */
wire t_13281,  t_13282;
/* u0_4776 Output nets */
wire t_13283,  t_13284;
/* u0_4777 Output nets */
wire t_13285,  t_13286;
/* u0_4778 Output nets */
wire t_13287,  t_13288;
/* u0_4779 Output nets */
wire t_13289,  t_13290;
/* u0_4780 Output nets */
wire t_13291,  t_13292;
/* u0_4781 Output nets */
wire t_13293,  t_13294;
/* u0_4782 Output nets */
wire t_13295,  t_13296;
/* u0_4783 Output nets */
wire t_13297,  t_13298;
/* u0_4784 Output nets */
wire t_13299,  t_13300;
/* u0_4785 Output nets */
wire t_13301,  t_13302;
/* u0_4786 Output nets */
wire t_13303,  t_13304;
/* u0_4787 Output nets */
wire t_13305,  t_13306;
/* u0_4788 Output nets */
wire t_13307,  t_13308;
/* u0_4789 Output nets */
wire t_13309,  t_13310;
/* u0_4790 Output nets */
wire t_13311,  t_13312;
/* u0_4791 Output nets */
wire t_13313,  t_13314;
/* u0_4792 Output nets */
wire t_13315,  t_13316;
/* u0_4793 Output nets */
wire t_13317,  t_13318;
/* u0_4794 Output nets */
wire t_13319,  t_13320;
/* u0_4795 Output nets */
wire t_13321,  t_13322;
/* u0_4796 Output nets */
wire t_13323,  t_13324;
/* u0_4797 Output nets */
wire t_13325,  t_13326;
/* u0_4798 Output nets */
wire t_13327,  t_13328;
/* u0_4799 Output nets */
wire t_13329,  t_13330;
/* u0_4800 Output nets */
wire t_13331,  t_13332;
/* u0_4801 Output nets */
wire t_13333,  t_13334;
/* u0_4802 Output nets */
wire t_13335,  t_13336;
/* u0_4803 Output nets */
wire t_13337,  t_13338;
/* u0_4804 Output nets */
wire t_13339,  t_13340;
/* u0_4805 Output nets */
wire t_13341,  t_13342;
/* u0_4806 Output nets */
wire t_13343,  t_13344;
/* u0_4807 Output nets */
wire t_13345,  t_13346;
/* u0_4808 Output nets */
wire t_13347,  t_13348;
/* u0_4809 Output nets */
wire t_13349,  t_13350;
/* u0_4810 Output nets */
wire t_13351,  t_13352;
/* u0_4811 Output nets */
wire t_13353,  t_13354;
/* u0_4812 Output nets */
wire t_13355,  t_13356;
/* u0_4813 Output nets */
wire t_13357,  t_13358;
/* u0_4814 Output nets */
wire t_13359,  t_13360;
/* u0_4815 Output nets */
wire t_13361,  t_13362;
/* u0_4816 Output nets */
wire t_13363,  t_13364;
/* u0_4817 Output nets */
wire t_13365,  t_13366;
/* u0_4818 Output nets */
wire t_13367,  t_13368;
/* u0_4819 Output nets */
wire t_13369,  t_13370;
/* u0_4820 Output nets */
wire t_13371,  t_13372;
/* u0_4821 Output nets */
wire t_13373,  t_13374;
/* u0_4822 Output nets */
wire t_13375,  t_13376;
/* u0_4823 Output nets */
wire t_13377,  t_13378;
/* u0_4824 Output nets */
wire t_13379,  t_13380;
/* u0_4825 Output nets */
wire t_13381,  t_13382;
/* u0_4826 Output nets */
wire t_13383,  t_13384;
/* u0_4827 Output nets */
wire t_13385,  t_13386;
/* u0_4828 Output nets */
wire t_13387,  t_13388;
/* u0_4829 Output nets */
wire t_13389,  t_13390;
/* u0_4830 Output nets */
wire t_13391,  t_13392;
/* u0_4831 Output nets */
wire t_13393,  t_13394;
/* u0_4832 Output nets */
wire t_13395,  t_13396;
/* u0_4833 Output nets */
wire t_13397,  t_13398;
/* u0_4834 Output nets */
wire t_13399,  t_13400;
/* u0_4835 Output nets */
wire t_13401,  t_13402;
/* u0_4836 Output nets */
wire t_13403,  t_13404;
/* u0_4837 Output nets */
wire t_13405,  t_13406;
/* u0_4838 Output nets */
wire t_13407,  t_13408;
/* u0_4839 Output nets */
wire t_13409,  t_13410;
/* u0_4840 Output nets */
wire t_13411,  t_13412;
/* u0_4841 Output nets */
wire t_13413,  t_13414;
/* u0_4842 Output nets */
wire t_13415,  t_13416;
/* u0_4843 Output nets */
wire t_13417,  t_13418;
/* u0_4844 Output nets */
wire t_13419,  t_13420;
/* u0_4845 Output nets */
wire t_13421,  t_13422;
/* u0_4846 Output nets */
wire t_13423,  t_13424;
/* u0_4847 Output nets */
wire t_13425,  t_13426;
/* u0_4848 Output nets */
wire t_13427,  t_13428;
/* u0_4849 Output nets */
wire t_13429,  t_13430;
/* u0_4850 Output nets */
wire t_13431,  t_13432;
/* u0_4851 Output nets */
wire t_13433,  t_13434;
/* u0_4852 Output nets */
wire t_13435;

/* compress stage 6 */
half_adder u0_4614(.a(t_12402), .b(t_11462), .o(t_12959), .cout(t_12960));
half_adder u0_4615(.a(t_12404), .b(t_11464), .o(t_12961), .cout(t_12962));
half_adder u0_4616(.a(t_12406), .b(t_12407), .o(t_12963), .cout(t_12964));
half_adder u0_4617(.a(t_12408), .b(t_12409), .o(t_12965), .cout(t_12966));
half_adder u0_4618(.a(t_12410), .b(t_12411), .o(t_12967), .cout(t_12968));
half_adder u0_4619(.a(t_12412), .b(t_11472), .o(t_12969), .cout(t_12970));
half_adder u0_4620(.a(t_12414), .b(t_12415), .o(t_12971), .cout(t_12972));
half_adder u0_4621(.a(t_12416), .b(t_12417), .o(t_12973), .cout(t_12974));
half_adder u0_4622(.a(t_12418), .b(t_12419), .o(t_12975), .cout(t_12976));
half_adder u0_4623(.a(t_12420), .b(t_12421), .o(t_12977), .cout(t_12978));
half_adder u0_4624(.a(t_12422), .b(t_12423), .o(t_12979), .cout(t_12980));
half_adder u0_4625(.a(t_12424), .b(t_12425), .o(t_12981), .cout(t_12982));
half_adder u0_4626(.a(t_12426), .b(t_12427), .o(t_12983), .cout(t_12984));
half_adder u0_4627(.a(t_12428), .b(t_12429), .o(t_12985), .cout(t_12986));
half_adder u0_4628(.a(t_12430), .b(t_11490), .o(t_12987), .cout(t_12988));
half_adder u0_4629(.a(t_12432), .b(t_12433), .o(t_12989), .cout(t_12990));
half_adder u0_4630(.a(t_12434), .b(t_11494), .o(t_12991), .cout(t_12992));
half_adder u0_4631(.a(t_12436), .b(t_12437), .o(t_12993), .cout(t_12994));
half_adder u0_4632(.a(t_12438), .b(t_12439), .o(t_12995), .cout(t_12996));
half_adder u0_4633(.a(t_12440), .b(t_12441), .o(t_12997), .cout(t_12998));
half_adder u0_4634(.a(t_12442), .b(t_12443), .o(t_12999), .cout(t_13000));
half_adder u0_4635(.a(t_12444), .b(t_12445), .o(t_13001), .cout(t_13002));
half_adder u0_4636(.a(t_12446), .b(t_12447), .o(t_13003), .cout(t_13004));
half_adder u0_4637(.a(t_12448), .b(t_12449), .o(t_13005), .cout(t_13006));
half_adder u0_4638(.a(t_12450), .b(t_12451), .o(t_13007), .cout(t_13008));
half_adder u0_4639(.a(t_12452), .b(t_12453), .o(t_13009), .cout(t_13010));
half_adder u0_4640(.a(t_12454), .b(t_12455), .o(t_13011), .cout(t_13012));
half_adder u0_4641(.a(t_12456), .b(t_12457), .o(t_13013), .cout(t_13014));
half_adder u0_4642(.a(t_12458), .b(t_12459), .o(t_13015), .cout(t_13016));
half_adder u0_4643(.a(t_12460), .b(t_12461), .o(t_13017), .cout(t_13018));
half_adder u0_4644(.a(t_12462), .b(t_12463), .o(t_13019), .cout(t_13020));
half_adder u0_4645(.a(t_12464), .b(t_12465), .o(t_13021), .cout(t_13022));
half_adder u0_4646(.a(t_12466), .b(t_12467), .o(t_13023), .cout(t_13024));
half_adder u0_4647(.a(t_12468), .b(t_11530), .o(t_13025), .cout(t_13026));
half_adder u0_4648(.a(t_12470), .b(t_12471), .o(t_13027), .cout(t_13028));
half_adder u0_4649(.a(t_12472), .b(t_12473), .o(t_13029), .cout(t_13030));
half_adder u0_4650(.a(t_12474), .b(t_12475), .o(t_13031), .cout(t_13032));
half_adder u0_4651(.a(t_12476), .b(t_11541), .o(t_13033), .cout(t_13034));
half_adder u0_4652(.a(t_12478), .b(t_12479), .o(t_13035), .cout(t_13036));
half_adder u0_4653(.a(t_12480), .b(t_12481), .o(t_13037), .cout(t_13038));
half_adder u0_4654(.a(t_12482), .b(t_12483), .o(t_13039), .cout(t_13040));
half_adder u0_4655(.a(t_12484), .b(t_12485), .o(t_13041), .cout(t_13042));
half_adder u0_4656(.a(t_12486), .b(t_12487), .o(t_13043), .cout(t_13044));
half_adder u0_4657(.a(t_12488), .b(t_12489), .o(t_13045), .cout(t_13046));
half_adder u0_4658(.a(t_12490), .b(t_12491), .o(t_13047), .cout(t_13048));
half_adder u0_4659(.a(t_12492), .b(t_12493), .o(t_13049), .cout(t_13050));
half_adder u0_4660(.a(t_12494), .b(t_12495), .o(t_13051), .cout(t_13052));
half_adder u0_4661(.a(t_12496), .b(t_12497), .o(t_13053), .cout(t_13054));
half_adder u0_4662(.a(t_12498), .b(t_12499), .o(t_13055), .cout(t_13056));
half_adder u0_4663(.a(t_12500), .b(t_12501), .o(t_13057), .cout(t_13058));
half_adder u0_4664(.a(t_12502), .b(t_12503), .o(t_13059), .cout(t_13060));
half_adder u0_4665(.a(t_12504), .b(t_12505), .o(t_13061), .cout(t_13062));
half_adder u0_4666(.a(t_12506), .b(t_12507), .o(t_13063), .cout(t_13064));
half_adder u0_4667(.a(t_12508), .b(t_12509), .o(t_13065), .cout(t_13066));
half_adder u0_4668(.a(t_12510), .b(t_12511), .o(t_13067), .cout(t_13068));
half_adder u0_4669(.a(t_12512), .b(t_12513), .o(t_13069), .cout(t_13070));
half_adder u0_4670(.a(t_12514), .b(t_12515), .o(t_13071), .cout(t_13072));
half_adder u0_4671(.a(t_12516), .b(t_12517), .o(t_13073), .cout(t_13074));
half_adder u0_4672(.a(t_12518), .b(t_12519), .o(t_13075), .cout(t_13076));
half_adder u0_4673(.a(t_12520), .b(t_12521), .o(t_13077), .cout(t_13078));
half_adder u0_4674(.a(t_12522), .b(t_12523), .o(t_13079), .cout(t_13080));
half_adder u0_4675(.a(t_12524), .b(t_12525), .o(t_13081), .cout(t_13082));
half_adder u0_4676(.a(t_12526), .b(t_12527), .o(t_13083), .cout(t_13084));
half_adder u0_4677(.a(t_12528), .b(t_12529), .o(t_13085), .cout(t_13086));
half_adder u0_4678(.a(t_12530), .b(t_12531), .o(t_13087), .cout(t_13088));
half_adder u0_4679(.a(t_12532), .b(t_12533), .o(t_13089), .cout(t_13090));
half_adder u0_4680(.a(t_12534), .b(t_12535), .o(t_13091), .cout(t_13092));
half_adder u0_4681(.a(t_12536), .b(t_12537), .o(t_13093), .cout(t_13094));
half_adder u0_4682(.a(t_12538), .b(t_12539), .o(t_13095), .cout(t_13096));
half_adder u0_4683(.a(t_12540), .b(t_12541), .o(t_13097), .cout(t_13098));
half_adder u0_4684(.a(t_12542), .b(t_12543), .o(t_13099), .cout(t_13100));
half_adder u0_4685(.a(t_12544), .b(t_12545), .o(t_13101), .cout(t_13102));
half_adder u0_4686(.a(t_12546), .b(t_12547), .o(t_13103), .cout(t_13104));
half_adder u0_4687(.a(t_12548), .b(t_12549), .o(t_13105), .cout(t_13106));
compressor_3_2 u1_4688(.a(t_12552), .b(t_12554), .cin(t_11675), .o(t_13107), .cout(t_13108));
half_adder u0_4689(.a(t_12555), .b(t_12556), .o(t_13109), .cout(t_13110));
half_adder u0_4690(.a(t_12557), .b(t_12558), .o(t_13111), .cout(t_13112));
compressor_3_2 u1_4691(.a(t_12561), .b(t_12563), .cin(t_11695), .o(t_13113), .cout(t_13114));
half_adder u0_4692(.a(t_12564), .b(t_12565), .o(t_13115), .cout(t_13116));
half_adder u0_4693(.a(t_12566), .b(t_12567), .o(t_13117), .cout(t_13118));
half_adder u0_4694(.a(t_12568), .b(t_12569), .o(t_13119), .cout(t_13120));
half_adder u0_4695(.a(t_12570), .b(t_12571), .o(t_13121), .cout(t_13122));
half_adder u0_4696(.a(t_12574), .b(t_12576), .o(t_13123), .cout(t_13124));
half_adder u0_4697(.a(t_12577), .b(t_12579), .o(t_13125), .cout(t_13126));
half_adder u0_4698(.a(t_12580), .b(t_12582), .o(t_13127), .cout(t_13128));
half_adder u0_4699(.a(t_12583), .b(t_12585), .o(t_13129), .cout(t_13130));
half_adder u0_4700(.a(t_12586), .b(t_12588), .o(t_13131), .cout(t_13132));
half_adder u0_4701(.a(t_12589), .b(t_12591), .o(t_13133), .cout(t_13134));
half_adder u0_4702(.a(t_12592), .b(t_12594), .o(t_13135), .cout(t_13136));
half_adder u0_4703(.a(t_12595), .b(t_12597), .o(t_13137), .cout(t_13138));
half_adder u0_4704(.a(t_12598), .b(t_12600), .o(t_13139), .cout(t_13140));
half_adder u0_4705(.a(t_12601), .b(t_12603), .o(t_13141), .cout(t_13142));
compressor_3_2 u1_4706(.a(t_12604), .b(t_12606), .cin(t_11775), .o(t_13143), .cout(t_13144));
half_adder u0_4707(.a(t_12607), .b(t_12608), .o(t_13145), .cout(t_13146));
half_adder u0_4708(.a(t_12609), .b(t_12611), .o(t_13147), .cout(t_13148));
half_adder u0_4709(.a(t_12612), .b(t_12614), .o(t_13149), .cout(t_13150));
half_adder u0_4710(.a(t_12615), .b(t_12617), .o(t_13151), .cout(t_13152));
compressor_3_2 u1_4711(.a(t_12618), .b(t_12620), .cin(t_11801), .o(t_13153), .cout(t_13154));
compressor_3_2 u1_4712(.a(t_12621), .b(t_12622), .cin(t_11809), .o(t_13155), .cout(t_13156));
half_adder u0_4713(.a(t_12625), .b(t_12627), .o(t_13157), .cout(t_13158));
half_adder u0_4714(.a(t_12628), .b(t_12630), .o(t_13159), .cout(t_13160));
compressor_3_2 u1_4715(.a(t_12631), .b(t_12633), .cin(t_11833), .o(t_13161), .cout(t_13162));
half_adder u0_4716(.a(t_12634), .b(t_12636), .o(t_13163), .cout(t_13164));
half_adder u0_4717(.a(t_12637), .b(t_12639), .o(t_13165), .cout(t_13166));
compressor_3_2 u1_4718(.a(t_12640), .b(t_12642), .cin(t_11850), .o(t_13167), .cout(t_13168));
compressor_3_2 u1_4719(.a(t_12643), .b(t_12645), .cin(t_11853), .o(t_13169), .cout(t_13170));
half_adder u0_4720(.a(t_12646), .b(t_12647), .o(t_13171), .cout(t_13172));
half_adder u0_4721(.a(t_12648), .b(t_12650), .o(t_13173), .cout(t_13174));
half_adder u0_4722(.a(t_12651), .b(t_12653), .o(t_13175), .cout(t_13176));
half_adder u0_4723(.a(t_12654), .b(t_12656), .o(t_13177), .cout(t_13178));
half_adder u0_4724(.a(t_12657), .b(t_12659), .o(t_13179), .cout(t_13180));
half_adder u0_4725(.a(t_12660), .b(t_12662), .o(t_13181), .cout(t_13182));
compressor_3_2 u1_4726(.a(t_12663), .b(t_12665), .cin(t_11897), .o(t_13183), .cout(t_13184));
compressor_3_2 u1_4727(.a(t_12666), .b(t_12668), .cin(t_11903), .o(t_13185), .cout(t_13186));
half_adder u0_4728(.a(t_12669), .b(t_12671), .o(t_13187), .cout(t_13188));
half_adder u0_4729(.a(t_12672), .b(t_12674), .o(t_13189), .cout(t_13190));
compressor_3_2 u1_4730(.a(t_12675), .b(t_12677), .cin(t_11921), .o(t_13191), .cout(t_13192));
half_adder u0_4731(.a(t_12678), .b(t_12680), .o(t_13193), .cout(t_13194));
compressor_3_2 u1_4732(.a(t_12681), .b(t_12683), .cin(t_11933), .o(t_13195), .cout(t_13196));
half_adder u0_4733(.a(t_12684), .b(t_12686), .o(t_13197), .cout(t_13198));
half_adder u0_4734(.a(t_12687), .b(t_12689), .o(t_13199), .cout(t_13200));
half_adder u0_4735(.a(t_12690), .b(t_12692), .o(t_13201), .cout(t_13202));
half_adder u0_4736(.a(t_12693), .b(t_12695), .o(t_13203), .cout(t_13204));
compressor_3_2 u1_4737(.a(t_12696), .b(t_12698), .cin(t_11963), .o(t_13205), .cout(t_13206));
compressor_3_2 u1_4738(.a(t_12699), .b(t_12701), .cin(t_11969), .o(t_13207), .cout(t_13208));
half_adder u0_4739(.a(t_12702), .b(t_12704), .o(t_13209), .cout(t_13210));
half_adder u0_4740(.a(t_12705), .b(t_12707), .o(t_13211), .cout(t_13212));
half_adder u0_4741(.a(t_12708), .b(t_12710), .o(t_13213), .cout(t_13214));
half_adder u0_4742(.a(t_12711), .b(t_12713), .o(t_13215), .cout(t_13216));
half_adder u0_4743(.a(t_12714), .b(t_12716), .o(t_13217), .cout(t_13218));
half_adder u0_4744(.a(t_12717), .b(t_12719), .o(t_13219), .cout(t_13220));
half_adder u0_4745(.a(t_12720), .b(t_12722), .o(t_13221), .cout(t_13222));
half_adder u0_4746(.a(t_12723), .b(t_12725), .o(t_13223), .cout(t_13224));
compressor_3_2 u1_4747(.a(t_12726), .b(t_12728), .cin(t_12022), .o(t_13225), .cout(t_13226));
compressor_3_2 u1_4748(.a(t_12729), .b(t_12731), .cin(t_12025), .o(t_13227), .cout(t_13228));
half_adder u0_4749(.a(t_12732), .b(t_12733), .o(t_13229), .cout(t_13230));
half_adder u0_4750(.a(t_12734), .b(t_12736), .o(t_13231), .cout(t_13232));
half_adder u0_4751(.a(t_12737), .b(t_12739), .o(t_13233), .cout(t_13234));
half_adder u0_4752(.a(t_12740), .b(t_12742), .o(t_13235), .cout(t_13236));
half_adder u0_4753(.a(t_12743), .b(t_12745), .o(t_13237), .cout(t_13238));
half_adder u0_4754(.a(t_12746), .b(t_12748), .o(t_13239), .cout(t_13240));
half_adder u0_4755(.a(t_12749), .b(t_12751), .o(t_13241), .cout(t_13242));
half_adder u0_4756(.a(t_12752), .b(t_12754), .o(t_13243), .cout(t_13244));
half_adder u0_4757(.a(t_12755), .b(t_12757), .o(t_13245), .cout(t_13246));
half_adder u0_4758(.a(t_12758), .b(t_12760), .o(t_13247), .cout(t_13248));
half_adder u0_4759(.a(t_12761), .b(t_12763), .o(t_13249), .cout(t_13250));
half_adder u0_4760(.a(t_12764), .b(t_12766), .o(t_13251), .cout(t_13252));
half_adder u0_4761(.a(t_12767), .b(t_12769), .o(t_13253), .cout(t_13254));
half_adder u0_4762(.a(t_12770), .b(t_12772), .o(t_13255), .cout(t_13256));
half_adder u0_4763(.a(t_12773), .b(t_12775), .o(t_13257), .cout(t_13258));
half_adder u0_4764(.a(t_12776), .b(t_12778), .o(t_13259), .cout(t_13260));
compressor_3_2 u1_4765(.a(t_12779), .b(t_12781), .cin(t_12111), .o(t_13261), .cout(t_13262));
half_adder u0_4766(.a(t_12782), .b(t_12783), .o(t_13263), .cout(t_13264));
half_adder u0_4767(.a(t_12784), .b(t_12785), .o(t_13265), .cout(t_13266));
half_adder u0_4768(.a(t_12786), .b(t_12787), .o(t_13267), .cout(t_13268));
compressor_3_2 u1_4769(.a(t_12790), .b(t_12792), .cin(t_12136), .o(t_13269), .cout(t_13270));
compressor_3_2 u1_4770(.a(t_12793), .b(t_12794), .cin(t_12141), .o(t_13271), .cout(t_13272));
half_adder u0_4771(.a(t_12795), .b(t_12796), .o(t_13273), .cout(t_13274));
half_adder u0_4772(.a(t_12797), .b(t_12798), .o(t_13275), .cout(t_13276));
half_adder u0_4773(.a(t_12799), .b(t_12800), .o(t_13277), .cout(t_13278));
half_adder u0_4774(.a(t_12801), .b(t_12802), .o(t_13279), .cout(t_13280));
half_adder u0_4775(.a(t_12803), .b(t_12804), .o(t_13281), .cout(t_13282));
half_adder u0_4776(.a(t_12805), .b(t_12806), .o(t_13283), .cout(t_13284));
half_adder u0_4777(.a(t_12807), .b(t_12808), .o(t_13285), .cout(t_13286));
half_adder u0_4778(.a(t_12809), .b(t_12810), .o(t_13287), .cout(t_13288));
half_adder u0_4779(.a(t_12811), .b(t_12812), .o(t_13289), .cout(t_13290));
half_adder u0_4780(.a(t_12813), .b(t_12814), .o(t_13291), .cout(t_13292));
half_adder u0_4781(.a(t_12815), .b(t_12816), .o(t_13293), .cout(t_13294));
half_adder u0_4782(.a(t_12817), .b(t_12818), .o(t_13295), .cout(t_13296));
half_adder u0_4783(.a(t_12819), .b(t_12820), .o(t_13297), .cout(t_13298));
half_adder u0_4784(.a(t_12821), .b(t_12822), .o(t_13299), .cout(t_13300));
half_adder u0_4785(.a(t_12823), .b(t_12824), .o(t_13301), .cout(t_13302));
half_adder u0_4786(.a(t_12825), .b(t_12826), .o(t_13303), .cout(t_13304));
half_adder u0_4787(.a(t_12827), .b(t_12828), .o(t_13305), .cout(t_13306));
half_adder u0_4788(.a(t_12829), .b(t_12830), .o(t_13307), .cout(t_13308));
half_adder u0_4789(.a(t_12831), .b(t_12832), .o(t_13309), .cout(t_13310));
half_adder u0_4790(.a(t_12833), .b(t_12834), .o(t_13311), .cout(t_13312));
half_adder u0_4791(.a(t_12835), .b(t_12836), .o(t_13313), .cout(t_13314));
half_adder u0_4792(.a(t_12837), .b(t_12838), .o(t_13315), .cout(t_13316));
half_adder u0_4793(.a(t_12839), .b(t_12840), .o(t_13317), .cout(t_13318));
half_adder u0_4794(.a(t_12841), .b(t_12842), .o(t_13319), .cout(t_13320));
half_adder u0_4795(.a(t_12843), .b(t_12844), .o(t_13321), .cout(t_13322));
half_adder u0_4796(.a(t_12845), .b(t_12846), .o(t_13323), .cout(t_13324));
half_adder u0_4797(.a(t_12847), .b(t_12848), .o(t_13325), .cout(t_13326));
half_adder u0_4798(.a(t_12849), .b(t_12850), .o(t_13327), .cout(t_13328));
half_adder u0_4799(.a(t_12851), .b(t_12852), .o(t_13329), .cout(t_13330));
half_adder u0_4800(.a(t_12853), .b(t_12854), .o(t_13331), .cout(t_13332));
half_adder u0_4801(.a(t_12855), .b(t_12856), .o(t_13333), .cout(t_13334));
half_adder u0_4802(.a(t_12857), .b(t_12858), .o(t_13335), .cout(t_13336));
half_adder u0_4803(.a(t_12859), .b(t_12860), .o(t_13337), .cout(t_13338));
half_adder u0_4804(.a(t_12861), .b(t_12862), .o(t_13339), .cout(t_13340));
half_adder u0_4805(.a(t_12863), .b(t_12864), .o(t_13341), .cout(t_13342));
half_adder u0_4806(.a(t_12865), .b(t_12866), .o(t_13343), .cout(t_13344));
half_adder u0_4807(.a(t_12867), .b(t_12868), .o(t_13345), .cout(t_13346));
half_adder u0_4808(.a(t_12869), .b(t_12870), .o(t_13347), .cout(t_13348));
half_adder u0_4809(.a(t_12871), .b(t_12872), .o(t_13349), .cout(t_13350));
half_adder u0_4810(.a(t_12873), .b(t_12874), .o(t_13351), .cout(t_13352));
half_adder u0_4811(.a(t_12875), .b(t_12876), .o(t_13353), .cout(t_13354));
half_adder u0_4812(.a(t_12877), .b(t_12878), .o(t_13355), .cout(t_13356));
half_adder u0_4813(.a(t_12879), .b(t_12880), .o(t_13357), .cout(t_13358));
half_adder u0_4814(.a(t_12881), .b(t_12882), .o(t_13359), .cout(t_13360));
half_adder u0_4815(.a(t_12883), .b(t_12884), .o(t_13361), .cout(t_13362));
half_adder u0_4816(.a(t_12885), .b(t_12886), .o(t_13363), .cout(t_13364));
half_adder u0_4817(.a(t_12887), .b(t_12888), .o(t_13365), .cout(t_13366));
half_adder u0_4818(.a(t_12889), .b(t_12890), .o(t_13367), .cout(t_13368));
half_adder u0_4819(.a(t_12891), .b(t_12892), .o(t_13369), .cout(t_13370));
half_adder u0_4820(.a(t_12893), .b(t_12894), .o(t_13371), .cout(t_13372));
half_adder u0_4821(.a(t_12895), .b(t_12896), .o(t_13373), .cout(t_13374));
half_adder u0_4822(.a(t_12897), .b(t_12898), .o(t_13375), .cout(t_13376));
half_adder u0_4823(.a(t_12899), .b(t_12900), .o(t_13377), .cout(t_13378));
half_adder u0_4824(.a(t_12901), .b(t_12902), .o(t_13379), .cout(t_13380));
half_adder u0_4825(.a(t_12903), .b(t_12904), .o(t_13381), .cout(t_13382));
half_adder u0_4826(.a(t_12905), .b(t_12906), .o(t_13383), .cout(t_13384));
half_adder u0_4827(.a(t_12907), .b(t_12908), .o(t_13385), .cout(t_13386));
half_adder u0_4828(.a(t_12909), .b(t_12910), .o(t_13387), .cout(t_13388));
half_adder u0_4829(.a(t_12911), .b(t_12912), .o(t_13389), .cout(t_13390));
half_adder u0_4830(.a(t_12913), .b(t_12914), .o(t_13391), .cout(t_13392));
half_adder u0_4831(.a(t_12915), .b(t_12916), .o(t_13393), .cout(t_13394));
half_adder u0_4832(.a(t_12917), .b(t_12918), .o(t_13395), .cout(t_13396));
half_adder u0_4833(.a(t_12919), .b(t_12920), .o(t_13397), .cout(t_13398));
half_adder u0_4834(.a(t_12921), .b(t_12922), .o(t_13399), .cout(t_13400));
half_adder u0_4835(.a(t_12923), .b(t_12924), .o(t_13401), .cout(t_13402));
half_adder u0_4836(.a(t_12925), .b(t_12926), .o(t_13403), .cout(t_13404));
half_adder u0_4837(.a(t_12927), .b(t_12928), .o(t_13405), .cout(t_13406));
half_adder u0_4838(.a(t_12929), .b(t_12930), .o(t_13407), .cout(t_13408));
half_adder u0_4839(.a(t_12931), .b(t_12932), .o(t_13409), .cout(t_13410));
half_adder u0_4840(.a(t_12933), .b(t_12934), .o(t_13411), .cout(t_13412));
half_adder u0_4841(.a(t_12935), .b(t_12936), .o(t_13413), .cout(t_13414));
half_adder u0_4842(.a(t_12937), .b(t_12938), .o(t_13415), .cout(t_13416));
half_adder u0_4843(.a(t_12939), .b(t_12940), .o(t_13417), .cout(t_13418));
half_adder u0_4844(.a(t_12941), .b(t_12942), .o(t_13419), .cout(t_13420));
half_adder u0_4845(.a(t_12943), .b(t_12944), .o(t_13421), .cout(t_13422));
half_adder u0_4846(.a(t_12945), .b(t_12946), .o(t_13423), .cout(t_13424));
half_adder u0_4847(.a(t_12947), .b(t_12948), .o(t_13425), .cout(t_13426));
half_adder u0_4848(.a(t_12949), .b(t_12950), .o(t_13427), .cout(t_13428));
half_adder u0_4849(.a(t_12951), .b(t_12952), .o(t_13429), .cout(t_13430));
half_adder u0_4850(.a(t_12953), .b(t_12954), .o(t_13431), .cout(t_13432));
half_adder u0_4851(.a(t_12955), .b(t_12956), .o(t_13433), .cout(t_13434));
half_adder u0_4852(.a(t_12957), .b(t_12958), .o(t_13435), .cout());

/* Output nets Compression result */
assign compress_a = {
 t_13435, t_13433, t_13431, t_13429,
 t_13427, t_13425, t_13423, t_13421,
 t_13419, t_13417, t_13415, t_13413,
 t_13411, t_13409, t_13407, t_13405,
 t_13403, t_13401, t_13399, t_13397,
 t_13395, t_13393, t_13391, t_13389,
 t_13387, t_13385, t_13383, t_13381,
 t_13379, t_13377, t_13375, t_13373,
 t_13371, t_13369, t_13367, t_13365,
 t_13363, t_13361, t_13359, t_13357,
 t_13355, t_13353, t_13351, t_13349,
 t_13347, t_13345, t_13343, t_13341,
 t_13339, t_13337, t_13335, t_13333,
 t_13331, t_13329, t_13327, t_13325,
 t_13323, t_13321, t_13319, t_13317,
 t_13315, t_13313, t_13311, t_13309,
 t_13307, t_13305, t_13303, t_13301,
 t_13299, t_13297, t_13295, t_13293,
 t_13291, t_13289, t_13287, t_13285,
 t_13283, t_13281, t_13279, t_13277,
 t_13275, t_13273, t_13271, t_13269,
 t_12789, t_13267, t_13265, t_13263,
 t_13261, t_13259, t_13257, t_13255,
 t_13253, t_13251, t_13249, t_13247,
 t_13245, t_13243, t_13241, t_13239,
 t_13237, t_13235, t_13233, t_13231,
 t_13229, t_13227, t_13225, t_13223,
 t_13221, t_13219, t_13217, t_13215,
 t_13213, t_13211, t_13209, t_13207,
 t_13205, t_13203, t_13201, t_13199,
 t_13197, t_13195, t_13193, t_13191,
 t_13189, t_13187, t_13185, t_13183,
 t_13181, t_13179, t_13177, t_13175,
 t_13173, t_13171, t_13169, t_13167,
 t_13165, t_13163, t_13161, t_13159,
 t_13157, t_12624, t_13155, t_13153,
 t_13151, t_13149, t_13147, t_13145,
 t_13143, t_13141, t_13139, t_13137,
 t_13135, t_13133, t_13131, t_13129,
 t_13127, t_13125, t_13123, t_12573,
 t_13121, t_13119, t_13117, t_13115,
 t_13113, t_12560, t_13111, t_13109,
 t_13107, t_12551, t_13105, t_13103,
 t_13101, t_13099, t_13097, t_13095,
 t_13093, t_13091, t_13089, t_13087,
 t_13085, t_13083, t_13081, t_13079,
 t_13077, t_13075, t_13073, t_13071,
 t_13069, t_13067, t_13065, t_13063,
 t_13061, t_13059, t_13057, t_13055,
 t_13053, t_13051, t_13049, t_13047,
 t_13045, t_13043, t_13041, t_13039,
 t_13037, t_13035, t_12477, t_13033,
 t_13031, t_13029, t_13027, t_12469,
 t_13025, t_13023, t_13021, t_13019,
 t_13017, t_13015, t_13013, t_13011,
 t_13009, t_13007, t_13005, t_13003,
 t_13001, t_12999, t_12997, t_12995,
 t_12993, t_12435, t_12991, t_12989,
 t_12431, t_12987, t_12985, t_12983,
 t_12981, t_12979, t_12977, t_12975,
 t_12973, t_12971, t_12413, t_12969,
 t_12967, t_12965, t_12963, t_12405,
 t_12961, t_12403, t_12959, t_12401,
 t_11460,  t_9728,  t_6441,     t_0
};
assign compress_b = {
 t_13434, t_13432, t_13430, t_13428,
 t_13426, t_13424, t_13422, t_13420,
 t_13418, t_13416, t_13414, t_13412,
 t_13410, t_13408, t_13406, t_13404,
 t_13402, t_13400, t_13398, t_13396,
 t_13394, t_13392, t_13390, t_13388,
 t_13386, t_13384, t_13382, t_13380,
 t_13378, t_13376, t_13374, t_13372,
 t_13370, t_13368, t_13366, t_13364,
 t_13362, t_13360, t_13358, t_13356,
 t_13354, t_13352, t_13350, t_13348,
 t_13346, t_13344, t_13342, t_13340,
 t_13338, t_13336, t_13334, t_13332,
 t_13330, t_13328, t_13326, t_13324,
 t_13322, t_13320, t_13318, t_13316,
 t_13314, t_13312, t_13310, t_13308,
 t_13306, t_13304, t_13302, t_13300,
 t_13298, t_13296, t_13294, t_13292,
 t_13290, t_13288, t_13286, t_13284,
 t_13282, t_13280, t_13278, t_13276,
 t_13274, t_13272, t_13270,    1'b0,
 t_13268, t_13266, t_13264, t_13262,
 t_13260, t_13258, t_13256, t_13254,
 t_13252, t_13250, t_13248, t_13246,
 t_13244, t_13242, t_13240, t_13238,
 t_13236, t_13234, t_13232, t_13230,
 t_13228, t_13226, t_13224, t_13222,
 t_13220, t_13218, t_13216, t_13214,
 t_13212, t_13210, t_13208, t_13206,
 t_13204, t_13202, t_13200, t_13198,
 t_13196, t_13194, t_13192, t_13190,
 t_13188, t_13186, t_13184, t_13182,
 t_13180, t_13178, t_13176, t_13174,
 t_13172, t_13170, t_13168, t_13166,
 t_13164, t_13162, t_13160, t_13158,
    1'b0, t_13156, t_13154, t_13152,
 t_13150, t_13148, t_13146, t_13144,
 t_13142, t_13140, t_13138, t_13136,
 t_13134, t_13132, t_13130, t_13128,
 t_13126, t_13124,    1'b0, t_13122,
 t_13120, t_13118, t_13116, t_13114,
    1'b0, t_13112, t_13110, t_13108,
    1'b0, t_13106, t_13104, t_13102,
 t_13100, t_13098, t_13096, t_13094,
 t_13092, t_13090, t_13088, t_13086,
 t_13084, t_13082, t_13080, t_13078,
 t_13076, t_13074, t_13072, t_13070,
 t_13068, t_13066, t_13064, t_13062,
 t_13060, t_13058, t_13056, t_13054,
 t_13052, t_13050, t_13048, t_13046,
 t_13044, t_13042, t_13040, t_13038,
 t_13036,    1'b0, t_13034, t_13032,
 t_13030, t_13028,    1'b0, t_13026,
 t_13024, t_13022, t_13020, t_13018,
 t_13016, t_13014, t_13012, t_13010,
 t_13008, t_13006, t_13004, t_13002,
 t_13000, t_12998, t_12996, t_12994,
    1'b0, t_12992, t_12990,    1'b0,
 t_12988, t_12986, t_12984, t_12982,
 t_12980, t_12978, t_12976, t_12974,
 t_12972,    1'b0, t_12970, t_12968,
 t_12966, t_12964,    1'b0, t_12962,
    1'b0, t_12960,    1'b0,    1'b0,
    1'b0,    1'b0,    1'b0,    1'b0
};

endmodule

/********************************************************************************/

module booth_coder(
//inputs
	sign,
	a,
	b,
//outputs
	partial_products,
	carry
);

parameter width = 8;

input wire sign;
input wire [width-1:0] a;
input wire [width-1:0] b;
output wire [(width+2)*(width/2+1)-1:0] partial_products;
output reg [width/2-1:0] carry;

reg [(width+2)*(width/2)-1:0] codingdata;
wire [width:0] b_ = {sign&b[width-1], b};
wire [width:0] a_temp = {a, 1'b0};

generate
	genvar i;
	for (i=0; i<width; i=i+2)
	begin: encoder
		always @ (*)
		begin
			case (a_temp[i+2:i])
			3'b0, 3'd7: begin
				codingdata[`INDEX] = {1'b1, {(width+1){1'b0}}};
				carry[i/2] = 1'b0;
			end
			3'd1, 3'd2: begin
				codingdata[`INDEX] = {~b_[width], b_};
				carry[i/2] = 1'b0;
			end
			3'd3: begin
				codingdata[`INDEX] = {~b_[width], b, 1'b0};
				carry[i/2] = 1'b0;
			end
			3'd4: begin
				codingdata[`INDEX] = {b_[width], ~b, 1'b1};
				carry[i/2] = 1'b1;
			end
			3'd5, 3'd6: begin
				codingdata[`INDEX] = {b_[width], ~b_};
				carry[i/2] = 1'b1;
			end
			default: begin
				codingdata[`INDEX] = {(width+2){1'b0}};
				carry[i/2] = 1'b0;
			end
			endcase
		end
	end
endgenerate

function [255:0] sign_sum(input integer n);
integer i;
begin
	for (sign_sum=0, i=0; i<n; i=i+2)
		sign_sum = sign_sum + ({256{1'b1}} << (n-i-2));
	sign_sum = sign_sum << 3;
end
endfunction

wire [width+1:0] signsum = sign_sum(width);
wire [width-1:0] unsign_correct = {width{ a[width-1]&(~sign) }} & b;
wire [width+1:0] extra_product = {signsum[width+1:2]+unsign_correct, signsum[1:0]};

assign partial_products = {extra_product, codingdata};

endmodule

module multer(
//inputs
    sign,
    A,
    B,
//outputs
    P
);

parameter width = 8;

input wire sign;
input wire [width-1:0] A;
input wire [width-1:0] B;
output wire [2*width-1:0] P;

wire [(width+2)*(width/2+1)-1:0] partial_products;
wire [width/2-1:0] carry;
wire [2*width-1:0] compress_a;
wire [2*width-1:0] compress_b;

booth_coder encoder(.sign(sign), .a(A), .b(B), .partial_products(partial_products), .carry(carry));
defparam
    encoder.width=width;

generate
	case (width)
		32 : _32_wallace_tree compressor(.partial_products(partial_products), .carry(carry), .compress_a(compress_a), .compress_b(compress_b));
		64 : _64_wallace_tree compressor(.partial_products(partial_products), .carry(carry), .compress_a(compress_a), .compress_b(compress_b));
		128: _128_wallace_tree compressor(.partial_products(partial_products), .carry(carry), .compress_a(compress_a), .compress_b(compress_b));
		default: _32_wallace_tree compressor(.partial_products(partial_products), .carry(carry), .compress_a(compress_a), .compress_b(compress_b));
	endcase
endgenerate

assign P = compress_a + compress_b;

endmodule

`undef INDEX
