`timescale 1ns / 1ps
`define INDEX (width+2)*(i/2+1)-1:(width+2)*i/2

module half_adder(
//inputs
	a,
	b,
//outputs
	o,
	cout
);

input wire a;
input wire b;
output wire o;
output wire cout;

`ifdef GSCL45NM
HAX1 HALFADD(.A(a),.B(b),.YS(o),.YC(cout));
`else
assign o = a^b;
assign cout = a&b;
`endif

endmodule

module compressor_3_2(
//inputs
	a,
	b,
	cin,
//outputs
	o,
	cout
);
input wire a;
input wire b;
input wire cin;
output wire o;
output wire cout;

`ifdef GSCL45NM
FAX1 FULLADD(.A(a),.B(b),.C(cin),.YS(o),.YC(cout));
`else
wire s = a^b;
wire g = a&b;

assign o = s^cin;
assign cout = s ? cin : g;
`endif

endmodule

module compressor_4_2(
//inputs
	a,
	b,
	c,
	d,
	cin,
//outputs
	o,
	co,
	cout
);

input wire a;
input wire b;
input wire c;
input wire d;
input wire cin;
output wire o;
output wire co;
output wire cout;
`ifdef FPGA_VERSION
wire carry;

compressor_3_2 FULLADD1(a,b,c,carry,cout);
compressor_3_2 FULLADD2(carry,d,cin,o,co);
`elsif GSCL45NM
wire carry;

FAX1 FULLADD1(.A(a),.B(b),.C(c),.YS(carry),.YC(cout));
FAX1 FULLADD2(.A(carry),.B(d),.C(cin),.YS(o),.YC(co));
`else
wire tmp1, tmp2, tmp3, tmp4, tmp5, tmp6;

assign tmp1 = ~(a&b);
assign tmp2 = ~(c&d);
assign tmp3 = ~((a|b)&tmp1);
assign tmp4 = ~((c|d)&tmp2);
assign tmp5 = ~((tmp1|tmp2)&(tmp3|tmp4));
assign tmp6 = tmp3^tmp4;
assign cout = ~(tmp1&tmp2);
assign co = tmp5|(tmp6&cin);
assign o = tmp6^cin;
`endif

endmodule

/********************************************************************************/

module _32_wallace_tree(
//inputs
	partial_products,
	carry,
//outputs
	compress_a,
	compress_b
);

localparam width = 32;

input wire [(width+2)*(width/2+1)-1:0] partial_products;
input wire [width/2-1:0] carry;
output wire [2*width-1:0] compress_a;
output wire [2*width-1:0] compress_b;

/* Input nets */
wire  s_0_0,  s_0_1,  s_1_0,  s_2_0,  s_2_1,  s_2_2;  
wire  s_3_0,  s_3_1,  s_4_0,  s_4_1,  s_4_2,  s_4_3;  
wire  s_5_0,  s_5_1,  s_5_2,  s_6_0,  s_6_1,  s_6_2;  
wire  s_6_3,  s_6_4,  s_7_0,  s_7_1,  s_7_2,  s_7_3;  
wire  s_8_0,  s_8_1,  s_8_2,  s_8_3,  s_8_4,  s_8_5;  
wire  s_9_0,  s_9_1,  s_9_2,  s_9_3,  s_9_4, s_10_0;  
wire s_10_1, s_10_2, s_10_3, s_10_4, s_10_5, s_10_6;  
wire s_11_0, s_11_1, s_11_2, s_11_3, s_11_4, s_11_5;  
wire s_12_0, s_12_1, s_12_2, s_12_3, s_12_4, s_12_5;  
wire s_12_6, s_12_7, s_13_0, s_13_1, s_13_2, s_13_3;  
wire s_13_4, s_13_5, s_13_6, s_14_0, s_14_1, s_14_2;  
wire s_14_3, s_14_4, s_14_5, s_14_6, s_14_7, s_14_8;  
wire s_15_0, s_15_1, s_15_2, s_15_3, s_15_4, s_15_5;  
wire s_15_6, s_15_7, s_16_0, s_16_1, s_16_2, s_16_3;  
wire s_16_4, s_16_5, s_16_6, s_16_7, s_16_8, s_16_9;  
wire s_17_0, s_17_1, s_17_2, s_17_3, s_17_4, s_17_5;  
wire s_17_6, s_17_7, s_17_8, s_18_0, s_18_1, s_18_2;  
wire s_18_3, s_18_4, s_18_5, s_18_6, s_18_7, s_18_8;  
wire s_18_9, s_18_10, s_19_0, s_19_1, s_19_2, s_19_3;  
wire s_19_4, s_19_5, s_19_6, s_19_7, s_19_8, s_19_9;  
wire s_20_0, s_20_1, s_20_2, s_20_3, s_20_4, s_20_5;  
wire s_20_6, s_20_7, s_20_8, s_20_9, s_20_10, s_20_11;  
wire s_21_0, s_21_1, s_21_2, s_21_3, s_21_4, s_21_5;  
wire s_21_6, s_21_7, s_21_8, s_21_9, s_21_10, s_22_0;  
wire s_22_1, s_22_2, s_22_3, s_22_4, s_22_5, s_22_6;  
wire s_22_7, s_22_8, s_22_9, s_22_10, s_22_11, s_22_12;  
wire s_23_0, s_23_1, s_23_2, s_23_3, s_23_4, s_23_5;  
wire s_23_6, s_23_7, s_23_8, s_23_9, s_23_10, s_23_11;  
wire s_24_0, s_24_1, s_24_2, s_24_3, s_24_4, s_24_5;  
wire s_24_6, s_24_7, s_24_8, s_24_9, s_24_10, s_24_11;  
wire s_24_12, s_24_13, s_25_0, s_25_1, s_25_2, s_25_3;  
wire s_25_4, s_25_5, s_25_6, s_25_7, s_25_8, s_25_9;  
wire s_25_10, s_25_11, s_25_12, s_26_0, s_26_1, s_26_2;  
wire s_26_3, s_26_4, s_26_5, s_26_6, s_26_7, s_26_8;  
wire s_26_9, s_26_10, s_26_11, s_26_12, s_26_13, s_26_14;  
wire s_27_0, s_27_1, s_27_2, s_27_3, s_27_4, s_27_5;  
wire s_27_6, s_27_7, s_27_8, s_27_9, s_27_10, s_27_11;  
wire s_27_12, s_27_13, s_28_0, s_28_1, s_28_2, s_28_3;  
wire s_28_4, s_28_5, s_28_6, s_28_7, s_28_8, s_28_9;  
wire s_28_10, s_28_11, s_28_12, s_28_13, s_28_14, s_28_15;  
wire s_29_0, s_29_1, s_29_2, s_29_3, s_29_4, s_29_5;  
wire s_29_6, s_29_7, s_29_8, s_29_9, s_29_10, s_29_11;  
wire s_29_12, s_29_13, s_29_14, s_30_0, s_30_1, s_30_2;  
wire s_30_3, s_30_4, s_30_5, s_30_6, s_30_7, s_30_8;  
wire s_30_9, s_30_10, s_30_11, s_30_12, s_30_13, s_30_14;  
wire s_30_15, s_30_16, s_31_0, s_31_1, s_31_2, s_31_3;  
wire s_31_4, s_31_5, s_31_6, s_31_7, s_31_8, s_31_9;  
wire s_31_10, s_31_11, s_31_12, s_31_13, s_31_14, s_31_15;  
wire s_32_0, s_32_1, s_32_2, s_32_3, s_32_4, s_32_5;  
wire s_32_6, s_32_7, s_32_8, s_32_9, s_32_10, s_32_11;  
wire s_32_12, s_32_13, s_32_14, s_32_15, s_32_16, s_33_0;  
wire s_33_1, s_33_2, s_33_3, s_33_4, s_33_5, s_33_6;  
wire s_33_7, s_33_8, s_33_9, s_33_10, s_33_11, s_33_12;  
wire s_33_13, s_33_14, s_33_15, s_33_16, s_34_0, s_34_1;  
wire s_34_2, s_34_3, s_34_4, s_34_5, s_34_6, s_34_7;  
wire s_34_8, s_34_9, s_34_10, s_34_11, s_34_12, s_34_13;  
wire s_34_14, s_34_15, s_35_0, s_35_1, s_35_2, s_35_3;  
wire s_35_4, s_35_5, s_35_6, s_35_7, s_35_8, s_35_9;  
wire s_35_10, s_35_11, s_35_12, s_35_13, s_35_14, s_35_15;  
wire s_36_0, s_36_1, s_36_2, s_36_3, s_36_4, s_36_5;  
wire s_36_6, s_36_7, s_36_8, s_36_9, s_36_10, s_36_11;  
wire s_36_12, s_36_13, s_36_14, s_37_0, s_37_1, s_37_2;  
wire s_37_3, s_37_4, s_37_5, s_37_6, s_37_7, s_37_8;  
wire s_37_9, s_37_10, s_37_11, s_37_12, s_37_13, s_37_14;  
wire s_38_0, s_38_1, s_38_2, s_38_3, s_38_4, s_38_5;  
wire s_38_6, s_38_7, s_38_8, s_38_9, s_38_10, s_38_11;  
wire s_38_12, s_38_13, s_39_0, s_39_1, s_39_2, s_39_3;  
wire s_39_4, s_39_5, s_39_6, s_39_7, s_39_8, s_39_9;  
wire s_39_10, s_39_11, s_39_12, s_39_13, s_40_0, s_40_1;  
wire s_40_2, s_40_3, s_40_4, s_40_5, s_40_6, s_40_7;  
wire s_40_8, s_40_9, s_40_10, s_40_11, s_40_12, s_41_0;  
wire s_41_1, s_41_2, s_41_3, s_41_4, s_41_5, s_41_6;  
wire s_41_7, s_41_8, s_41_9, s_41_10, s_41_11, s_41_12;  
wire s_42_0, s_42_1, s_42_2, s_42_3, s_42_4, s_42_5;  
wire s_42_6, s_42_7, s_42_8, s_42_9, s_42_10, s_42_11;  
wire s_43_0, s_43_1, s_43_2, s_43_3, s_43_4, s_43_5;  
wire s_43_6, s_43_7, s_43_8, s_43_9, s_43_10, s_43_11;  
wire s_44_0, s_44_1, s_44_2, s_44_3, s_44_4, s_44_5;  
wire s_44_6, s_44_7, s_44_8, s_44_9, s_44_10, s_45_0;  
wire s_45_1, s_45_2, s_45_3, s_45_4, s_45_5, s_45_6;  
wire s_45_7, s_45_8, s_45_9, s_45_10, s_46_0, s_46_1;  
wire s_46_2, s_46_3, s_46_4, s_46_5, s_46_6, s_46_7;  
wire s_46_8, s_46_9, s_47_0, s_47_1, s_47_2, s_47_3;  
wire s_47_4, s_47_5, s_47_6, s_47_7, s_47_8, s_47_9;  
wire s_48_0, s_48_1, s_48_2, s_48_3, s_48_4, s_48_5;  
wire s_48_6, s_48_7, s_48_8, s_49_0, s_49_1, s_49_2;  
wire s_49_3, s_49_4, s_49_5, s_49_6, s_49_7, s_49_8;  
wire s_50_0, s_50_1, s_50_2, s_50_3, s_50_4, s_50_5;  
wire s_50_6, s_50_7, s_51_0, s_51_1, s_51_2, s_51_3;  
wire s_51_4, s_51_5, s_51_6, s_51_7, s_52_0, s_52_1;  
wire s_52_2, s_52_3, s_52_4, s_52_5, s_52_6, s_53_0;  
wire s_53_1, s_53_2, s_53_3, s_53_4, s_53_5, s_53_6;  
wire s_54_0, s_54_1, s_54_2, s_54_3, s_54_4, s_54_5;  
wire s_55_0, s_55_1, s_55_2, s_55_3, s_55_4, s_55_5;  
wire s_56_0, s_56_1, s_56_2, s_56_3, s_56_4, s_57_0;  
wire s_57_1, s_57_2, s_57_3, s_57_4, s_58_0, s_58_1;  
wire s_58_2, s_58_3, s_59_0, s_59_1, s_59_2, s_59_3;  
wire s_60_0, s_60_1, s_60_2, s_61_0, s_61_1, s_61_2;  
wire s_62_0, s_62_1, s_63_0, s_63_1;  

assign {
 s_30_16,  s_28_15,  s_26_14,  s_24_13,  s_22_12,  s_20_11, 
 s_18_10,   s_16_9,   s_14_8,   s_12_7,   s_10_6,    s_8_5, 
   s_6_4,    s_4_3,    s_2_2,    s_0_1  
} = carry;

assign {
  s_33_0,   s_32_0,   s_31_0,   s_30_0,   s_29_0,   s_28_0, 
  s_27_0,   s_26_0,   s_25_0,   s_24_0,   s_23_0,   s_22_0, 
  s_21_0,   s_20_0,   s_19_0,   s_18_0,   s_17_0,   s_16_0, 
  s_15_0,   s_14_0,   s_13_0,   s_12_0,   s_11_0,   s_10_0, 
   s_9_0,    s_8_0,    s_7_0,    s_6_0,    s_5_0,    s_4_0, 
   s_3_0,    s_2_0,    s_1_0,    s_0_0  
} = partial_products[(width+2)*(0+1)-1:(width+2)*0];

assign {
  s_35_0,   s_34_0,   s_33_1,   s_32_1,   s_31_1,   s_30_1, 
  s_29_1,   s_28_1,   s_27_1,   s_26_1,   s_25_1,   s_24_1, 
  s_23_1,   s_22_1,   s_21_1,   s_20_1,   s_19_1,   s_18_1, 
  s_17_1,   s_16_1,   s_15_1,   s_14_1,   s_13_1,   s_12_1, 
  s_11_1,   s_10_1,    s_9_1,    s_8_1,    s_7_1,    s_6_1, 
   s_5_1,    s_4_1,    s_3_1,    s_2_1  
} = partial_products[(width+2)*(1+1)-1:(width+2)*1];

assign {
  s_37_0,   s_36_0,   s_35_1,   s_34_1,   s_33_2,   s_32_2, 
  s_31_2,   s_30_2,   s_29_2,   s_28_2,   s_27_2,   s_26_2, 
  s_25_2,   s_24_2,   s_23_2,   s_22_2,   s_21_2,   s_20_2, 
  s_19_2,   s_18_2,   s_17_2,   s_16_2,   s_15_2,   s_14_2, 
  s_13_2,   s_12_2,   s_11_2,   s_10_2,    s_9_2,    s_8_2, 
   s_7_2,    s_6_2,    s_5_2,    s_4_2  
} = partial_products[(width+2)*(2+1)-1:(width+2)*2];

assign {
  s_39_0,   s_38_0,   s_37_1,   s_36_1,   s_35_2,   s_34_2, 
  s_33_3,   s_32_3,   s_31_3,   s_30_3,   s_29_3,   s_28_3, 
  s_27_3,   s_26_3,   s_25_3,   s_24_3,   s_23_3,   s_22_3, 
  s_21_3,   s_20_3,   s_19_3,   s_18_3,   s_17_3,   s_16_3, 
  s_15_3,   s_14_3,   s_13_3,   s_12_3,   s_11_3,   s_10_3, 
   s_9_3,    s_8_3,    s_7_3,    s_6_3  
} = partial_products[(width+2)*(3+1)-1:(width+2)*3];

assign {
  s_41_0,   s_40_0,   s_39_1,   s_38_1,   s_37_2,   s_36_2, 
  s_35_3,   s_34_3,   s_33_4,   s_32_4,   s_31_4,   s_30_4, 
  s_29_4,   s_28_4,   s_27_4,   s_26_4,   s_25_4,   s_24_4, 
  s_23_4,   s_22_4,   s_21_4,   s_20_4,   s_19_4,   s_18_4, 
  s_17_4,   s_16_4,   s_15_4,   s_14_4,   s_13_4,   s_12_4, 
  s_11_4,   s_10_4,    s_9_4,    s_8_4  
} = partial_products[(width+2)*(4+1)-1:(width+2)*4];

assign {
  s_43_0,   s_42_0,   s_41_1,   s_40_1,   s_39_2,   s_38_2, 
  s_37_3,   s_36_3,   s_35_4,   s_34_4,   s_33_5,   s_32_5, 
  s_31_5,   s_30_5,   s_29_5,   s_28_5,   s_27_5,   s_26_5, 
  s_25_5,   s_24_5,   s_23_5,   s_22_5,   s_21_5,   s_20_5, 
  s_19_5,   s_18_5,   s_17_5,   s_16_5,   s_15_5,   s_14_5, 
  s_13_5,   s_12_5,   s_11_5,   s_10_5  
} = partial_products[(width+2)*(5+1)-1:(width+2)*5];

assign {
  s_45_0,   s_44_0,   s_43_1,   s_42_1,   s_41_2,   s_40_2, 
  s_39_3,   s_38_3,   s_37_4,   s_36_4,   s_35_5,   s_34_5, 
  s_33_6,   s_32_6,   s_31_6,   s_30_6,   s_29_6,   s_28_6, 
  s_27_6,   s_26_6,   s_25_6,   s_24_6,   s_23_6,   s_22_6, 
  s_21_6,   s_20_6,   s_19_6,   s_18_6,   s_17_6,   s_16_6, 
  s_15_6,   s_14_6,   s_13_6,   s_12_6  
} = partial_products[(width+2)*(6+1)-1:(width+2)*6];

assign {
  s_47_0,   s_46_0,   s_45_1,   s_44_1,   s_43_2,   s_42_2, 
  s_41_3,   s_40_3,   s_39_4,   s_38_4,   s_37_5,   s_36_5, 
  s_35_6,   s_34_6,   s_33_7,   s_32_7,   s_31_7,   s_30_7, 
  s_29_7,   s_28_7,   s_27_7,   s_26_7,   s_25_7,   s_24_7, 
  s_23_7,   s_22_7,   s_21_7,   s_20_7,   s_19_7,   s_18_7, 
  s_17_7,   s_16_7,   s_15_7,   s_14_7  
} = partial_products[(width+2)*(7+1)-1:(width+2)*7];

assign {
  s_49_0,   s_48_0,   s_47_1,   s_46_1,   s_45_2,   s_44_2, 
  s_43_3,   s_42_3,   s_41_4,   s_40_4,   s_39_5,   s_38_5, 
  s_37_6,   s_36_6,   s_35_7,   s_34_7,   s_33_8,   s_32_8, 
  s_31_8,   s_30_8,   s_29_8,   s_28_8,   s_27_8,   s_26_8, 
  s_25_8,   s_24_8,   s_23_8,   s_22_8,   s_21_8,   s_20_8, 
  s_19_8,   s_18_8,   s_17_8,   s_16_8  
} = partial_products[(width+2)*(8+1)-1:(width+2)*8];

assign {
  s_51_0,   s_50_0,   s_49_1,   s_48_1,   s_47_2,   s_46_2, 
  s_45_3,   s_44_3,   s_43_4,   s_42_4,   s_41_5,   s_40_5, 
  s_39_6,   s_38_6,   s_37_7,   s_36_7,   s_35_8,   s_34_8, 
  s_33_9,   s_32_9,   s_31_9,   s_30_9,   s_29_9,   s_28_9, 
  s_27_9,   s_26_9,   s_25_9,   s_24_9,   s_23_9,   s_22_9, 
  s_21_9,   s_20_9,   s_19_9,   s_18_9  
} = partial_products[(width+2)*(9+1)-1:(width+2)*9];

assign {
  s_53_0,   s_52_0,   s_51_1,   s_50_1,   s_49_2,   s_48_2, 
  s_47_3,   s_46_3,   s_45_4,   s_44_4,   s_43_5,   s_42_5, 
  s_41_6,   s_40_6,   s_39_7,   s_38_7,   s_37_8,   s_36_8, 
  s_35_9,   s_34_9,  s_33_10,  s_32_10,  s_31_10,  s_30_10, 
 s_29_10,  s_28_10,  s_27_10,  s_26_10,  s_25_10,  s_24_10, 
 s_23_10,  s_22_10,  s_21_10,  s_20_10  
} = partial_products[(width+2)*(10+1)-1:(width+2)*10];

assign {
  s_55_0,   s_54_0,   s_53_1,   s_52_1,   s_51_2,   s_50_2, 
  s_49_3,   s_48_3,   s_47_4,   s_46_4,   s_45_5,   s_44_5, 
  s_43_6,   s_42_6,   s_41_7,   s_40_7,   s_39_8,   s_38_8, 
  s_37_9,   s_36_9,  s_35_10,  s_34_10,  s_33_11,  s_32_11, 
 s_31_11,  s_30_11,  s_29_11,  s_28_11,  s_27_11,  s_26_11, 
 s_25_11,  s_24_11,  s_23_11,  s_22_11  
} = partial_products[(width+2)*(11+1)-1:(width+2)*11];

assign {
  s_57_0,   s_56_0,   s_55_1,   s_54_1,   s_53_2,   s_52_2, 
  s_51_3,   s_50_3,   s_49_4,   s_48_4,   s_47_5,   s_46_5, 
  s_45_6,   s_44_6,   s_43_7,   s_42_7,   s_41_8,   s_40_8, 
  s_39_9,   s_38_9,  s_37_10,  s_36_10,  s_35_11,  s_34_11, 
 s_33_12,  s_32_12,  s_31_12,  s_30_12,  s_29_12,  s_28_12, 
 s_27_12,  s_26_12,  s_25_12,  s_24_12  
} = partial_products[(width+2)*(12+1)-1:(width+2)*12];

assign {
  s_59_0,   s_58_0,   s_57_1,   s_56_1,   s_55_2,   s_54_2, 
  s_53_3,   s_52_3,   s_51_4,   s_50_4,   s_49_5,   s_48_5, 
  s_47_6,   s_46_6,   s_45_7,   s_44_7,   s_43_8,   s_42_8, 
  s_41_9,   s_40_9,  s_39_10,  s_38_10,  s_37_11,  s_36_11, 
 s_35_12,  s_34_12,  s_33_13,  s_32_13,  s_31_13,  s_30_13, 
 s_29_13,  s_28_13,  s_27_13,  s_26_13  
} = partial_products[(width+2)*(13+1)-1:(width+2)*13];

assign {
  s_61_0,   s_60_0,   s_59_1,   s_58_1,   s_57_2,   s_56_2, 
  s_55_3,   s_54_3,   s_53_4,   s_52_4,   s_51_5,   s_50_5, 
  s_49_6,   s_48_6,   s_47_7,   s_46_7,   s_45_8,   s_44_8, 
  s_43_9,   s_42_9,  s_41_10,  s_40_10,  s_39_11,  s_38_11, 
 s_37_12,  s_36_12,  s_35_13,  s_34_13,  s_33_14,  s_32_14, 
 s_31_14,  s_30_14,  s_29_14,  s_28_14  
} = partial_products[(width+2)*(14+1)-1:(width+2)*14];

assign {
  s_63_0,   s_62_0,   s_61_1,   s_60_1,   s_59_2,   s_58_2, 
  s_57_3,   s_56_3,   s_55_4,   s_54_4,   s_53_5,   s_52_5, 
  s_51_6,   s_50_6,   s_49_7,   s_48_7,   s_47_8,   s_46_8, 
  s_45_9,   s_44_9,  s_43_10,  s_42_10,  s_41_11,  s_40_11, 
 s_39_12,  s_38_12,  s_37_13,  s_36_13,  s_35_14,  s_34_14, 
 s_33_15,  s_32_15,  s_31_15,  s_30_15  
} = partial_products[(width+2)*(15+1)-1:(width+2)*15];

assign {
  s_63_1,   s_62_1,   s_61_2,   s_60_2,   s_59_3,   s_58_3, 
  s_57_4,   s_56_4,   s_55_5,   s_54_5,   s_53_6,   s_52_6, 
  s_51_7,   s_50_7,   s_49_8,   s_48_8,   s_47_9,   s_46_9, 
 s_45_10,  s_44_10,  s_43_11,  s_42_11,  s_41_12,  s_40_12, 
 s_39_13,  s_38_13,  s_37_14,  s_36_14,  s_35_15,  s_34_15, 
 s_33_16,  s_32_16  
} = partial_products[(width+2)*(width/2+1)-1:(width+2)*width/2+2];

/* u0_1 Output nets */
wire    t_0,   t_1;  
/* u1_2 Output nets */
wire    t_2,   t_3;  
/* u0_3 Output nets */
wire    t_4,   t_5;  
/* u1_4 Output nets */
wire    t_6,   t_7;  
/* u1_5 Output nets */
wire    t_8,   t_9;  
/* u2_6 Output nets */
wire   t_10,  t_11,  t_12;  
/* u2_7 Output nets */
wire   t_13,  t_14,  t_15;  
/* u2_8 Output nets */
wire   t_16,  t_17,  t_18;  
/* u0_9 Output nets */
wire   t_19,  t_20;  
/* u2_10 Output nets */
wire   t_21,  t_22,  t_23;  
/* u2_11 Output nets */
wire   t_24,  t_25,  t_26;  
/* u1_12 Output nets */
wire   t_27,  t_28;  
/* u2_13 Output nets */
wire   t_29,  t_30,  t_31;  
/* u0_14 Output nets */
wire   t_32,  t_33;  
/* u2_15 Output nets */
wire   t_34,  t_35,  t_36;  
/* u1_16 Output nets */
wire   t_37,  t_38;  
/* u2_17 Output nets */
wire   t_39,  t_40,  t_41;  
/* u1_18 Output nets */
wire   t_42,  t_43;  
/* u2_19 Output nets */
wire   t_44,  t_45,  t_46;  
/* u2_20 Output nets */
wire   t_47,  t_48,  t_49;  
/* u2_21 Output nets */
wire   t_50,  t_51,  t_52;  
/* u2_22 Output nets */
wire   t_53,  t_54,  t_55;  
/* u2_23 Output nets */
wire   t_56,  t_57,  t_58;  
/* u2_24 Output nets */
wire   t_59,  t_60,  t_61;  
/* u0_25 Output nets */
wire   t_62,  t_63;  
/* u2_26 Output nets */
wire   t_64,  t_65,  t_66;  
/* u2_27 Output nets */
wire   t_67,  t_68,  t_69;  
/* u2_28 Output nets */
wire   t_70,  t_71,  t_72;  
/* u2_29 Output nets */
wire   t_73,  t_74,  t_75;  
/* u1_30 Output nets */
wire   t_76,  t_77;  
/* u2_31 Output nets */
wire   t_78,  t_79,  t_80;  
/* u2_32 Output nets */
wire   t_81,  t_82,  t_83;  
/* u0_33 Output nets */
wire   t_84,  t_85;  
/* u2_34 Output nets */
wire   t_86,  t_87,  t_88;  
/* u2_35 Output nets */
wire   t_89,  t_90,  t_91;  
/* u1_36 Output nets */
wire   t_92,  t_93;  
/* u2_37 Output nets */
wire   t_94,  t_95,  t_96;  
/* u2_38 Output nets */
wire   t_97,  t_98,  t_99;  
/* u1_39 Output nets */
wire  t_100, t_101;  
/* u2_40 Output nets */
wire  t_102, t_103, t_104;  
/* u2_41 Output nets */
wire  t_105, t_106, t_107;  
/* u2_42 Output nets */
wire  t_108, t_109, t_110;  
/* u2_43 Output nets */
wire  t_111, t_112, t_113;  
/* u2_44 Output nets */
wire  t_114, t_115, t_116;  
/* u2_45 Output nets */
wire  t_117, t_118, t_119;  
/* u2_46 Output nets */
wire  t_120, t_121, t_122;  
/* u2_47 Output nets */
wire  t_123, t_124, t_125;  
/* u2_48 Output nets */
wire  t_126, t_127, t_128;  
/* u0_49 Output nets */
wire  t_129, t_130;  
/* u2_50 Output nets */
wire  t_131, t_132, t_133;  
/* u2_51 Output nets */
wire  t_134, t_135, t_136;  
/* u2_52 Output nets */
wire  t_137, t_138, t_139;  
/* u2_53 Output nets */
wire  t_140, t_141, t_142;  
/* u2_54 Output nets */
wire  t_143, t_144, t_145;  
/* u2_55 Output nets */
wire  t_146, t_147, t_148;  
/* u1_56 Output nets */
wire  t_149, t_150;  
/* u2_57 Output nets */
wire  t_151, t_152, t_153;  
/* u2_58 Output nets */
wire  t_154, t_155, t_156;  
/* u2_59 Output nets */
wire  t_157, t_158, t_159;  
/* u0_60 Output nets */
wire  t_160, t_161;  
/* u2_61 Output nets */
wire  t_162, t_163, t_164;  
/* u2_62 Output nets */
wire  t_165, t_166, t_167;  
/* u2_63 Output nets */
wire  t_168, t_169, t_170;  
/* u1_64 Output nets */
wire  t_171, t_172;  
/* u2_65 Output nets */
wire  t_173, t_174, t_175;  
/* u2_66 Output nets */
wire  t_176, t_177, t_178;  
/* u2_67 Output nets */
wire  t_179, t_180, t_181;  
/* u1_68 Output nets */
wire  t_182, t_183;  
/* u2_69 Output nets */
wire  t_184, t_185, t_186;  
/* u2_70 Output nets */
wire  t_187, t_188, t_189;  
/* u2_71 Output nets */
wire  t_190, t_191, t_192;  
/* u2_72 Output nets */
wire  t_193, t_194, t_195;  
/* u2_73 Output nets */
wire  t_196, t_197, t_198;  
/* u2_74 Output nets */
wire  t_199, t_200, t_201;  
/* u2_75 Output nets */
wire  t_202, t_203, t_204;  
/* u2_76 Output nets */
wire  t_205, t_206, t_207;  
/* u2_77 Output nets */
wire  t_208, t_209, t_210;  
/* u2_78 Output nets */
wire  t_211, t_212, t_213;  
/* u2_79 Output nets */
wire  t_214, t_215, t_216;  
/* u2_80 Output nets */
wire  t_217, t_218, t_219;  
/* u2_81 Output nets */
wire  t_220, t_221, t_222;  
/* u2_82 Output nets */
wire  t_223, t_224, t_225;  
/* u2_83 Output nets */
wire  t_226, t_227, t_228;  
/* u2_84 Output nets */
wire  t_229, t_230, t_231;  
/* u2_85 Output nets */
wire  t_232, t_233, t_234;  
/* u2_86 Output nets */
wire  t_235, t_236, t_237;  
/* u2_87 Output nets */
wire  t_238, t_239, t_240;  
/* u2_88 Output nets */
wire  t_241, t_242, t_243;  
/* u2_89 Output nets */
wire  t_244, t_245, t_246;  
/* u2_90 Output nets */
wire  t_247, t_248, t_249;  
/* u2_91 Output nets */
wire  t_250, t_251, t_252;  
/* u2_92 Output nets */
wire  t_253, t_254, t_255;  
/* u2_93 Output nets */
wire  t_256, t_257, t_258;  
/* u2_94 Output nets */
wire  t_259, t_260, t_261;  
/* u2_95 Output nets */
wire  t_262, t_263, t_264;  
/* u1_96 Output nets */
wire  t_265, t_266;  
/* u2_97 Output nets */
wire  t_267, t_268, t_269;  
/* u2_98 Output nets */
wire  t_270, t_271, t_272;  
/* u2_99 Output nets */
wire  t_273, t_274, t_275;  
/* u1_100 Output nets */
wire  t_276, t_277;  
/* u2_101 Output nets */
wire  t_278, t_279, t_280;  
/* u2_102 Output nets */
wire  t_281, t_282, t_283;  
/* u2_103 Output nets */
wire  t_284, t_285, t_286;  
/* u0_104 Output nets */
wire  t_287, t_288;  
/* u2_105 Output nets */
wire  t_289, t_290, t_291;  
/* u2_106 Output nets */
wire  t_292, t_293, t_294;  
/* u2_107 Output nets */
wire  t_295, t_296, t_297;  
/* u0_108 Output nets */
wire  t_298, t_299;  
/* u2_109 Output nets */
wire  t_300, t_301, t_302;  
/* u2_110 Output nets */
wire  t_303, t_304, t_305;  
/* u2_111 Output nets */
wire  t_306, t_307, t_308;  
/* u2_112 Output nets */
wire  t_309, t_310, t_311;  
/* u2_113 Output nets */
wire  t_312, t_313, t_314;  
/* u2_114 Output nets */
wire  t_315, t_316, t_317;  
/* u2_115 Output nets */
wire  t_318, t_319, t_320;  
/* u2_116 Output nets */
wire  t_321, t_322, t_323;  
/* u2_117 Output nets */
wire  t_324, t_325, t_326;  
/* u2_118 Output nets */
wire  t_327, t_328, t_329;  
/* u2_119 Output nets */
wire  t_330, t_331, t_332;  
/* u2_120 Output nets */
wire  t_333, t_334, t_335;  
/* u2_121 Output nets */
wire  t_336, t_337, t_338;  
/* u2_122 Output nets */
wire  t_339, t_340, t_341;  
/* u1_123 Output nets */
wire  t_342, t_343;  
/* u2_124 Output nets */
wire  t_344, t_345, t_346;  
/* u2_125 Output nets */
wire  t_347, t_348, t_349;  
/* u1_126 Output nets */
wire  t_350, t_351;  
/* u2_127 Output nets */
wire  t_352, t_353, t_354;  
/* u2_128 Output nets */
wire  t_355, t_356, t_357;  
/* u0_129 Output nets */
wire  t_358, t_359;  
/* u2_130 Output nets */
wire  t_360, t_361, t_362;  
/* u2_131 Output nets */
wire  t_363, t_364, t_365;  
/* u0_132 Output nets */
wire  t_366, t_367;  
/* u2_133 Output nets */
wire  t_368, t_369, t_370;  
/* u2_134 Output nets */
wire  t_371, t_372, t_373;  
/* u2_135 Output nets */
wire  t_374, t_375, t_376;  
/* u2_136 Output nets */
wire  t_377, t_378, t_379;  
/* u2_137 Output nets */
wire  t_380, t_381, t_382;  
/* u2_138 Output nets */
wire  t_383, t_384, t_385;  
/* u2_139 Output nets */
wire  t_386, t_387, t_388;  
/* u2_140 Output nets */
wire  t_389, t_390, t_391;  
/* u2_141 Output nets */
wire  t_392, t_393, t_394;  
/* u1_142 Output nets */
wire  t_395, t_396;  
/* u2_143 Output nets */
wire  t_397, t_398, t_399;  
/* u1_144 Output nets */
wire  t_400, t_401;  
/* u2_145 Output nets */
wire  t_402, t_403, t_404;  
/* u0_146 Output nets */
wire  t_405, t_406;  
/* u2_147 Output nets */
wire  t_407, t_408, t_409;  
/* u0_148 Output nets */
wire  t_410, t_411;  
/* u2_149 Output nets */
wire  t_412, t_413, t_414;  
/* u2_150 Output nets */
wire  t_415, t_416, t_417;  
/* u2_151 Output nets */
wire  t_418, t_419, t_420;  
/* u2_152 Output nets */
wire  t_421, t_422, t_423;  
/* u1_153 Output nets */
wire  t_424, t_425;  
/* u1_154 Output nets */
wire  t_426, t_427;  
/* u0_155 Output nets */
wire  t_428, t_429;  
/* u0_156 Output nets */
wire  t_430;  

/* compress stage 1 */
half_adder u0_1(.a(s_0_1), .b(s_0_0), .o(t_0), .cout(t_1)); 
compressor_3_2 u1_2(.a(s_2_2), .b(s_2_1), .cin(s_2_0), .o(t_2), .cout(t_3)); 
half_adder u0_3(.a(s_3_1), .b(s_3_0), .o(t_4), .cout(t_5)); 
compressor_3_2 u1_4(.a(s_4_2), .b(s_4_1), .cin(s_4_0), .o(t_6), .cout(t_7)); 
compressor_3_2 u1_5(.a(s_5_2), .b(s_5_1), .cin(s_5_0), .o(t_8), .cout(t_9)); 
compressor_4_2 u2_6(.a(s_6_4), .b(s_6_3), .c(s_6_2), .d(s_6_1), .cin(s_6_0), .o(t_10), .co(t_11), .cout(t_12)); 
compressor_4_2 u2_7(.a(s_7_3), .b(s_7_2), .c(s_7_1), .d(s_7_0), .cin(t_12), .o(t_13), .co(t_14), .cout(t_15)); 
compressor_4_2 u2_8(.a(s_8_3), .b(s_8_2), .c(s_8_1), .d(s_8_0), .cin(t_15), .o(t_16), .co(t_17), .cout(t_18)); 
half_adder u0_9(.a(s_8_5), .b(s_8_4), .o(t_19), .cout(t_20)); 
compressor_4_2 u2_10(.a(s_9_3), .b(s_9_2), .c(s_9_1), .d(s_9_0), .cin(t_18), .o(t_21), .co(t_22), .cout(t_23)); 
compressor_4_2 u2_11(.a(s_10_3), .b(s_10_2), .c(s_10_1), .d(s_10_0), .cin(t_23), .o(t_24), .co(t_25), .cout(t_26)); 
compressor_3_2 u1_12(.a(s_10_6), .b(s_10_5), .cin(s_10_4), .o(t_27), .cout(t_28)); 
compressor_4_2 u2_13(.a(s_11_3), .b(s_11_2), .c(s_11_1), .d(s_11_0), .cin(t_26), .o(t_29), .co(t_30), .cout(t_31)); 
half_adder u0_14(.a(s_11_5), .b(s_11_4), .o(t_32), .cout(t_33)); 
compressor_4_2 u2_15(.a(s_12_3), .b(s_12_2), .c(s_12_1), .d(s_12_0), .cin(t_31), .o(t_34), .co(t_35), .cout(t_36)); 
compressor_3_2 u1_16(.a(s_12_6), .b(s_12_5), .cin(s_12_4), .o(t_37), .cout(t_38)); 
compressor_4_2 u2_17(.a(s_13_3), .b(s_13_2), .c(s_13_1), .d(s_13_0), .cin(t_36), .o(t_39), .co(t_40), .cout(t_41)); 
compressor_3_2 u1_18(.a(s_13_6), .b(s_13_5), .cin(s_13_4), .o(t_42), .cout(t_43)); 
compressor_4_2 u2_19(.a(s_14_3), .b(s_14_2), .c(s_14_1), .d(s_14_0), .cin(t_41), .o(t_44), .co(t_45), .cout(t_46)); 
compressor_4_2 u2_20(.a(s_14_8), .b(s_14_7), .c(s_14_6), .d(s_14_5), .cin(s_14_4), .o(t_47), .co(t_48), .cout(t_49)); 
compressor_4_2 u2_21(.a(s_15_3), .b(s_15_2), .c(s_15_1), .d(s_15_0), .cin(t_46), .o(t_50), .co(t_51), .cout(t_52)); 
compressor_4_2 u2_22(.a(s_15_7), .b(s_15_6), .c(s_15_5), .d(s_15_4), .cin(t_49), .o(t_53), .co(t_54), .cout(t_55)); 
compressor_4_2 u2_23(.a(s_16_3), .b(s_16_2), .c(s_16_1), .d(s_16_0), .cin(t_52), .o(t_56), .co(t_57), .cout(t_58)); 
compressor_4_2 u2_24(.a(s_16_7), .b(s_16_6), .c(s_16_5), .d(s_16_4), .cin(t_55), .o(t_59), .co(t_60), .cout(t_61)); 
half_adder u0_25(.a(s_16_9), .b(s_16_8), .o(t_62), .cout(t_63)); 
compressor_4_2 u2_26(.a(s_17_3), .b(s_17_2), .c(s_17_1), .d(s_17_0), .cin(t_58), .o(t_64), .co(t_65), .cout(t_66)); 
compressor_4_2 u2_27(.a(s_17_7), .b(s_17_6), .c(s_17_5), .d(s_17_4), .cin(t_61), .o(t_67), .co(t_68), .cout(t_69)); 
compressor_4_2 u2_28(.a(s_18_3), .b(s_18_2), .c(s_18_1), .d(s_18_0), .cin(t_66), .o(t_70), .co(t_71), .cout(t_72)); 
compressor_4_2 u2_29(.a(s_18_7), .b(s_18_6), .c(s_18_5), .d(s_18_4), .cin(t_69), .o(t_73), .co(t_74), .cout(t_75)); 
compressor_3_2 u1_30(.a(s_18_10), .b(s_18_9), .cin(s_18_8), .o(t_76), .cout(t_77)); 
compressor_4_2 u2_31(.a(s_19_3), .b(s_19_2), .c(s_19_1), .d(s_19_0), .cin(t_72), .o(t_78), .co(t_79), .cout(t_80)); 
compressor_4_2 u2_32(.a(s_19_7), .b(s_19_6), .c(s_19_5), .d(s_19_4), .cin(t_75), .o(t_81), .co(t_82), .cout(t_83)); 
half_adder u0_33(.a(s_19_9), .b(s_19_8), .o(t_84), .cout(t_85)); 
compressor_4_2 u2_34(.a(s_20_3), .b(s_20_2), .c(s_20_1), .d(s_20_0), .cin(t_80), .o(t_86), .co(t_87), .cout(t_88)); 
compressor_4_2 u2_35(.a(s_20_7), .b(s_20_6), .c(s_20_5), .d(s_20_4), .cin(t_83), .o(t_89), .co(t_90), .cout(t_91)); 
compressor_3_2 u1_36(.a(s_20_10), .b(s_20_9), .cin(s_20_8), .o(t_92), .cout(t_93)); 
compressor_4_2 u2_37(.a(s_21_3), .b(s_21_2), .c(s_21_1), .d(s_21_0), .cin(t_88), .o(t_94), .co(t_95), .cout(t_96)); 
compressor_4_2 u2_38(.a(s_21_7), .b(s_21_6), .c(s_21_5), .d(s_21_4), .cin(t_91), .o(t_97), .co(t_98), .cout(t_99)); 
compressor_3_2 u1_39(.a(s_21_10), .b(s_21_9), .cin(s_21_8), .o(t_100), .cout(t_101)); 
compressor_4_2 u2_40(.a(s_22_3), .b(s_22_2), .c(s_22_1), .d(s_22_0), .cin(t_96), .o(t_102), .co(t_103), .cout(t_104)); 
compressor_4_2 u2_41(.a(s_22_7), .b(s_22_6), .c(s_22_5), .d(s_22_4), .cin(t_99), .o(t_105), .co(t_106), .cout(t_107)); 
compressor_4_2 u2_42(.a(s_22_12), .b(s_22_11), .c(s_22_10), .d(s_22_9), .cin(s_22_8), .o(t_108), .co(t_109), .cout(t_110)); 
compressor_4_2 u2_43(.a(s_23_3), .b(s_23_2), .c(s_23_1), .d(s_23_0), .cin(t_104), .o(t_111), .co(t_112), .cout(t_113)); 
compressor_4_2 u2_44(.a(s_23_7), .b(s_23_6), .c(s_23_5), .d(s_23_4), .cin(t_107), .o(t_114), .co(t_115), .cout(t_116)); 
compressor_4_2 u2_45(.a(s_23_11), .b(s_23_10), .c(s_23_9), .d(s_23_8), .cin(t_110), .o(t_117), .co(t_118), .cout(t_119)); 
compressor_4_2 u2_46(.a(s_24_3), .b(s_24_2), .c(s_24_1), .d(s_24_0), .cin(t_113), .o(t_120), .co(t_121), .cout(t_122)); 
compressor_4_2 u2_47(.a(s_24_7), .b(s_24_6), .c(s_24_5), .d(s_24_4), .cin(t_116), .o(t_123), .co(t_124), .cout(t_125)); 
compressor_4_2 u2_48(.a(s_24_11), .b(s_24_10), .c(s_24_9), .d(s_24_8), .cin(t_119), .o(t_126), .co(t_127), .cout(t_128)); 
half_adder u0_49(.a(s_24_13), .b(s_24_12), .o(t_129), .cout(t_130)); 
compressor_4_2 u2_50(.a(s_25_3), .b(s_25_2), .c(s_25_1), .d(s_25_0), .cin(t_122), .o(t_131), .co(t_132), .cout(t_133)); 
compressor_4_2 u2_51(.a(s_25_7), .b(s_25_6), .c(s_25_5), .d(s_25_4), .cin(t_125), .o(t_134), .co(t_135), .cout(t_136)); 
compressor_4_2 u2_52(.a(s_25_11), .b(s_25_10), .c(s_25_9), .d(s_25_8), .cin(t_128), .o(t_137), .co(t_138), .cout(t_139)); 
compressor_4_2 u2_53(.a(s_26_3), .b(s_26_2), .c(s_26_1), .d(s_26_0), .cin(t_133), .o(t_140), .co(t_141), .cout(t_142)); 
compressor_4_2 u2_54(.a(s_26_7), .b(s_26_6), .c(s_26_5), .d(s_26_4), .cin(t_136), .o(t_143), .co(t_144), .cout(t_145)); 
compressor_4_2 u2_55(.a(s_26_11), .b(s_26_10), .c(s_26_9), .d(s_26_8), .cin(t_139), .o(t_146), .co(t_147), .cout(t_148)); 
compressor_3_2 u1_56(.a(s_26_14), .b(s_26_13), .cin(s_26_12), .o(t_149), .cout(t_150)); 
compressor_4_2 u2_57(.a(s_27_3), .b(s_27_2), .c(s_27_1), .d(s_27_0), .cin(t_142), .o(t_151), .co(t_152), .cout(t_153)); 
compressor_4_2 u2_58(.a(s_27_7), .b(s_27_6), .c(s_27_5), .d(s_27_4), .cin(t_145), .o(t_154), .co(t_155), .cout(t_156)); 
compressor_4_2 u2_59(.a(s_27_11), .b(s_27_10), .c(s_27_9), .d(s_27_8), .cin(t_148), .o(t_157), .co(t_158), .cout(t_159)); 
half_adder u0_60(.a(s_27_13), .b(s_27_12), .o(t_160), .cout(t_161)); 
compressor_4_2 u2_61(.a(s_28_3), .b(s_28_2), .c(s_28_1), .d(s_28_0), .cin(t_153), .o(t_162), .co(t_163), .cout(t_164)); 
compressor_4_2 u2_62(.a(s_28_7), .b(s_28_6), .c(s_28_5), .d(s_28_4), .cin(t_156), .o(t_165), .co(t_166), .cout(t_167)); 
compressor_4_2 u2_63(.a(s_28_11), .b(s_28_10), .c(s_28_9), .d(s_28_8), .cin(t_159), .o(t_168), .co(t_169), .cout(t_170)); 
compressor_3_2 u1_64(.a(s_28_14), .b(s_28_13), .cin(s_28_12), .o(t_171), .cout(t_172)); 
compressor_4_2 u2_65(.a(s_29_3), .b(s_29_2), .c(s_29_1), .d(s_29_0), .cin(t_164), .o(t_173), .co(t_174), .cout(t_175)); 
compressor_4_2 u2_66(.a(s_29_7), .b(s_29_6), .c(s_29_5), .d(s_29_4), .cin(t_167), .o(t_176), .co(t_177), .cout(t_178)); 
compressor_4_2 u2_67(.a(s_29_11), .b(s_29_10), .c(s_29_9), .d(s_29_8), .cin(t_170), .o(t_179), .co(t_180), .cout(t_181)); 
compressor_3_2 u1_68(.a(s_29_14), .b(s_29_13), .cin(s_29_12), .o(t_182), .cout(t_183)); 
compressor_4_2 u2_69(.a(s_30_3), .b(s_30_2), .c(s_30_1), .d(s_30_0), .cin(t_175), .o(t_184), .co(t_185), .cout(t_186)); 
compressor_4_2 u2_70(.a(s_30_7), .b(s_30_6), .c(s_30_5), .d(s_30_4), .cin(t_178), .o(t_187), .co(t_188), .cout(t_189)); 
compressor_4_2 u2_71(.a(s_30_11), .b(s_30_10), .c(s_30_9), .d(s_30_8), .cin(t_181), .o(t_190), .co(t_191), .cout(t_192)); 
compressor_4_2 u2_72(.a(s_30_16), .b(s_30_15), .c(s_30_14), .d(s_30_13), .cin(s_30_12), .o(t_193), .co(t_194), .cout(t_195)); 
compressor_4_2 u2_73(.a(s_31_3), .b(s_31_2), .c(s_31_1), .d(s_31_0), .cin(t_186), .o(t_196), .co(t_197), .cout(t_198)); 
compressor_4_2 u2_74(.a(s_31_7), .b(s_31_6), .c(s_31_5), .d(s_31_4), .cin(t_189), .o(t_199), .co(t_200), .cout(t_201)); 
compressor_4_2 u2_75(.a(s_31_11), .b(s_31_10), .c(s_31_9), .d(s_31_8), .cin(t_192), .o(t_202), .co(t_203), .cout(t_204)); 
compressor_4_2 u2_76(.a(s_31_15), .b(s_31_14), .c(s_31_13), .d(s_31_12), .cin(t_195), .o(t_205), .co(t_206), .cout(t_207)); 
compressor_4_2 u2_77(.a(s_32_3), .b(s_32_2), .c(s_32_1), .d(s_32_0), .cin(t_198), .o(t_208), .co(t_209), .cout(t_210)); 
compressor_4_2 u2_78(.a(s_32_7), .b(s_32_6), .c(s_32_5), .d(s_32_4), .cin(t_201), .o(t_211), .co(t_212), .cout(t_213)); 
compressor_4_2 u2_79(.a(s_32_11), .b(s_32_10), .c(s_32_9), .d(s_32_8), .cin(t_204), .o(t_214), .co(t_215), .cout(t_216)); 
compressor_4_2 u2_80(.a(s_32_15), .b(s_32_14), .c(s_32_13), .d(s_32_12), .cin(t_207), .o(t_217), .co(t_218), .cout(t_219)); 
compressor_4_2 u2_81(.a(s_33_3), .b(s_33_2), .c(s_33_1), .d(s_33_0), .cin(t_210), .o(t_220), .co(t_221), .cout(t_222)); 
compressor_4_2 u2_82(.a(s_33_7), .b(s_33_6), .c(s_33_5), .d(s_33_4), .cin(t_213), .o(t_223), .co(t_224), .cout(t_225)); 
compressor_4_2 u2_83(.a(s_33_11), .b(s_33_10), .c(s_33_9), .d(s_33_8), .cin(t_216), .o(t_226), .co(t_227), .cout(t_228)); 
compressor_4_2 u2_84(.a(s_33_15), .b(s_33_14), .c(s_33_13), .d(s_33_12), .cin(t_219), .o(t_229), .co(t_230), .cout(t_231)); 
compressor_4_2 u2_85(.a(s_34_3), .b(s_34_2), .c(s_34_1), .d(s_34_0), .cin(t_222), .o(t_232), .co(t_233), .cout(t_234)); 
compressor_4_2 u2_86(.a(s_34_7), .b(s_34_6), .c(s_34_5), .d(s_34_4), .cin(t_225), .o(t_235), .co(t_236), .cout(t_237)); 
compressor_4_2 u2_87(.a(s_34_11), .b(s_34_10), .c(s_34_9), .d(s_34_8), .cin(t_228), .o(t_238), .co(t_239), .cout(t_240)); 
compressor_4_2 u2_88(.a(s_34_15), .b(s_34_14), .c(s_34_13), .d(s_34_12), .cin(t_231), .o(t_241), .co(t_242), .cout(t_243)); 
compressor_4_2 u2_89(.a(s_35_3), .b(s_35_2), .c(s_35_1), .d(s_35_0), .cin(t_234), .o(t_244), .co(t_245), .cout(t_246)); 
compressor_4_2 u2_90(.a(s_35_7), .b(s_35_6), .c(s_35_5), .d(s_35_4), .cin(t_237), .o(t_247), .co(t_248), .cout(t_249)); 
compressor_4_2 u2_91(.a(s_35_11), .b(s_35_10), .c(s_35_9), .d(s_35_8), .cin(t_240), .o(t_250), .co(t_251), .cout(t_252)); 
compressor_4_2 u2_92(.a(s_35_15), .b(s_35_14), .c(s_35_13), .d(s_35_12), .cin(t_243), .o(t_253), .co(t_254), .cout(t_255)); 
compressor_4_2 u2_93(.a(s_36_3), .b(s_36_2), .c(s_36_1), .d(s_36_0), .cin(t_246), .o(t_256), .co(t_257), .cout(t_258)); 
compressor_4_2 u2_94(.a(s_36_7), .b(s_36_6), .c(s_36_5), .d(s_36_4), .cin(t_249), .o(t_259), .co(t_260), .cout(t_261)); 
compressor_4_2 u2_95(.a(s_36_11), .b(s_36_10), .c(s_36_9), .d(s_36_8), .cin(t_252), .o(t_262), .co(t_263), .cout(t_264)); 
compressor_3_2 u1_96(.a(s_36_13), .b(s_36_12), .cin(t_255), .o(t_265), .cout(t_266)); 
compressor_4_2 u2_97(.a(s_37_3), .b(s_37_2), .c(s_37_1), .d(s_37_0), .cin(t_258), .o(t_267), .co(t_268), .cout(t_269)); 
compressor_4_2 u2_98(.a(s_37_7), .b(s_37_6), .c(s_37_5), .d(s_37_4), .cin(t_261), .o(t_270), .co(t_271), .cout(t_272)); 
compressor_4_2 u2_99(.a(s_37_11), .b(s_37_10), .c(s_37_9), .d(s_37_8), .cin(t_264), .o(t_273), .co(t_274), .cout(t_275)); 
compressor_3_2 u1_100(.a(s_37_14), .b(s_37_13), .cin(s_37_12), .o(t_276), .cout(t_277)); 
compressor_4_2 u2_101(.a(s_38_3), .b(s_38_2), .c(s_38_1), .d(s_38_0), .cin(t_269), .o(t_278), .co(t_279), .cout(t_280)); 
compressor_4_2 u2_102(.a(s_38_7), .b(s_38_6), .c(s_38_5), .d(s_38_4), .cin(t_272), .o(t_281), .co(t_282), .cout(t_283)); 
compressor_4_2 u2_103(.a(s_38_11), .b(s_38_10), .c(s_38_9), .d(s_38_8), .cin(t_275), .o(t_284), .co(t_285), .cout(t_286)); 
half_adder u0_104(.a(s_38_13), .b(s_38_12), .o(t_287), .cout(t_288)); 
compressor_4_2 u2_105(.a(s_39_3), .b(s_39_2), .c(s_39_1), .d(s_39_0), .cin(t_280), .o(t_289), .co(t_290), .cout(t_291)); 
compressor_4_2 u2_106(.a(s_39_7), .b(s_39_6), .c(s_39_5), .d(s_39_4), .cin(t_283), .o(t_292), .co(t_293), .cout(t_294)); 
compressor_4_2 u2_107(.a(s_39_11), .b(s_39_10), .c(s_39_9), .d(s_39_8), .cin(t_286), .o(t_295), .co(t_296), .cout(t_297)); 
half_adder u0_108(.a(s_39_13), .b(s_39_12), .o(t_298), .cout(t_299)); 
compressor_4_2 u2_109(.a(s_40_3), .b(s_40_2), .c(s_40_1), .d(s_40_0), .cin(t_291), .o(t_300), .co(t_301), .cout(t_302)); 
compressor_4_2 u2_110(.a(s_40_7), .b(s_40_6), .c(s_40_5), .d(s_40_4), .cin(t_294), .o(t_303), .co(t_304), .cout(t_305)); 
compressor_4_2 u2_111(.a(s_40_11), .b(s_40_10), .c(s_40_9), .d(s_40_8), .cin(t_297), .o(t_306), .co(t_307), .cout(t_308)); 
compressor_4_2 u2_112(.a(s_41_3), .b(s_41_2), .c(s_41_1), .d(s_41_0), .cin(t_302), .o(t_309), .co(t_310), .cout(t_311)); 
compressor_4_2 u2_113(.a(s_41_7), .b(s_41_6), .c(s_41_5), .d(s_41_4), .cin(t_305), .o(t_312), .co(t_313), .cout(t_314)); 
compressor_4_2 u2_114(.a(s_41_11), .b(s_41_10), .c(s_41_9), .d(s_41_8), .cin(t_308), .o(t_315), .co(t_316), .cout(t_317)); 
compressor_4_2 u2_115(.a(s_42_3), .b(s_42_2), .c(s_42_1), .d(s_42_0), .cin(t_311), .o(t_318), .co(t_319), .cout(t_320)); 
compressor_4_2 u2_116(.a(s_42_7), .b(s_42_6), .c(s_42_5), .d(s_42_4), .cin(t_314), .o(t_321), .co(t_322), .cout(t_323)); 
compressor_4_2 u2_117(.a(s_42_11), .b(s_42_10), .c(s_42_9), .d(s_42_8), .cin(t_317), .o(t_324), .co(t_325), .cout(t_326)); 
compressor_4_2 u2_118(.a(s_43_3), .b(s_43_2), .c(s_43_1), .d(s_43_0), .cin(t_320), .o(t_327), .co(t_328), .cout(t_329)); 
compressor_4_2 u2_119(.a(s_43_7), .b(s_43_6), .c(s_43_5), .d(s_43_4), .cin(t_323), .o(t_330), .co(t_331), .cout(t_332)); 
compressor_4_2 u2_120(.a(s_43_11), .b(s_43_10), .c(s_43_9), .d(s_43_8), .cin(t_326), .o(t_333), .co(t_334), .cout(t_335)); 
compressor_4_2 u2_121(.a(s_44_3), .b(s_44_2), .c(s_44_1), .d(s_44_0), .cin(t_329), .o(t_336), .co(t_337), .cout(t_338)); 
compressor_4_2 u2_122(.a(s_44_7), .b(s_44_6), .c(s_44_5), .d(s_44_4), .cin(t_332), .o(t_339), .co(t_340), .cout(t_341)); 
compressor_3_2 u1_123(.a(s_44_9), .b(s_44_8), .cin(t_335), .o(t_342), .cout(t_343)); 
compressor_4_2 u2_124(.a(s_45_3), .b(s_45_2), .c(s_45_1), .d(s_45_0), .cin(t_338), .o(t_344), .co(t_345), .cout(t_346)); 
compressor_4_2 u2_125(.a(s_45_7), .b(s_45_6), .c(s_45_5), .d(s_45_4), .cin(t_341), .o(t_347), .co(t_348), .cout(t_349)); 
compressor_3_2 u1_126(.a(s_45_10), .b(s_45_9), .cin(s_45_8), .o(t_350), .cout(t_351)); 
compressor_4_2 u2_127(.a(s_46_3), .b(s_46_2), .c(s_46_1), .d(s_46_0), .cin(t_346), .o(t_352), .co(t_353), .cout(t_354)); 
compressor_4_2 u2_128(.a(s_46_7), .b(s_46_6), .c(s_46_5), .d(s_46_4), .cin(t_349), .o(t_355), .co(t_356), .cout(t_357)); 
half_adder u0_129(.a(s_46_9), .b(s_46_8), .o(t_358), .cout(t_359)); 
compressor_4_2 u2_130(.a(s_47_3), .b(s_47_2), .c(s_47_1), .d(s_47_0), .cin(t_354), .o(t_360), .co(t_361), .cout(t_362)); 
compressor_4_2 u2_131(.a(s_47_7), .b(s_47_6), .c(s_47_5), .d(s_47_4), .cin(t_357), .o(t_363), .co(t_364), .cout(t_365)); 
half_adder u0_132(.a(s_47_9), .b(s_47_8), .o(t_366), .cout(t_367)); 
compressor_4_2 u2_133(.a(s_48_3), .b(s_48_2), .c(s_48_1), .d(s_48_0), .cin(t_362), .o(t_368), .co(t_369), .cout(t_370)); 
compressor_4_2 u2_134(.a(s_48_7), .b(s_48_6), .c(s_48_5), .d(s_48_4), .cin(t_365), .o(t_371), .co(t_372), .cout(t_373)); 
compressor_4_2 u2_135(.a(s_49_3), .b(s_49_2), .c(s_49_1), .d(s_49_0), .cin(t_370), .o(t_374), .co(t_375), .cout(t_376)); 
compressor_4_2 u2_136(.a(s_49_7), .b(s_49_6), .c(s_49_5), .d(s_49_4), .cin(t_373), .o(t_377), .co(t_378), .cout(t_379)); 
compressor_4_2 u2_137(.a(s_50_3), .b(s_50_2), .c(s_50_1), .d(s_50_0), .cin(t_376), .o(t_380), .co(t_381), .cout(t_382)); 
compressor_4_2 u2_138(.a(s_50_7), .b(s_50_6), .c(s_50_5), .d(s_50_4), .cin(t_379), .o(t_383), .co(t_384), .cout(t_385)); 
compressor_4_2 u2_139(.a(s_51_3), .b(s_51_2), .c(s_51_1), .d(s_51_0), .cin(t_382), .o(t_386), .co(t_387), .cout(t_388)); 
compressor_4_2 u2_140(.a(s_51_7), .b(s_51_6), .c(s_51_5), .d(s_51_4), .cin(t_385), .o(t_389), .co(t_390), .cout(t_391)); 
compressor_4_2 u2_141(.a(s_52_3), .b(s_52_2), .c(s_52_1), .d(s_52_0), .cin(t_388), .o(t_392), .co(t_393), .cout(t_394)); 
compressor_3_2 u1_142(.a(s_52_5), .b(s_52_4), .cin(t_391), .o(t_395), .cout(t_396)); 
compressor_4_2 u2_143(.a(s_53_3), .b(s_53_2), .c(s_53_1), .d(s_53_0), .cin(t_394), .o(t_397), .co(t_398), .cout(t_399)); 
compressor_3_2 u1_144(.a(s_53_6), .b(s_53_5), .cin(s_53_4), .o(t_400), .cout(t_401)); 
compressor_4_2 u2_145(.a(s_54_3), .b(s_54_2), .c(s_54_1), .d(s_54_0), .cin(t_399), .o(t_402), .co(t_403), .cout(t_404)); 
half_adder u0_146(.a(s_54_5), .b(s_54_4), .o(t_405), .cout(t_406)); 
compressor_4_2 u2_147(.a(s_55_3), .b(s_55_2), .c(s_55_1), .d(s_55_0), .cin(t_404), .o(t_407), .co(t_408), .cout(t_409)); 
half_adder u0_148(.a(s_55_5), .b(s_55_4), .o(t_410), .cout(t_411)); 
compressor_4_2 u2_149(.a(s_56_3), .b(s_56_2), .c(s_56_1), .d(s_56_0), .cin(t_409), .o(t_412), .co(t_413), .cout(t_414)); 
compressor_4_2 u2_150(.a(s_57_3), .b(s_57_2), .c(s_57_1), .d(s_57_0), .cin(t_414), .o(t_415), .co(t_416), .cout(t_417)); 
compressor_4_2 u2_151(.a(s_58_3), .b(s_58_2), .c(s_58_1), .d(s_58_0), .cin(t_417), .o(t_418), .co(t_419), .cout(t_420)); 
compressor_4_2 u2_152(.a(s_59_3), .b(s_59_2), .c(s_59_1), .d(s_59_0), .cin(t_420), .o(t_421), .co(t_422), .cout(t_423)); 
compressor_3_2 u1_153(.a(s_60_1), .b(s_60_0), .cin(t_423), .o(t_424), .cout(t_425)); 
compressor_3_2 u1_154(.a(s_61_2), .b(s_61_1), .cin(s_61_0), .o(t_426), .cout(t_427)); 
half_adder u0_155(.a(s_62_1), .b(s_62_0), .o(t_428), .cout(t_429)); 
half_adder u0_156(.a(s_63_1), .b(s_63_0), .o(t_430), .cout()); 

/* u0_157 Output nets */
wire  t_431, t_432;  
/* u0_158 Output nets */
wire  t_433, t_434;  
/* u1_159 Output nets */
wire  t_435, t_436;  
/* u0_160 Output nets */
wire  t_437, t_438;  
/* u0_161 Output nets */
wire  t_439, t_440;  
/* u0_162 Output nets */
wire  t_441, t_442;  
/* u1_163 Output nets */
wire  t_443, t_444;  
/* u1_164 Output nets */
wire  t_445, t_446;  
/* u1_165 Output nets */
wire  t_447, t_448;  
/* u1_166 Output nets */
wire  t_449, t_450;  
/* u2_167 Output nets */
wire  t_451, t_452, t_453;  
/* u2_168 Output nets */
wire  t_454, t_455, t_456;  
/* u2_169 Output nets */
wire  t_457, t_458, t_459;  
/* u2_170 Output nets */
wire  t_460, t_461, t_462;  
/* u2_171 Output nets */
wire  t_463, t_464, t_465;  
/* u2_172 Output nets */
wire  t_466, t_467, t_468;  
/* u0_173 Output nets */
wire  t_469, t_470;  
/* u2_174 Output nets */
wire  t_471, t_472, t_473;  
/* u2_175 Output nets */
wire  t_474, t_475, t_476;  
/* u0_176 Output nets */
wire  t_477, t_478;  
/* u2_177 Output nets */
wire  t_479, t_480, t_481;  
/* u1_178 Output nets */
wire  t_482, t_483;  
/* u2_179 Output nets */
wire  t_484, t_485, t_486;  
/* u0_180 Output nets */
wire  t_487, t_488;  
/* u2_181 Output nets */
wire  t_489, t_490, t_491;  
/* u0_182 Output nets */
wire  t_492, t_493;  
/* u2_183 Output nets */
wire  t_494, t_495, t_496;  
/* u0_184 Output nets */
wire  t_497, t_498;  
/* u2_185 Output nets */
wire  t_499, t_500, t_501;  
/* u1_186 Output nets */
wire  t_502, t_503;  
/* u2_187 Output nets */
wire  t_504, t_505, t_506;  
/* u1_188 Output nets */
wire  t_507, t_508;  
/* u2_189 Output nets */
wire  t_509, t_510, t_511;  
/* u1_190 Output nets */
wire  t_512, t_513;  
/* u2_191 Output nets */
wire  t_514, t_515, t_516;  
/* u1_192 Output nets */
wire  t_517, t_518;  
/* u2_193 Output nets */
wire  t_519, t_520, t_521;  
/* u2_194 Output nets */
wire  t_522, t_523, t_524;  
/* u2_195 Output nets */
wire  t_525, t_526, t_527;  
/* u2_196 Output nets */
wire  t_528, t_529, t_530;  
/* u2_197 Output nets */
wire  t_531, t_532, t_533;  
/* u2_198 Output nets */
wire  t_534, t_535, t_536;  
/* u2_199 Output nets */
wire  t_537, t_538, t_539;  
/* u2_200 Output nets */
wire  t_540, t_541, t_542;  
/* u2_201 Output nets */
wire  t_543, t_544, t_545;  
/* u2_202 Output nets */
wire  t_546, t_547, t_548;  
/* u2_203 Output nets */
wire  t_549, t_550, t_551;  
/* u2_204 Output nets */
wire  t_552, t_553, t_554;  
/* u2_205 Output nets */
wire  t_555, t_556, t_557;  
/* u2_206 Output nets */
wire  t_558, t_559, t_560;  
/* u2_207 Output nets */
wire  t_561, t_562, t_563;  
/* u2_208 Output nets */
wire  t_564, t_565, t_566;  
/* u2_209 Output nets */
wire  t_567, t_568, t_569;  
/* u2_210 Output nets */
wire  t_570, t_571, t_572;  
/* u2_211 Output nets */
wire  t_573, t_574, t_575;  
/* u2_212 Output nets */
wire  t_576, t_577, t_578;  
/* u2_213 Output nets */
wire  t_579, t_580, t_581;  
/* u2_214 Output nets */
wire  t_582, t_583, t_584;  
/* u2_215 Output nets */
wire  t_585, t_586, t_587;  
/* u2_216 Output nets */
wire  t_588, t_589, t_590;  
/* u2_217 Output nets */
wire  t_591, t_592, t_593;  
/* u2_218 Output nets */
wire  t_594, t_595, t_596;  
/* u2_219 Output nets */
wire  t_597, t_598, t_599;  
/* u1_220 Output nets */
wire  t_600, t_601;  
/* u2_221 Output nets */
wire  t_602, t_603, t_604;  
/* u0_222 Output nets */
wire  t_605, t_606;  
/* u2_223 Output nets */
wire  t_607, t_608, t_609;  
/* u0_224 Output nets */
wire  t_610, t_611;  
/* u2_225 Output nets */
wire  t_612, t_613, t_614;  
/* u1_226 Output nets */
wire  t_615, t_616;  
/* u2_227 Output nets */
wire  t_617, t_618, t_619;  
/* u0_228 Output nets */
wire  t_620, t_621;  
/* u2_229 Output nets */
wire  t_622, t_623, t_624;  
/* u0_230 Output nets */
wire  t_625, t_626;  
/* u2_231 Output nets */
wire  t_627, t_628, t_629;  
/* u0_232 Output nets */
wire  t_630, t_631;  
/* u2_233 Output nets */
wire  t_632, t_633, t_634;  
/* u0_234 Output nets */
wire  t_635, t_636;  
/* u2_235 Output nets */
wire  t_637, t_638, t_639;  
/* u2_236 Output nets */
wire  t_640, t_641, t_642;  
/* u2_237 Output nets */
wire  t_643, t_644, t_645;  
/* u2_238 Output nets */
wire  t_646, t_647, t_648;  
/* u2_239 Output nets */
wire  t_649, t_650, t_651;  
/* u2_240 Output nets */
wire  t_652, t_653, t_654;  
/* u2_241 Output nets */
wire  t_655, t_656, t_657;  
/* u2_242 Output nets */
wire  t_658, t_659, t_660;  
/* u1_243 Output nets */
wire  t_661, t_662;  
/* u0_244 Output nets */
wire  t_663, t_664;  
/* u0_245 Output nets */
wire  t_665, t_666;  
/* u1_246 Output nets */
wire  t_667, t_668;  
/* u0_247 Output nets */
wire  t_669, t_670;  
/* u0_248 Output nets */
wire  t_671, t_672;  
/* u0_249 Output nets */
wire  t_673;  

/* compress stage 2 */
half_adder u0_157(.a(t_1), .b(s_1_0), .o(t_431), .cout(t_432)); 
half_adder u0_158(.a(t_4), .b(t_3), .o(t_433), .cout(t_434)); 
compressor_3_2 u1_159(.a(t_6), .b(t_5), .cin(s_4_3), .o(t_435), .cout(t_436)); 
half_adder u0_160(.a(t_8), .b(t_7), .o(t_437), .cout(t_438)); 
half_adder u0_161(.a(t_10), .b(t_9), .o(t_439), .cout(t_440)); 
half_adder u0_162(.a(t_13), .b(t_11), .o(t_441), .cout(t_442)); 
compressor_3_2 u1_163(.a(t_19), .b(t_16), .cin(t_14), .o(t_443), .cout(t_444)); 
compressor_3_2 u1_164(.a(t_20), .b(t_17), .cin(s_9_4), .o(t_445), .cout(t_446)); 
compressor_3_2 u1_165(.a(t_27), .b(t_24), .cin(t_22), .o(t_447), .cout(t_448)); 
compressor_3_2 u1_166(.a(t_29), .b(t_28), .cin(t_25), .o(t_449), .cout(t_450)); 
compressor_4_2 u2_167(.a(t_37), .b(t_34), .c(t_33), .d(t_30), .cin(s_12_7), .o(t_451), .co(t_452), .cout(t_453)); 
compressor_4_2 u2_168(.a(t_42), .b(t_39), .c(t_38), .d(t_35), .cin(t_453), .o(t_454), .co(t_455), .cout(t_456)); 
compressor_4_2 u2_169(.a(t_47), .b(t_44), .c(t_43), .d(t_40), .cin(t_456), .o(t_457), .co(t_458), .cout(t_459)); 
compressor_4_2 u2_170(.a(t_53), .b(t_50), .c(t_48), .d(t_45), .cin(t_459), .o(t_460), .co(t_461), .cout(t_462)); 
compressor_4_2 u2_171(.a(t_59), .b(t_56), .c(t_54), .d(t_51), .cin(t_462), .o(t_463), .co(t_464), .cout(t_465)); 
compressor_4_2 u2_172(.a(t_63), .b(t_60), .c(t_57), .d(s_17_8), .cin(t_465), .o(t_466), .co(t_467), .cout(t_468)); 
half_adder u0_173(.a(t_67), .b(t_64), .o(t_469), .cout(t_470)); 
compressor_4_2 u2_174(.a(t_73), .b(t_70), .c(t_68), .d(t_65), .cin(t_468), .o(t_471), .co(t_472), .cout(t_473)); 
compressor_4_2 u2_175(.a(t_78), .b(t_77), .c(t_74), .d(t_71), .cin(t_473), .o(t_474), .co(t_475), .cout(t_476)); 
half_adder u0_176(.a(t_84), .b(t_81), .o(t_477), .cout(t_478)); 
compressor_4_2 u2_177(.a(t_85), .b(t_82), .c(t_79), .d(s_20_11), .cin(t_476), .o(t_479), .co(t_480), .cout(t_481)); 
compressor_3_2 u1_178(.a(t_92), .b(t_89), .cin(t_86), .o(t_482), .cout(t_483)); 
compressor_4_2 u2_179(.a(t_94), .b(t_93), .c(t_90), .d(t_87), .cin(t_481), .o(t_484), .co(t_485), .cout(t_486)); 
half_adder u0_180(.a(t_100), .b(t_97), .o(t_487), .cout(t_488)); 
compressor_4_2 u2_181(.a(t_102), .b(t_101), .c(t_98), .d(t_95), .cin(t_486), .o(t_489), .co(t_490), .cout(t_491)); 
half_adder u0_182(.a(t_108), .b(t_105), .o(t_492), .cout(t_493)); 
compressor_4_2 u2_183(.a(t_111), .b(t_109), .c(t_106), .d(t_103), .cin(t_491), .o(t_494), .co(t_495), .cout(t_496)); 
half_adder u0_184(.a(t_117), .b(t_114), .o(t_497), .cout(t_498)); 
compressor_4_2 u2_185(.a(t_120), .b(t_118), .c(t_115), .d(t_112), .cin(t_496), .o(t_499), .co(t_500), .cout(t_501)); 
compressor_3_2 u1_186(.a(t_129), .b(t_126), .cin(t_123), .o(t_502), .cout(t_503)); 
compressor_4_2 u2_187(.a(t_127), .b(t_124), .c(t_121), .d(s_25_12), .cin(t_501), .o(t_504), .co(t_505), .cout(t_506)); 
compressor_3_2 u1_188(.a(t_134), .b(t_131), .cin(t_130), .o(t_507), .cout(t_508)); 
compressor_4_2 u2_189(.a(t_140), .b(t_138), .c(t_135), .d(t_132), .cin(t_506), .o(t_509), .co(t_510), .cout(t_511)); 
compressor_3_2 u1_190(.a(t_149), .b(t_146), .cin(t_143), .o(t_512), .cout(t_513)); 
compressor_4_2 u2_191(.a(t_150), .b(t_147), .c(t_144), .d(t_141), .cin(t_511), .o(t_514), .co(t_515), .cout(t_516)); 
compressor_3_2 u1_192(.a(t_157), .b(t_154), .cin(t_151), .o(t_517), .cout(t_518)); 
compressor_4_2 u2_193(.a(t_158), .b(t_155), .c(t_152), .d(s_28_15), .cin(t_516), .o(t_519), .co(t_520), .cout(t_521)); 
compressor_4_2 u2_194(.a(t_171), .b(t_168), .c(t_165), .d(t_162), .cin(t_161), .o(t_522), .co(t_523), .cout(t_524)); 
compressor_4_2 u2_195(.a(t_172), .b(t_169), .c(t_166), .d(t_163), .cin(t_521), .o(t_525), .co(t_526), .cout(t_527)); 
compressor_4_2 u2_196(.a(t_182), .b(t_179), .c(t_176), .d(t_173), .cin(t_524), .o(t_528), .co(t_529), .cout(t_530)); 
compressor_4_2 u2_197(.a(t_183), .b(t_180), .c(t_177), .d(t_174), .cin(t_527), .o(t_531), .co(t_532), .cout(t_533)); 
compressor_4_2 u2_198(.a(t_193), .b(t_190), .c(t_187), .d(t_184), .cin(t_530), .o(t_534), .co(t_535), .cout(t_536)); 
compressor_4_2 u2_199(.a(t_194), .b(t_191), .c(t_188), .d(t_185), .cin(t_533), .o(t_537), .co(t_538), .cout(t_539)); 
compressor_4_2 u2_200(.a(t_205), .b(t_202), .c(t_199), .d(t_196), .cin(t_536), .o(t_540), .co(t_541), .cout(t_542)); 
compressor_4_2 u2_201(.a(t_203), .b(t_200), .c(t_197), .d(s_32_16), .cin(t_539), .o(t_543), .co(t_544), .cout(t_545)); 
compressor_4_2 u2_202(.a(t_214), .b(t_211), .c(t_208), .d(t_206), .cin(t_542), .o(t_546), .co(t_547), .cout(t_548)); 
compressor_4_2 u2_203(.a(t_215), .b(t_212), .c(t_209), .d(s_33_16), .cin(t_545), .o(t_549), .co(t_550), .cout(t_551)); 
compressor_4_2 u2_204(.a(t_226), .b(t_223), .c(t_220), .d(t_218), .cin(t_548), .o(t_552), .co(t_553), .cout(t_554)); 
compressor_4_2 u2_205(.a(t_230), .b(t_227), .c(t_224), .d(t_221), .cin(t_551), .o(t_555), .co(t_556), .cout(t_557)); 
compressor_4_2 u2_206(.a(t_241), .b(t_238), .c(t_235), .d(t_232), .cin(t_554), .o(t_558), .co(t_559), .cout(t_560)); 
compressor_4_2 u2_207(.a(t_242), .b(t_239), .c(t_236), .d(t_233), .cin(t_557), .o(t_561), .co(t_562), .cout(t_563)); 
compressor_4_2 u2_208(.a(t_253), .b(t_250), .c(t_247), .d(t_244), .cin(t_560), .o(t_564), .co(t_565), .cout(t_566)); 
compressor_4_2 u2_209(.a(t_251), .b(t_248), .c(t_245), .d(s_36_14), .cin(t_563), .o(t_567), .co(t_568), .cout(t_569)); 
compressor_4_2 u2_210(.a(t_262), .b(t_259), .c(t_256), .d(t_254), .cin(t_566), .o(t_570), .co(t_571), .cout(t_572)); 
compressor_4_2 u2_211(.a(t_266), .b(t_263), .c(t_260), .d(t_257), .cin(t_569), .o(t_573), .co(t_574), .cout(t_575)); 
compressor_4_2 u2_212(.a(t_276), .b(t_273), .c(t_270), .d(t_267), .cin(t_572), .o(t_576), .co(t_577), .cout(t_578)); 
compressor_4_2 u2_213(.a(t_277), .b(t_274), .c(t_271), .d(t_268), .cin(t_575), .o(t_579), .co(t_580), .cout(t_581)); 
compressor_4_2 u2_214(.a(t_287), .b(t_284), .c(t_281), .d(t_278), .cin(t_578), .o(t_582), .co(t_583), .cout(t_584)); 
compressor_4_2 u2_215(.a(t_288), .b(t_285), .c(t_282), .d(t_279), .cin(t_581), .o(t_585), .co(t_586), .cout(t_587)); 
compressor_4_2 u2_216(.a(t_298), .b(t_295), .c(t_292), .d(t_289), .cin(t_584), .o(t_588), .co(t_589), .cout(t_590)); 
compressor_4_2 u2_217(.a(t_296), .b(t_293), .c(t_290), .d(s_40_12), .cin(t_587), .o(t_591), .co(t_592), .cout(t_593)); 
compressor_4_2 u2_218(.a(t_306), .b(t_303), .c(t_300), .d(t_299), .cin(t_590), .o(t_594), .co(t_595), .cout(t_596)); 
compressor_4_2 u2_219(.a(t_307), .b(t_304), .c(t_301), .d(s_41_12), .cin(t_593), .o(t_597), .co(t_598), .cout(t_599)); 
compressor_3_2 u1_220(.a(t_312), .b(t_309), .cin(t_596), .o(t_600), .cout(t_601)); 
compressor_4_2 u2_221(.a(t_318), .b(t_316), .c(t_313), .d(t_310), .cin(t_599), .o(t_602), .co(t_603), .cout(t_604)); 
half_adder u0_222(.a(t_324), .b(t_321), .o(t_605), .cout(t_606)); 
compressor_4_2 u2_223(.a(t_327), .b(t_325), .c(t_322), .d(t_319), .cin(t_604), .o(t_607), .co(t_608), .cout(t_609)); 
half_adder u0_224(.a(t_333), .b(t_330), .o(t_610), .cout(t_611)); 
compressor_4_2 u2_225(.a(t_334), .b(t_331), .c(t_328), .d(s_44_10), .cin(t_609), .o(t_612), .co(t_613), .cout(t_614)); 
compressor_3_2 u1_226(.a(t_342), .b(t_339), .cin(t_336), .o(t_615), .cout(t_616)); 
compressor_4_2 u2_227(.a(t_344), .b(t_343), .c(t_340), .d(t_337), .cin(t_614), .o(t_617), .co(t_618), .cout(t_619)); 
half_adder u0_228(.a(t_350), .b(t_347), .o(t_620), .cout(t_621)); 
compressor_4_2 u2_229(.a(t_352), .b(t_351), .c(t_348), .d(t_345), .cin(t_619), .o(t_622), .co(t_623), .cout(t_624)); 
half_adder u0_230(.a(t_358), .b(t_355), .o(t_625), .cout(t_626)); 
compressor_4_2 u2_231(.a(t_360), .b(t_359), .c(t_356), .d(t_353), .cin(t_624), .o(t_627), .co(t_628), .cout(t_629)); 
half_adder u0_232(.a(t_366), .b(t_363), .o(t_630), .cout(t_631)); 
compressor_4_2 u2_233(.a(t_367), .b(t_364), .c(t_361), .d(s_48_8), .cin(t_629), .o(t_632), .co(t_633), .cout(t_634)); 
half_adder u0_234(.a(t_371), .b(t_368), .o(t_635), .cout(t_636)); 
compressor_4_2 u2_235(.a(t_374), .b(t_372), .c(t_369), .d(s_49_8), .cin(t_634), .o(t_637), .co(t_638), .cout(t_639)); 
compressor_4_2 u2_236(.a(t_383), .b(t_380), .c(t_378), .d(t_375), .cin(t_639), .o(t_640), .co(t_641), .cout(t_642)); 
compressor_4_2 u2_237(.a(t_389), .b(t_386), .c(t_384), .d(t_381), .cin(t_642), .o(t_643), .co(t_644), .cout(t_645)); 
compressor_4_2 u2_238(.a(t_392), .b(t_390), .c(t_387), .d(s_52_6), .cin(t_645), .o(t_646), .co(t_647), .cout(t_648)); 
compressor_4_2 u2_239(.a(t_400), .b(t_397), .c(t_396), .d(t_393), .cin(t_648), .o(t_649), .co(t_650), .cout(t_651)); 
compressor_4_2 u2_240(.a(t_405), .b(t_402), .c(t_401), .d(t_398), .cin(t_651), .o(t_652), .co(t_653), .cout(t_654)); 
compressor_4_2 u2_241(.a(t_410), .b(t_407), .c(t_406), .d(t_403), .cin(t_654), .o(t_655), .co(t_656), .cout(t_657)); 
compressor_4_2 u2_242(.a(t_412), .b(t_411), .c(t_408), .d(s_56_4), .cin(t_657), .o(t_658), .co(t_659), .cout(t_660)); 
compressor_3_2 u1_243(.a(t_413), .b(s_57_4), .cin(t_660), .o(t_661), .cout(t_662)); 
half_adder u0_244(.a(t_418), .b(t_416), .o(t_663), .cout(t_664)); 
half_adder u0_245(.a(t_421), .b(t_419), .o(t_665), .cout(t_666)); 
compressor_3_2 u1_246(.a(t_424), .b(t_422), .cin(s_60_2), .o(t_667), .cout(t_668)); 
half_adder u0_247(.a(t_426), .b(t_425), .o(t_669), .cout(t_670)); 
half_adder u0_248(.a(t_428), .b(t_427), .o(t_671), .cout(t_672)); 
half_adder u0_249(.a(t_430), .b(t_429), .o(t_673), .cout()); 

/* u0_250 Output nets */
wire  t_674, t_675;  
/* u0_251 Output nets */
wire  t_676, t_677;  
/* u0_252 Output nets */
wire  t_678, t_679;  
/* u0_253 Output nets */
wire  t_680, t_681;  
/* u0_254 Output nets */
wire  t_682, t_683;  
/* u0_255 Output nets */
wire  t_684, t_685;  
/* u1_256 Output nets */
wire  t_686, t_687;  
/* u0_257 Output nets */
wire  t_688, t_689;  
/* u1_258 Output nets */
wire  t_690, t_691;  
/* u0_259 Output nets */
wire  t_692, t_693;  
/* u0_260 Output nets */
wire  t_694, t_695;  
/* u0_261 Output nets */
wire  t_696, t_697;  
/* u0_262 Output nets */
wire  t_698, t_699;  
/* u1_263 Output nets */
wire  t_700, t_701;  
/* u1_264 Output nets */
wire  t_702, t_703;  
/* u1_265 Output nets */
wire  t_704, t_705;  
/* u1_266 Output nets */
wire  t_706, t_707;  
/* u1_267 Output nets */
wire  t_708, t_709;  
/* u1_268 Output nets */
wire  t_710, t_711;  
/* u1_269 Output nets */
wire  t_712, t_713;  
/* u1_270 Output nets */
wire  t_714, t_715;  
/* u1_271 Output nets */
wire  t_716, t_717;  
/* u2_272 Output nets */
wire  t_718, t_719, t_720;  
/* u2_273 Output nets */
wire  t_721, t_722, t_723;  
/* u2_274 Output nets */
wire  t_724, t_725, t_726;  
/* u2_275 Output nets */
wire  t_727, t_728, t_729;  
/* u2_276 Output nets */
wire  t_730, t_731, t_732;  
/* u2_277 Output nets */
wire  t_733, t_734, t_735;  
/* u2_278 Output nets */
wire  t_736, t_737, t_738;  
/* u2_279 Output nets */
wire  t_739, t_740, t_741;  
/* u2_280 Output nets */
wire  t_742, t_743, t_744;  
/* u2_281 Output nets */
wire  t_745, t_746, t_747;  
/* u2_282 Output nets */
wire  t_748, t_749, t_750;  
/* u2_283 Output nets */
wire  t_751, t_752, t_753;  
/* u2_284 Output nets */
wire  t_754, t_755, t_756;  
/* u2_285 Output nets */
wire  t_757, t_758, t_759;  
/* u2_286 Output nets */
wire  t_760, t_761, t_762;  
/* u2_287 Output nets */
wire  t_763, t_764, t_765;  
/* u2_288 Output nets */
wire  t_766, t_767, t_768;  
/* u2_289 Output nets */
wire  t_769, t_770, t_771;  
/* u2_290 Output nets */
wire  t_772, t_773, t_774;  
/* u2_291 Output nets */
wire  t_775, t_776, t_777;  
/* u2_292 Output nets */
wire  t_778, t_779, t_780;  
/* u2_293 Output nets */
wire  t_781, t_782, t_783;  
/* u2_294 Output nets */
wire  t_784, t_785, t_786;  
/* u2_295 Output nets */
wire  t_787, t_788, t_789;  
/* u2_296 Output nets */
wire  t_790, t_791, t_792;  
/* u1_297 Output nets */
wire  t_793, t_794;  
/* u0_298 Output nets */
wire  t_795, t_796;  
/* u1_299 Output nets */
wire  t_797, t_798;  
/* u0_300 Output nets */
wire  t_799, t_800;  
/* u0_301 Output nets */
wire  t_801, t_802;  
/* u0_302 Output nets */
wire  t_803, t_804;  
/* u0_303 Output nets */
wire  t_805, t_806;  
/* u1_304 Output nets */
wire  t_807, t_808;  
/* u0_305 Output nets */
wire  t_809, t_810;  
/* u0_306 Output nets */
wire  t_811, t_812;  
/* u0_307 Output nets */
wire  t_813, t_814;  
/* u0_308 Output nets */
wire  t_815, t_816;  
/* u0_309 Output nets */
wire  t_817, t_818;  
/* u0_310 Output nets */
wire  t_819;  

/* compress stage 3 */
half_adder u0_250(.a(t_432), .b(t_2), .o(t_674), .cout(t_675)); 
half_adder u0_251(.a(t_435), .b(t_434), .o(t_676), .cout(t_677)); 
half_adder u0_252(.a(t_437), .b(t_436), .o(t_678), .cout(t_679)); 
half_adder u0_253(.a(t_439), .b(t_438), .o(t_680), .cout(t_681)); 
half_adder u0_254(.a(t_441), .b(t_440), .o(t_682), .cout(t_683)); 
half_adder u0_255(.a(t_443), .b(t_442), .o(t_684), .cout(t_685)); 
compressor_3_2 u1_256(.a(t_445), .b(t_444), .cin(t_21), .o(t_686), .cout(t_687)); 
half_adder u0_257(.a(t_447), .b(t_446), .o(t_688), .cout(t_689)); 
compressor_3_2 u1_258(.a(t_449), .b(t_448), .cin(t_32), .o(t_690), .cout(t_691)); 
half_adder u0_259(.a(t_451), .b(t_450), .o(t_692), .cout(t_693)); 
half_adder u0_260(.a(t_454), .b(t_452), .o(t_694), .cout(t_695)); 
half_adder u0_261(.a(t_457), .b(t_455), .o(t_696), .cout(t_697)); 
half_adder u0_262(.a(t_460), .b(t_458), .o(t_698), .cout(t_699)); 
compressor_3_2 u1_263(.a(t_463), .b(t_461), .cin(t_62), .o(t_700), .cout(t_701)); 
compressor_3_2 u1_264(.a(t_469), .b(t_466), .cin(t_464), .o(t_702), .cout(t_703)); 
compressor_3_2 u1_265(.a(t_470), .b(t_467), .cin(t_76), .o(t_704), .cout(t_705)); 
compressor_3_2 u1_266(.a(t_477), .b(t_474), .cin(t_472), .o(t_706), .cout(t_707)); 
compressor_3_2 u1_267(.a(t_479), .b(t_478), .cin(t_475), .o(t_708), .cout(t_709)); 
compressor_3_2 u1_268(.a(t_484), .b(t_483), .cin(t_480), .o(t_710), .cout(t_711)); 
compressor_3_2 u1_269(.a(t_489), .b(t_488), .cin(t_485), .o(t_712), .cout(t_713)); 
compressor_3_2 u1_270(.a(t_494), .b(t_493), .cin(t_490), .o(t_714), .cout(t_715)); 
compressor_3_2 u1_271(.a(t_499), .b(t_498), .cin(t_495), .o(t_716), .cout(t_717)); 
compressor_4_2 u2_272(.a(t_507), .b(t_504), .c(t_503), .d(t_500), .cin(t_137), .o(t_718), .co(t_719), .cout(t_720)); 
compressor_4_2 u2_273(.a(t_512), .b(t_509), .c(t_508), .d(t_505), .cin(t_720), .o(t_721), .co(t_722), .cout(t_723)); 
compressor_4_2 u2_274(.a(t_514), .b(t_513), .c(t_510), .d(t_160), .cin(t_723), .o(t_724), .co(t_725), .cout(t_726)); 
compressor_4_2 u2_275(.a(t_522), .b(t_519), .c(t_518), .d(t_515), .cin(t_726), .o(t_727), .co(t_728), .cout(t_729)); 
compressor_4_2 u2_276(.a(t_528), .b(t_525), .c(t_523), .d(t_520), .cin(t_729), .o(t_730), .co(t_731), .cout(t_732)); 
compressor_4_2 u2_277(.a(t_534), .b(t_531), .c(t_529), .d(t_526), .cin(t_732), .o(t_733), .co(t_734), .cout(t_735)); 
compressor_4_2 u2_278(.a(t_540), .b(t_537), .c(t_535), .d(t_532), .cin(t_735), .o(t_736), .co(t_737), .cout(t_738)); 
compressor_4_2 u2_279(.a(t_543), .b(t_541), .c(t_538), .d(t_217), .cin(t_738), .o(t_739), .co(t_740), .cout(t_741)); 
compressor_4_2 u2_280(.a(t_549), .b(t_547), .c(t_544), .d(t_229), .cin(t_741), .o(t_742), .co(t_743), .cout(t_744)); 
compressor_4_2 u2_281(.a(t_558), .b(t_555), .c(t_553), .d(t_550), .cin(t_744), .o(t_745), .co(t_746), .cout(t_747)); 
compressor_4_2 u2_282(.a(t_564), .b(t_561), .c(t_559), .d(t_556), .cin(t_747), .o(t_748), .co(t_749), .cout(t_750)); 
compressor_4_2 u2_283(.a(t_567), .b(t_565), .c(t_562), .d(t_265), .cin(t_750), .o(t_751), .co(t_752), .cout(t_753)); 
compressor_4_2 u2_284(.a(t_576), .b(t_573), .c(t_571), .d(t_568), .cin(t_753), .o(t_754), .co(t_755), .cout(t_756)); 
compressor_4_2 u2_285(.a(t_582), .b(t_579), .c(t_577), .d(t_574), .cin(t_756), .o(t_757), .co(t_758), .cout(t_759)); 
compressor_4_2 u2_286(.a(t_588), .b(t_585), .c(t_583), .d(t_580), .cin(t_759), .o(t_760), .co(t_761), .cout(t_762)); 
compressor_4_2 u2_287(.a(t_594), .b(t_591), .c(t_589), .d(t_586), .cin(t_762), .o(t_763), .co(t_764), .cout(t_765)); 
compressor_4_2 u2_288(.a(t_597), .b(t_595), .c(t_592), .d(t_315), .cin(t_765), .o(t_766), .co(t_767), .cout(t_768)); 
compressor_4_2 u2_289(.a(t_605), .b(t_602), .c(t_601), .d(t_598), .cin(t_768), .o(t_769), .co(t_770), .cout(t_771)); 
compressor_4_2 u2_290(.a(t_610), .b(t_607), .c(t_606), .d(t_603), .cin(t_771), .o(t_772), .co(t_773), .cout(t_774)); 
compressor_4_2 u2_291(.a(t_615), .b(t_612), .c(t_611), .d(t_608), .cin(t_774), .o(t_775), .co(t_776), .cout(t_777)); 
compressor_4_2 u2_292(.a(t_620), .b(t_617), .c(t_616), .d(t_613), .cin(t_777), .o(t_778), .co(t_779), .cout(t_780)); 
compressor_4_2 u2_293(.a(t_625), .b(t_622), .c(t_621), .d(t_618), .cin(t_780), .o(t_781), .co(t_782), .cout(t_783)); 
compressor_4_2 u2_294(.a(t_630), .b(t_627), .c(t_626), .d(t_623), .cin(t_783), .o(t_784), .co(t_785), .cout(t_786)); 
compressor_4_2 u2_295(.a(t_635), .b(t_632), .c(t_631), .d(t_628), .cin(t_786), .o(t_787), .co(t_788), .cout(t_789)); 
compressor_4_2 u2_296(.a(t_637), .b(t_636), .c(t_633), .d(t_377), .cin(t_789), .o(t_790), .co(t_791), .cout(t_792)); 
compressor_3_2 u1_297(.a(t_640), .b(t_638), .cin(t_792), .o(t_793), .cout(t_794)); 
half_adder u0_298(.a(t_643), .b(t_641), .o(t_795), .cout(t_796)); 
compressor_3_2 u1_299(.a(t_646), .b(t_644), .cin(t_395), .o(t_797), .cout(t_798)); 
half_adder u0_300(.a(t_649), .b(t_647), .o(t_799), .cout(t_800)); 
half_adder u0_301(.a(t_652), .b(t_650), .o(t_801), .cout(t_802)); 
half_adder u0_302(.a(t_655), .b(t_653), .o(t_803), .cout(t_804)); 
half_adder u0_303(.a(t_658), .b(t_656), .o(t_805), .cout(t_806)); 
compressor_3_2 u1_304(.a(t_661), .b(t_659), .cin(t_415), .o(t_807), .cout(t_808)); 
half_adder u0_305(.a(t_663), .b(t_662), .o(t_809), .cout(t_810)); 
half_adder u0_306(.a(t_665), .b(t_664), .o(t_811), .cout(t_812)); 
half_adder u0_307(.a(t_667), .b(t_666), .o(t_813), .cout(t_814)); 
half_adder u0_308(.a(t_669), .b(t_668), .o(t_815), .cout(t_816)); 
half_adder u0_309(.a(t_671), .b(t_670), .o(t_817), .cout(t_818)); 
half_adder u0_310(.a(t_673), .b(t_672), .o(t_819), .cout()); 

/* u0_311 Output nets */
wire  t_820, t_821;  
/* u0_312 Output nets */
wire  t_822, t_823;  
/* u0_313 Output nets */
wire  t_824, t_825;  
/* u0_314 Output nets */
wire  t_826, t_827;  
/* u0_315 Output nets */
wire  t_828, t_829;  
/* u0_316 Output nets */
wire  t_830, t_831;  
/* u0_317 Output nets */
wire  t_832, t_833;  
/* u0_318 Output nets */
wire  t_834, t_835;  
/* u0_319 Output nets */
wire  t_836, t_837;  
/* u0_320 Output nets */
wire  t_838, t_839;  
/* u0_321 Output nets */
wire  t_840, t_841;  
/* u0_322 Output nets */
wire  t_842, t_843;  
/* u0_323 Output nets */
wire  t_844, t_845;  
/* u0_324 Output nets */
wire  t_846, t_847;  
/* u1_325 Output nets */
wire  t_848, t_849;  
/* u0_326 Output nets */
wire  t_850, t_851;  
/* u1_327 Output nets */
wire  t_852, t_853;  
/* u1_328 Output nets */
wire  t_854, t_855;  
/* u1_329 Output nets */
wire  t_856, t_857;  
/* u1_330 Output nets */
wire  t_858, t_859;  
/* u1_331 Output nets */
wire  t_860, t_861;  
/* u0_332 Output nets */
wire  t_862, t_863;  
/* u0_333 Output nets */
wire  t_864, t_865;  
/* u1_334 Output nets */
wire  t_866, t_867;  
/* u0_335 Output nets */
wire  t_868, t_869;  
/* u0_336 Output nets */
wire  t_870, t_871;  
/* u0_337 Output nets */
wire  t_872, t_873;  
/* u0_338 Output nets */
wire  t_874, t_875;  
/* u1_339 Output nets */
wire  t_876, t_877;  
/* u1_340 Output nets */
wire  t_878, t_879;  
/* u0_341 Output nets */
wire  t_880, t_881;  
/* u0_342 Output nets */
wire  t_882, t_883;  
/* u1_343 Output nets */
wire  t_884, t_885;  
/* u0_344 Output nets */
wire  t_886, t_887;  
/* u0_345 Output nets */
wire  t_888, t_889;  
/* u0_346 Output nets */
wire  t_890, t_891;  
/* u0_347 Output nets */
wire  t_892, t_893;  
/* u1_348 Output nets */
wire  t_894, t_895;  
/* u0_349 Output nets */
wire  t_896, t_897;  
/* u0_350 Output nets */
wire  t_898, t_899;  
/* u0_351 Output nets */
wire  t_900, t_901;  
/* u0_352 Output nets */
wire  t_902, t_903;  
/* u0_353 Output nets */
wire  t_904, t_905;  
/* u0_354 Output nets */
wire  t_906, t_907;  
/* u0_355 Output nets */
wire  t_908, t_909;  
/* u0_356 Output nets */
wire  t_910, t_911;  
/* u0_357 Output nets */
wire  t_912, t_913;  
/* u0_358 Output nets */
wire  t_914, t_915;  
/* u0_359 Output nets */
wire  t_916, t_917;  
/* u0_360 Output nets */
wire  t_918, t_919;  
/* u0_361 Output nets */
wire  t_920, t_921;  
/* u0_362 Output nets */
wire  t_922, t_923;  
/* u0_363 Output nets */
wire  t_924, t_925;  
/* u0_364 Output nets */
wire  t_926, t_927;  
/* u0_365 Output nets */
wire  t_928, t_929;  
/* u0_366 Output nets */
wire  t_930, t_931;  
/* u0_367 Output nets */
wire  t_932, t_933;  
/* u0_368 Output nets */
wire  t_934, t_935;  
/* u0_369 Output nets */
wire  t_936, t_937;  
/* u0_370 Output nets */
wire  t_938;  

/* compress stage 4 */
half_adder u0_311(.a(t_675), .b(t_433), .o(t_820), .cout(t_821)); 
half_adder u0_312(.a(t_678), .b(t_677), .o(t_822), .cout(t_823)); 
half_adder u0_313(.a(t_680), .b(t_679), .o(t_824), .cout(t_825)); 
half_adder u0_314(.a(t_682), .b(t_681), .o(t_826), .cout(t_827)); 
half_adder u0_315(.a(t_684), .b(t_683), .o(t_828), .cout(t_829)); 
half_adder u0_316(.a(t_686), .b(t_685), .o(t_830), .cout(t_831)); 
half_adder u0_317(.a(t_688), .b(t_687), .o(t_832), .cout(t_833)); 
half_adder u0_318(.a(t_690), .b(t_689), .o(t_834), .cout(t_835)); 
half_adder u0_319(.a(t_692), .b(t_691), .o(t_836), .cout(t_837)); 
half_adder u0_320(.a(t_694), .b(t_693), .o(t_838), .cout(t_839)); 
half_adder u0_321(.a(t_696), .b(t_695), .o(t_840), .cout(t_841)); 
half_adder u0_322(.a(t_698), .b(t_697), .o(t_842), .cout(t_843)); 
half_adder u0_323(.a(t_700), .b(t_699), .o(t_844), .cout(t_845)); 
half_adder u0_324(.a(t_702), .b(t_701), .o(t_846), .cout(t_847)); 
compressor_3_2 u1_325(.a(t_704), .b(t_703), .cin(t_471), .o(t_848), .cout(t_849)); 
half_adder u0_326(.a(t_706), .b(t_705), .o(t_850), .cout(t_851)); 
compressor_3_2 u1_327(.a(t_708), .b(t_707), .cin(t_482), .o(t_852), .cout(t_853)); 
compressor_3_2 u1_328(.a(t_710), .b(t_709), .cin(t_487), .o(t_854), .cout(t_855)); 
compressor_3_2 u1_329(.a(t_712), .b(t_711), .cin(t_492), .o(t_856), .cout(t_857)); 
compressor_3_2 u1_330(.a(t_714), .b(t_713), .cin(t_497), .o(t_858), .cout(t_859)); 
compressor_3_2 u1_331(.a(t_716), .b(t_715), .cin(t_502), .o(t_860), .cout(t_861)); 
half_adder u0_332(.a(t_718), .b(t_717), .o(t_862), .cout(t_863)); 
half_adder u0_333(.a(t_721), .b(t_719), .o(t_864), .cout(t_865)); 
compressor_3_2 u1_334(.a(t_724), .b(t_722), .cin(t_517), .o(t_866), .cout(t_867)); 
half_adder u0_335(.a(t_727), .b(t_725), .o(t_868), .cout(t_869)); 
half_adder u0_336(.a(t_730), .b(t_728), .o(t_870), .cout(t_871)); 
half_adder u0_337(.a(t_733), .b(t_731), .o(t_872), .cout(t_873)); 
half_adder u0_338(.a(t_736), .b(t_734), .o(t_874), .cout(t_875)); 
compressor_3_2 u1_339(.a(t_739), .b(t_737), .cin(t_546), .o(t_876), .cout(t_877)); 
compressor_3_2 u1_340(.a(t_742), .b(t_740), .cin(t_552), .o(t_878), .cout(t_879)); 
half_adder u0_341(.a(t_745), .b(t_743), .o(t_880), .cout(t_881)); 
half_adder u0_342(.a(t_748), .b(t_746), .o(t_882), .cout(t_883)); 
compressor_3_2 u1_343(.a(t_751), .b(t_749), .cin(t_570), .o(t_884), .cout(t_885)); 
half_adder u0_344(.a(t_754), .b(t_752), .o(t_886), .cout(t_887)); 
half_adder u0_345(.a(t_757), .b(t_755), .o(t_888), .cout(t_889)); 
half_adder u0_346(.a(t_760), .b(t_758), .o(t_890), .cout(t_891)); 
half_adder u0_347(.a(t_763), .b(t_761), .o(t_892), .cout(t_893)); 
compressor_3_2 u1_348(.a(t_766), .b(t_764), .cin(t_600), .o(t_894), .cout(t_895)); 
half_adder u0_349(.a(t_769), .b(t_767), .o(t_896), .cout(t_897)); 
half_adder u0_350(.a(t_772), .b(t_770), .o(t_898), .cout(t_899)); 
half_adder u0_351(.a(t_775), .b(t_773), .o(t_900), .cout(t_901)); 
half_adder u0_352(.a(t_778), .b(t_776), .o(t_902), .cout(t_903)); 
half_adder u0_353(.a(t_781), .b(t_779), .o(t_904), .cout(t_905)); 
half_adder u0_354(.a(t_784), .b(t_782), .o(t_906), .cout(t_907)); 
half_adder u0_355(.a(t_787), .b(t_785), .o(t_908), .cout(t_909)); 
half_adder u0_356(.a(t_790), .b(t_788), .o(t_910), .cout(t_911)); 
half_adder u0_357(.a(t_793), .b(t_791), .o(t_912), .cout(t_913)); 
half_adder u0_358(.a(t_795), .b(t_794), .o(t_914), .cout(t_915)); 
half_adder u0_359(.a(t_797), .b(t_796), .o(t_916), .cout(t_917)); 
half_adder u0_360(.a(t_799), .b(t_798), .o(t_918), .cout(t_919)); 
half_adder u0_361(.a(t_801), .b(t_800), .o(t_920), .cout(t_921)); 
half_adder u0_362(.a(t_803), .b(t_802), .o(t_922), .cout(t_923)); 
half_adder u0_363(.a(t_805), .b(t_804), .o(t_924), .cout(t_925)); 
half_adder u0_364(.a(t_807), .b(t_806), .o(t_926), .cout(t_927)); 
half_adder u0_365(.a(t_809), .b(t_808), .o(t_928), .cout(t_929)); 
half_adder u0_366(.a(t_811), .b(t_810), .o(t_930), .cout(t_931)); 
half_adder u0_367(.a(t_813), .b(t_812), .o(t_932), .cout(t_933)); 
half_adder u0_368(.a(t_815), .b(t_814), .o(t_934), .cout(t_935)); 
half_adder u0_369(.a(t_817), .b(t_816), .o(t_936), .cout(t_937)); 
half_adder u0_370(.a(t_819), .b(t_818), .o(t_938), .cout()); 

/* Output nets Compression result */
assign compress_a = {
   t_937,   t_935,   t_933,   t_931,
   t_929,   t_927,   t_925,   t_923,
   t_921,   t_919,   t_917,   t_915,
   t_913,   t_911,   t_909,   t_907,
   t_905,   t_903,   t_901,   t_899,
   t_897,   t_895,   t_893,   t_891,
   t_889,   t_887,   t_885,   t_883,
   t_881,   t_879,   t_877,   t_875,
   t_873,   t_871,   t_869,   t_867,
   t_865,   t_863,   t_861,   t_859,
   t_857,   t_855,   t_853,   t_851,
   t_849,   t_847,   t_845,   t_843,
   t_841,   t_839,   t_837,   t_835,
   t_833,   t_831,   t_829,   t_827,
   t_825,   t_823,   t_822,   t_676,
   t_820,   t_674,   t_431,     t_0
};
assign compress_b = {
   t_938,   t_936,   t_934,   t_932,
   t_930,   t_928,   t_926,   t_924,
   t_922,   t_920,   t_918,   t_916,
   t_914,   t_912,   t_910,   t_908,
   t_906,   t_904,   t_902,   t_900,
   t_898,   t_896,   t_894,   t_892,
   t_890,   t_888,   t_886,   t_884,
   t_882,   t_880,   t_878,   t_876,
   t_874,   t_872,   t_870,   t_868,
   t_866,   t_864,   t_862,   t_860,
   t_858,   t_856,   t_854,   t_852,
   t_850,   t_848,   t_846,   t_844,
   t_842,   t_840,   t_838,   t_836,
   t_834,   t_832,   t_830,   t_828,
   t_826,   t_824,    1'b0,   t_821,
    1'b0,    1'b0,    1'b0,    1'b0
};

endmodule

/********************************************************************************/

module _64_wallace_tree(
//inputs
	partial_products,
	carry,
//outputs
	compress_a,
	compress_b
);

localparam width = 64;

input wire [(width+2)*(width/2+1)-1:0] partial_products;
input wire [width/2-1:0] carry;
output wire [2*width-1:0] compress_a;
output wire [2*width-1:0] compress_b;

/* Input nets */
wire    s_0_0,    s_0_1,    s_1_0,    s_2_0,    s_2_1,    s_2_2;
wire    s_3_0,    s_3_1,    s_4_0,    s_4_1,    s_4_2,    s_4_3;
wire    s_5_0,    s_5_1,    s_5_2,    s_6_0,    s_6_1,    s_6_2;
wire    s_6_3,    s_6_4,    s_7_0,    s_7_1,    s_7_2,    s_7_3;
wire    s_8_0,    s_8_1,    s_8_2,    s_8_3,    s_8_4,    s_8_5;
wire    s_9_0,    s_9_1,    s_9_2,    s_9_3,    s_9_4,   s_10_0;
wire   s_10_1,   s_10_2,   s_10_3,   s_10_4,   s_10_5,   s_10_6;
wire   s_11_0,   s_11_1,   s_11_2,   s_11_3,   s_11_4,   s_11_5;
wire   s_12_0,   s_12_1,   s_12_2,   s_12_3,   s_12_4,   s_12_5;
wire   s_12_6,   s_12_7,   s_13_0,   s_13_1,   s_13_2,   s_13_3;
wire   s_13_4,   s_13_5,   s_13_6,   s_14_0,   s_14_1,   s_14_2;
wire   s_14_3,   s_14_4,   s_14_5,   s_14_6,   s_14_7,   s_14_8;
wire   s_15_0,   s_15_1,   s_15_2,   s_15_3,   s_15_4,   s_15_5;
wire   s_15_6,   s_15_7,   s_16_0,   s_16_1,   s_16_2,   s_16_3;
wire   s_16_4,   s_16_5,   s_16_6,   s_16_7,   s_16_8,   s_16_9;
wire   s_17_0,   s_17_1,   s_17_2,   s_17_3,   s_17_4,   s_17_5;
wire   s_17_6,   s_17_7,   s_17_8,   s_18_0,   s_18_1,   s_18_2;
wire   s_18_3,   s_18_4,   s_18_5,   s_18_6,   s_18_7,   s_18_8;
wire   s_18_9,  s_18_10,   s_19_0,   s_19_1,   s_19_2,   s_19_3;
wire   s_19_4,   s_19_5,   s_19_6,   s_19_7,   s_19_8,   s_19_9;
wire   s_20_0,   s_20_1,   s_20_2,   s_20_3,   s_20_4,   s_20_5;
wire   s_20_6,   s_20_7,   s_20_8,   s_20_9,  s_20_10,  s_20_11;
wire   s_21_0,   s_21_1,   s_21_2,   s_21_3,   s_21_4,   s_21_5;
wire   s_21_6,   s_21_7,   s_21_8,   s_21_9,  s_21_10,   s_22_0;
wire   s_22_1,   s_22_2,   s_22_3,   s_22_4,   s_22_5,   s_22_6;
wire   s_22_7,   s_22_8,   s_22_9,  s_22_10,  s_22_11,  s_22_12;
wire   s_23_0,   s_23_1,   s_23_2,   s_23_3,   s_23_4,   s_23_5;
wire   s_23_6,   s_23_7,   s_23_8,   s_23_9,  s_23_10,  s_23_11;
wire   s_24_0,   s_24_1,   s_24_2,   s_24_3,   s_24_4,   s_24_5;
wire   s_24_6,   s_24_7,   s_24_8,   s_24_9,  s_24_10,  s_24_11;
wire  s_24_12,  s_24_13,   s_25_0,   s_25_1,   s_25_2,   s_25_3;
wire   s_25_4,   s_25_5,   s_25_6,   s_25_7,   s_25_8,   s_25_9;
wire  s_25_10,  s_25_11,  s_25_12,   s_26_0,   s_26_1,   s_26_2;
wire   s_26_3,   s_26_4,   s_26_5,   s_26_6,   s_26_7,   s_26_8;
wire   s_26_9,  s_26_10,  s_26_11,  s_26_12,  s_26_13,  s_26_14;
wire   s_27_0,   s_27_1,   s_27_2,   s_27_3,   s_27_4,   s_27_5;
wire   s_27_6,   s_27_7,   s_27_8,   s_27_9,  s_27_10,  s_27_11;
wire  s_27_12,  s_27_13,   s_28_0,   s_28_1,   s_28_2,   s_28_3;
wire   s_28_4,   s_28_5,   s_28_6,   s_28_7,   s_28_8,   s_28_9;
wire  s_28_10,  s_28_11,  s_28_12,  s_28_13,  s_28_14,  s_28_15;
wire   s_29_0,   s_29_1,   s_29_2,   s_29_3,   s_29_4,   s_29_5;
wire   s_29_6,   s_29_7,   s_29_8,   s_29_9,  s_29_10,  s_29_11;
wire  s_29_12,  s_29_13,  s_29_14,   s_30_0,   s_30_1,   s_30_2;
wire   s_30_3,   s_30_4,   s_30_5,   s_30_6,   s_30_7,   s_30_8;
wire   s_30_9,  s_30_10,  s_30_11,  s_30_12,  s_30_13,  s_30_14;
wire  s_30_15,  s_30_16,   s_31_0,   s_31_1,   s_31_2,   s_31_3;
wire   s_31_4,   s_31_5,   s_31_6,   s_31_7,   s_31_8,   s_31_9;
wire  s_31_10,  s_31_11,  s_31_12,  s_31_13,  s_31_14,  s_31_15;
wire   s_32_0,   s_32_1,   s_32_2,   s_32_3,   s_32_4,   s_32_5;
wire   s_32_6,   s_32_7,   s_32_8,   s_32_9,  s_32_10,  s_32_11;
wire  s_32_12,  s_32_13,  s_32_14,  s_32_15,  s_32_16,  s_32_17;
wire   s_33_0,   s_33_1,   s_33_2,   s_33_3,   s_33_4,   s_33_5;
wire   s_33_6,   s_33_7,   s_33_8,   s_33_9,  s_33_10,  s_33_11;
wire  s_33_12,  s_33_13,  s_33_14,  s_33_15,  s_33_16,   s_34_0;
wire   s_34_1,   s_34_2,   s_34_3,   s_34_4,   s_34_5,   s_34_6;
wire   s_34_7,   s_34_8,   s_34_9,  s_34_10,  s_34_11,  s_34_12;
wire  s_34_13,  s_34_14,  s_34_15,  s_34_16,  s_34_17,  s_34_18;
wire   s_35_0,   s_35_1,   s_35_2,   s_35_3,   s_35_4,   s_35_5;
wire   s_35_6,   s_35_7,   s_35_8,   s_35_9,  s_35_10,  s_35_11;
wire  s_35_12,  s_35_13,  s_35_14,  s_35_15,  s_35_16,  s_35_17;
wire   s_36_0,   s_36_1,   s_36_2,   s_36_3,   s_36_4,   s_36_5;
wire   s_36_6,   s_36_7,   s_36_8,   s_36_9,  s_36_10,  s_36_11;
wire  s_36_12,  s_36_13,  s_36_14,  s_36_15,  s_36_16,  s_36_17;
wire  s_36_18,  s_36_19,   s_37_0,   s_37_1,   s_37_2,   s_37_3;
wire   s_37_4,   s_37_5,   s_37_6,   s_37_7,   s_37_8,   s_37_9;
wire  s_37_10,  s_37_11,  s_37_12,  s_37_13,  s_37_14,  s_37_15;
wire  s_37_16,  s_37_17,  s_37_18,   s_38_0,   s_38_1,   s_38_2;
wire   s_38_3,   s_38_4,   s_38_5,   s_38_6,   s_38_7,   s_38_8;
wire   s_38_9,  s_38_10,  s_38_11,  s_38_12,  s_38_13,  s_38_14;
wire  s_38_15,  s_38_16,  s_38_17,  s_38_18,  s_38_19,  s_38_20;
wire   s_39_0,   s_39_1,   s_39_2,   s_39_3,   s_39_4,   s_39_5;
wire   s_39_6,   s_39_7,   s_39_8,   s_39_9,  s_39_10,  s_39_11;
wire  s_39_12,  s_39_13,  s_39_14,  s_39_15,  s_39_16,  s_39_17;
wire  s_39_18,  s_39_19,   s_40_0,   s_40_1,   s_40_2,   s_40_3;
wire   s_40_4,   s_40_5,   s_40_6,   s_40_7,   s_40_8,   s_40_9;
wire  s_40_10,  s_40_11,  s_40_12,  s_40_13,  s_40_14,  s_40_15;
wire  s_40_16,  s_40_17,  s_40_18,  s_40_19,  s_40_20,  s_40_21;
wire   s_41_0,   s_41_1,   s_41_2,   s_41_3,   s_41_4,   s_41_5;
wire   s_41_6,   s_41_7,   s_41_8,   s_41_9,  s_41_10,  s_41_11;
wire  s_41_12,  s_41_13,  s_41_14,  s_41_15,  s_41_16,  s_41_17;
wire  s_41_18,  s_41_19,  s_41_20,   s_42_0,   s_42_1,   s_42_2;
wire   s_42_3,   s_42_4,   s_42_5,   s_42_6,   s_42_7,   s_42_8;
wire   s_42_9,  s_42_10,  s_42_11,  s_42_12,  s_42_13,  s_42_14;
wire  s_42_15,  s_42_16,  s_42_17,  s_42_18,  s_42_19,  s_42_20;
wire  s_42_21,  s_42_22,   s_43_0,   s_43_1,   s_43_2,   s_43_3;
wire   s_43_4,   s_43_5,   s_43_6,   s_43_7,   s_43_8,   s_43_9;
wire  s_43_10,  s_43_11,  s_43_12,  s_43_13,  s_43_14,  s_43_15;
wire  s_43_16,  s_43_17,  s_43_18,  s_43_19,  s_43_20,  s_43_21;
wire   s_44_0,   s_44_1,   s_44_2,   s_44_3,   s_44_4,   s_44_5;
wire   s_44_6,   s_44_7,   s_44_8,   s_44_9,  s_44_10,  s_44_11;
wire  s_44_12,  s_44_13,  s_44_14,  s_44_15,  s_44_16,  s_44_17;
wire  s_44_18,  s_44_19,  s_44_20,  s_44_21,  s_44_22,  s_44_23;
wire   s_45_0,   s_45_1,   s_45_2,   s_45_3,   s_45_4,   s_45_5;
wire   s_45_6,   s_45_7,   s_45_8,   s_45_9,  s_45_10,  s_45_11;
wire  s_45_12,  s_45_13,  s_45_14,  s_45_15,  s_45_16,  s_45_17;
wire  s_45_18,  s_45_19,  s_45_20,  s_45_21,  s_45_22,   s_46_0;
wire   s_46_1,   s_46_2,   s_46_3,   s_46_4,   s_46_5,   s_46_6;
wire   s_46_7,   s_46_8,   s_46_9,  s_46_10,  s_46_11,  s_46_12;
wire  s_46_13,  s_46_14,  s_46_15,  s_46_16,  s_46_17,  s_46_18;
wire  s_46_19,  s_46_20,  s_46_21,  s_46_22,  s_46_23,  s_46_24;
wire   s_47_0,   s_47_1,   s_47_2,   s_47_3,   s_47_4,   s_47_5;
wire   s_47_6,   s_47_7,   s_47_8,   s_47_9,  s_47_10,  s_47_11;
wire  s_47_12,  s_47_13,  s_47_14,  s_47_15,  s_47_16,  s_47_17;
wire  s_47_18,  s_47_19,  s_47_20,  s_47_21,  s_47_22,  s_47_23;
wire   s_48_0,   s_48_1,   s_48_2,   s_48_3,   s_48_4,   s_48_5;
wire   s_48_6,   s_48_7,   s_48_8,   s_48_9,  s_48_10,  s_48_11;
wire  s_48_12,  s_48_13,  s_48_14,  s_48_15,  s_48_16,  s_48_17;
wire  s_48_18,  s_48_19,  s_48_20,  s_48_21,  s_48_22,  s_48_23;
wire  s_48_24,  s_48_25,   s_49_0,   s_49_1,   s_49_2,   s_49_3;
wire   s_49_4,   s_49_5,   s_49_6,   s_49_7,   s_49_8,   s_49_9;
wire  s_49_10,  s_49_11,  s_49_12,  s_49_13,  s_49_14,  s_49_15;
wire  s_49_16,  s_49_17,  s_49_18,  s_49_19,  s_49_20,  s_49_21;
wire  s_49_22,  s_49_23,  s_49_24,   s_50_0,   s_50_1,   s_50_2;
wire   s_50_3,   s_50_4,   s_50_5,   s_50_6,   s_50_7,   s_50_8;
wire   s_50_9,  s_50_10,  s_50_11,  s_50_12,  s_50_13,  s_50_14;
wire  s_50_15,  s_50_16,  s_50_17,  s_50_18,  s_50_19,  s_50_20;
wire  s_50_21,  s_50_22,  s_50_23,  s_50_24,  s_50_25,  s_50_26;
wire   s_51_0,   s_51_1,   s_51_2,   s_51_3,   s_51_4,   s_51_5;
wire   s_51_6,   s_51_7,   s_51_8,   s_51_9,  s_51_10,  s_51_11;
wire  s_51_12,  s_51_13,  s_51_14,  s_51_15,  s_51_16,  s_51_17;
wire  s_51_18,  s_51_19,  s_51_20,  s_51_21,  s_51_22,  s_51_23;
wire  s_51_24,  s_51_25,   s_52_0,   s_52_1,   s_52_2,   s_52_3;
wire   s_52_4,   s_52_5,   s_52_6,   s_52_7,   s_52_8,   s_52_9;
wire  s_52_10,  s_52_11,  s_52_12,  s_52_13,  s_52_14,  s_52_15;
wire  s_52_16,  s_52_17,  s_52_18,  s_52_19,  s_52_20,  s_52_21;
wire  s_52_22,  s_52_23,  s_52_24,  s_52_25,  s_52_26,  s_52_27;
wire   s_53_0,   s_53_1,   s_53_2,   s_53_3,   s_53_4,   s_53_5;
wire   s_53_6,   s_53_7,   s_53_8,   s_53_9,  s_53_10,  s_53_11;
wire  s_53_12,  s_53_13,  s_53_14,  s_53_15,  s_53_16,  s_53_17;
wire  s_53_18,  s_53_19,  s_53_20,  s_53_21,  s_53_22,  s_53_23;
wire  s_53_24,  s_53_25,  s_53_26,   s_54_0,   s_54_1,   s_54_2;
wire   s_54_3,   s_54_4,   s_54_5,   s_54_6,   s_54_7,   s_54_8;
wire   s_54_9,  s_54_10,  s_54_11,  s_54_12,  s_54_13,  s_54_14;
wire  s_54_15,  s_54_16,  s_54_17,  s_54_18,  s_54_19,  s_54_20;
wire  s_54_21,  s_54_22,  s_54_23,  s_54_24,  s_54_25,  s_54_26;
wire  s_54_27,  s_54_28,   s_55_0,   s_55_1,   s_55_2,   s_55_3;
wire   s_55_4,   s_55_5,   s_55_6,   s_55_7,   s_55_8,   s_55_9;
wire  s_55_10,  s_55_11,  s_55_12,  s_55_13,  s_55_14,  s_55_15;
wire  s_55_16,  s_55_17,  s_55_18,  s_55_19,  s_55_20,  s_55_21;
wire  s_55_22,  s_55_23,  s_55_24,  s_55_25,  s_55_26,  s_55_27;
wire   s_56_0,   s_56_1,   s_56_2,   s_56_3,   s_56_4,   s_56_5;
wire   s_56_6,   s_56_7,   s_56_8,   s_56_9,  s_56_10,  s_56_11;
wire  s_56_12,  s_56_13,  s_56_14,  s_56_15,  s_56_16,  s_56_17;
wire  s_56_18,  s_56_19,  s_56_20,  s_56_21,  s_56_22,  s_56_23;
wire  s_56_24,  s_56_25,  s_56_26,  s_56_27,  s_56_28,  s_56_29;
wire   s_57_0,   s_57_1,   s_57_2,   s_57_3,   s_57_4,   s_57_5;
wire   s_57_6,   s_57_7,   s_57_8,   s_57_9,  s_57_10,  s_57_11;
wire  s_57_12,  s_57_13,  s_57_14,  s_57_15,  s_57_16,  s_57_17;
wire  s_57_18,  s_57_19,  s_57_20,  s_57_21,  s_57_22,  s_57_23;
wire  s_57_24,  s_57_25,  s_57_26,  s_57_27,  s_57_28,   s_58_0;
wire   s_58_1,   s_58_2,   s_58_3,   s_58_4,   s_58_5,   s_58_6;
wire   s_58_7,   s_58_8,   s_58_9,  s_58_10,  s_58_11,  s_58_12;
wire  s_58_13,  s_58_14,  s_58_15,  s_58_16,  s_58_17,  s_58_18;
wire  s_58_19,  s_58_20,  s_58_21,  s_58_22,  s_58_23,  s_58_24;
wire  s_58_25,  s_58_26,  s_58_27,  s_58_28,  s_58_29,  s_58_30;
wire   s_59_0,   s_59_1,   s_59_2,   s_59_3,   s_59_4,   s_59_5;
wire   s_59_6,   s_59_7,   s_59_8,   s_59_9,  s_59_10,  s_59_11;
wire  s_59_12,  s_59_13,  s_59_14,  s_59_15,  s_59_16,  s_59_17;
wire  s_59_18,  s_59_19,  s_59_20,  s_59_21,  s_59_22,  s_59_23;
wire  s_59_24,  s_59_25,  s_59_26,  s_59_27,  s_59_28,  s_59_29;
wire   s_60_0,   s_60_1,   s_60_2,   s_60_3,   s_60_4,   s_60_5;
wire   s_60_6,   s_60_7,   s_60_8,   s_60_9,  s_60_10,  s_60_11;
wire  s_60_12,  s_60_13,  s_60_14,  s_60_15,  s_60_16,  s_60_17;
wire  s_60_18,  s_60_19,  s_60_20,  s_60_21,  s_60_22,  s_60_23;
wire  s_60_24,  s_60_25,  s_60_26,  s_60_27,  s_60_28,  s_60_29;
wire  s_60_30,  s_60_31,   s_61_0,   s_61_1,   s_61_2,   s_61_3;
wire   s_61_4,   s_61_5,   s_61_6,   s_61_7,   s_61_8,   s_61_9;
wire  s_61_10,  s_61_11,  s_61_12,  s_61_13,  s_61_14,  s_61_15;
wire  s_61_16,  s_61_17,  s_61_18,  s_61_19,  s_61_20,  s_61_21;
wire  s_61_22,  s_61_23,  s_61_24,  s_61_25,  s_61_26,  s_61_27;
wire  s_61_28,  s_61_29,  s_61_30,   s_62_0,   s_62_1,   s_62_2;
wire   s_62_3,   s_62_4,   s_62_5,   s_62_6,   s_62_7,   s_62_8;
wire   s_62_9,  s_62_10,  s_62_11,  s_62_12,  s_62_13,  s_62_14;
wire  s_62_15,  s_62_16,  s_62_17,  s_62_18,  s_62_19,  s_62_20;
wire  s_62_21,  s_62_22,  s_62_23,  s_62_24,  s_62_25,  s_62_26;
wire  s_62_27,  s_62_28,  s_62_29,  s_62_30,  s_62_31,  s_62_32;
wire   s_63_0,   s_63_1,   s_63_2,   s_63_3,   s_63_4,   s_63_5;
wire   s_63_6,   s_63_7,   s_63_8,   s_63_9,  s_63_10,  s_63_11;
wire  s_63_12,  s_63_13,  s_63_14,  s_63_15,  s_63_16,  s_63_17;
wire  s_63_18,  s_63_19,  s_63_20,  s_63_21,  s_63_22,  s_63_23;
wire  s_63_24,  s_63_25,  s_63_26,  s_63_27,  s_63_28,  s_63_29;
wire  s_63_30,  s_63_31,   s_64_0,   s_64_1,   s_64_2,   s_64_3;
wire   s_64_4,   s_64_5,   s_64_6,   s_64_7,   s_64_8,   s_64_9;
wire  s_64_10,  s_64_11,  s_64_12,  s_64_13,  s_64_14,  s_64_15;
wire  s_64_16,  s_64_17,  s_64_18,  s_64_19,  s_64_20,  s_64_21;
wire  s_64_22,  s_64_23,  s_64_24,  s_64_25,  s_64_26,  s_64_27;
wire  s_64_28,  s_64_29,  s_64_30,  s_64_31,  s_64_32,   s_65_0;
wire   s_65_1,   s_65_2,   s_65_3,   s_65_4,   s_65_5,   s_65_6;
wire   s_65_7,   s_65_8,   s_65_9,  s_65_10,  s_65_11,  s_65_12;
wire  s_65_13,  s_65_14,  s_65_15,  s_65_16,  s_65_17,  s_65_18;
wire  s_65_19,  s_65_20,  s_65_21,  s_65_22,  s_65_23,  s_65_24;
wire  s_65_25,  s_65_26,  s_65_27,  s_65_28,  s_65_29,  s_65_30;
wire  s_65_31,  s_65_32,   s_66_0,   s_66_1,   s_66_2,   s_66_3;
wire   s_66_4,   s_66_5,   s_66_6,   s_66_7,   s_66_8,   s_66_9;
wire  s_66_10,  s_66_11,  s_66_12,  s_66_13,  s_66_14,  s_66_15;
wire  s_66_16,  s_66_17,  s_66_18,  s_66_19,  s_66_20,  s_66_21;
wire  s_66_22,  s_66_23,  s_66_24,  s_66_25,  s_66_26,  s_66_27;
wire  s_66_28,  s_66_29,  s_66_30,  s_66_31,   s_67_0,   s_67_1;
wire   s_67_2,   s_67_3,   s_67_4,   s_67_5,   s_67_6,   s_67_7;
wire   s_67_8,   s_67_9,  s_67_10,  s_67_11,  s_67_12,  s_67_13;
wire  s_67_14,  s_67_15,  s_67_16,  s_67_17,  s_67_18,  s_67_19;
wire  s_67_20,  s_67_21,  s_67_22,  s_67_23,  s_67_24,  s_67_25;
wire  s_67_26,  s_67_27,  s_67_28,  s_67_29,  s_67_30,  s_67_31;
wire   s_68_0,   s_68_1,   s_68_2,   s_68_3,   s_68_4,   s_68_5;
wire   s_68_6,   s_68_7,   s_68_8,   s_68_9,  s_68_10,  s_68_11;
wire  s_68_12,  s_68_13,  s_68_14,  s_68_15,  s_68_16,  s_68_17;
wire  s_68_18,  s_68_19,  s_68_20,  s_68_21,  s_68_22,  s_68_23;
wire  s_68_24,  s_68_25,  s_68_26,  s_68_27,  s_68_28,  s_68_29;
wire  s_68_30,   s_69_0,   s_69_1,   s_69_2,   s_69_3,   s_69_4;
wire   s_69_5,   s_69_6,   s_69_7,   s_69_8,   s_69_9,  s_69_10;
wire  s_69_11,  s_69_12,  s_69_13,  s_69_14,  s_69_15,  s_69_16;
wire  s_69_17,  s_69_18,  s_69_19,  s_69_20,  s_69_21,  s_69_22;
wire  s_69_23,  s_69_24,  s_69_25,  s_69_26,  s_69_27,  s_69_28;
wire  s_69_29,  s_69_30,   s_70_0,   s_70_1,   s_70_2,   s_70_3;
wire   s_70_4,   s_70_5,   s_70_6,   s_70_7,   s_70_8,   s_70_9;
wire  s_70_10,  s_70_11,  s_70_12,  s_70_13,  s_70_14,  s_70_15;
wire  s_70_16,  s_70_17,  s_70_18,  s_70_19,  s_70_20,  s_70_21;
wire  s_70_22,  s_70_23,  s_70_24,  s_70_25,  s_70_26,  s_70_27;
wire  s_70_28,  s_70_29,   s_71_0,   s_71_1,   s_71_2,   s_71_3;
wire   s_71_4,   s_71_5,   s_71_6,   s_71_7,   s_71_8,   s_71_9;
wire  s_71_10,  s_71_11,  s_71_12,  s_71_13,  s_71_14,  s_71_15;
wire  s_71_16,  s_71_17,  s_71_18,  s_71_19,  s_71_20,  s_71_21;
wire  s_71_22,  s_71_23,  s_71_24,  s_71_25,  s_71_26,  s_71_27;
wire  s_71_28,  s_71_29,   s_72_0,   s_72_1,   s_72_2,   s_72_3;
wire   s_72_4,   s_72_5,   s_72_6,   s_72_7,   s_72_8,   s_72_9;
wire  s_72_10,  s_72_11,  s_72_12,  s_72_13,  s_72_14,  s_72_15;
wire  s_72_16,  s_72_17,  s_72_18,  s_72_19,  s_72_20,  s_72_21;
wire  s_72_22,  s_72_23,  s_72_24,  s_72_25,  s_72_26,  s_72_27;
wire  s_72_28,   s_73_0,   s_73_1,   s_73_2,   s_73_3,   s_73_4;
wire   s_73_5,   s_73_6,   s_73_7,   s_73_8,   s_73_9,  s_73_10;
wire  s_73_11,  s_73_12,  s_73_13,  s_73_14,  s_73_15,  s_73_16;
wire  s_73_17,  s_73_18,  s_73_19,  s_73_20,  s_73_21,  s_73_22;
wire  s_73_23,  s_73_24,  s_73_25,  s_73_26,  s_73_27,  s_73_28;
wire   s_74_0,   s_74_1,   s_74_2,   s_74_3,   s_74_4,   s_74_5;
wire   s_74_6,   s_74_7,   s_74_8,   s_74_9,  s_74_10,  s_74_11;
wire  s_74_12,  s_74_13,  s_74_14,  s_74_15,  s_74_16,  s_74_17;
wire  s_74_18,  s_74_19,  s_74_20,  s_74_21,  s_74_22,  s_74_23;
wire  s_74_24,  s_74_25,  s_74_26,  s_74_27,   s_75_0,   s_75_1;
wire   s_75_2,   s_75_3,   s_75_4,   s_75_5,   s_75_6,   s_75_7;
wire   s_75_8,   s_75_9,  s_75_10,  s_75_11,  s_75_12,  s_75_13;
wire  s_75_14,  s_75_15,  s_75_16,  s_75_17,  s_75_18,  s_75_19;
wire  s_75_20,  s_75_21,  s_75_22,  s_75_23,  s_75_24,  s_75_25;
wire  s_75_26,  s_75_27,   s_76_0,   s_76_1,   s_76_2,   s_76_3;
wire   s_76_4,   s_76_5,   s_76_6,   s_76_7,   s_76_8,   s_76_9;
wire  s_76_10,  s_76_11,  s_76_12,  s_76_13,  s_76_14,  s_76_15;
wire  s_76_16,  s_76_17,  s_76_18,  s_76_19,  s_76_20,  s_76_21;
wire  s_76_22,  s_76_23,  s_76_24,  s_76_25,  s_76_26,   s_77_0;
wire   s_77_1,   s_77_2,   s_77_3,   s_77_4,   s_77_5,   s_77_6;
wire   s_77_7,   s_77_8,   s_77_9,  s_77_10,  s_77_11,  s_77_12;
wire  s_77_13,  s_77_14,  s_77_15,  s_77_16,  s_77_17,  s_77_18;
wire  s_77_19,  s_77_20,  s_77_21,  s_77_22,  s_77_23,  s_77_24;
wire  s_77_25,  s_77_26,   s_78_0,   s_78_1,   s_78_2,   s_78_3;
wire   s_78_4,   s_78_5,   s_78_6,   s_78_7,   s_78_8,   s_78_9;
wire  s_78_10,  s_78_11,  s_78_12,  s_78_13,  s_78_14,  s_78_15;
wire  s_78_16,  s_78_17,  s_78_18,  s_78_19,  s_78_20,  s_78_21;
wire  s_78_22,  s_78_23,  s_78_24,  s_78_25,   s_79_0,   s_79_1;
wire   s_79_2,   s_79_3,   s_79_4,   s_79_5,   s_79_6,   s_79_7;
wire   s_79_8,   s_79_9,  s_79_10,  s_79_11,  s_79_12,  s_79_13;
wire  s_79_14,  s_79_15,  s_79_16,  s_79_17,  s_79_18,  s_79_19;
wire  s_79_20,  s_79_21,  s_79_22,  s_79_23,  s_79_24,  s_79_25;
wire   s_80_0,   s_80_1,   s_80_2,   s_80_3,   s_80_4,   s_80_5;
wire   s_80_6,   s_80_7,   s_80_8,   s_80_9,  s_80_10,  s_80_11;
wire  s_80_12,  s_80_13,  s_80_14,  s_80_15,  s_80_16,  s_80_17;
wire  s_80_18,  s_80_19,  s_80_20,  s_80_21,  s_80_22,  s_80_23;
wire  s_80_24,   s_81_0,   s_81_1,   s_81_2,   s_81_3,   s_81_4;
wire   s_81_5,   s_81_6,   s_81_7,   s_81_8,   s_81_9,  s_81_10;
wire  s_81_11,  s_81_12,  s_81_13,  s_81_14,  s_81_15,  s_81_16;
wire  s_81_17,  s_81_18,  s_81_19,  s_81_20,  s_81_21,  s_81_22;
wire  s_81_23,  s_81_24,   s_82_0,   s_82_1,   s_82_2,   s_82_3;
wire   s_82_4,   s_82_5,   s_82_6,   s_82_7,   s_82_8,   s_82_9;
wire  s_82_10,  s_82_11,  s_82_12,  s_82_13,  s_82_14,  s_82_15;
wire  s_82_16,  s_82_17,  s_82_18,  s_82_19,  s_82_20,  s_82_21;
wire  s_82_22,  s_82_23,   s_83_0,   s_83_1,   s_83_2,   s_83_3;
wire   s_83_4,   s_83_5,   s_83_6,   s_83_7,   s_83_8,   s_83_9;
wire  s_83_10,  s_83_11,  s_83_12,  s_83_13,  s_83_14,  s_83_15;
wire  s_83_16,  s_83_17,  s_83_18,  s_83_19,  s_83_20,  s_83_21;
wire  s_83_22,  s_83_23,   s_84_0,   s_84_1,   s_84_2,   s_84_3;
wire   s_84_4,   s_84_5,   s_84_6,   s_84_7,   s_84_8,   s_84_9;
wire  s_84_10,  s_84_11,  s_84_12,  s_84_13,  s_84_14,  s_84_15;
wire  s_84_16,  s_84_17,  s_84_18,  s_84_19,  s_84_20,  s_84_21;
wire  s_84_22,   s_85_0,   s_85_1,   s_85_2,   s_85_3,   s_85_4;
wire   s_85_5,   s_85_6,   s_85_7,   s_85_8,   s_85_9,  s_85_10;
wire  s_85_11,  s_85_12,  s_85_13,  s_85_14,  s_85_15,  s_85_16;
wire  s_85_17,  s_85_18,  s_85_19,  s_85_20,  s_85_21,  s_85_22;
wire   s_86_0,   s_86_1,   s_86_2,   s_86_3,   s_86_4,   s_86_5;
wire   s_86_6,   s_86_7,   s_86_8,   s_86_9,  s_86_10,  s_86_11;
wire  s_86_12,  s_86_13,  s_86_14,  s_86_15,  s_86_16,  s_86_17;
wire  s_86_18,  s_86_19,  s_86_20,  s_86_21,   s_87_0,   s_87_1;
wire   s_87_2,   s_87_3,   s_87_4,   s_87_5,   s_87_6,   s_87_7;
wire   s_87_8,   s_87_9,  s_87_10,  s_87_11,  s_87_12,  s_87_13;
wire  s_87_14,  s_87_15,  s_87_16,  s_87_17,  s_87_18,  s_87_19;
wire  s_87_20,  s_87_21,   s_88_0,   s_88_1,   s_88_2,   s_88_3;
wire   s_88_4,   s_88_5,   s_88_6,   s_88_7,   s_88_8,   s_88_9;
wire  s_88_10,  s_88_11,  s_88_12,  s_88_13,  s_88_14,  s_88_15;
wire  s_88_16,  s_88_17,  s_88_18,  s_88_19,  s_88_20,   s_89_0;
wire   s_89_1,   s_89_2,   s_89_3,   s_89_4,   s_89_5,   s_89_6;
wire   s_89_7,   s_89_8,   s_89_9,  s_89_10,  s_89_11,  s_89_12;
wire  s_89_13,  s_89_14,  s_89_15,  s_89_16,  s_89_17,  s_89_18;
wire  s_89_19,  s_89_20,   s_90_0,   s_90_1,   s_90_2,   s_90_3;
wire   s_90_4,   s_90_5,   s_90_6,   s_90_7,   s_90_8,   s_90_9;
wire  s_90_10,  s_90_11,  s_90_12,  s_90_13,  s_90_14,  s_90_15;
wire  s_90_16,  s_90_17,  s_90_18,  s_90_19,   s_91_0,   s_91_1;
wire   s_91_2,   s_91_3,   s_91_4,   s_91_5,   s_91_6,   s_91_7;
wire   s_91_8,   s_91_9,  s_91_10,  s_91_11,  s_91_12,  s_91_13;
wire  s_91_14,  s_91_15,  s_91_16,  s_91_17,  s_91_18,  s_91_19;
wire   s_92_0,   s_92_1,   s_92_2,   s_92_3,   s_92_4,   s_92_5;
wire   s_92_6,   s_92_7,   s_92_8,   s_92_9,  s_92_10,  s_92_11;
wire  s_92_12,  s_92_13,  s_92_14,  s_92_15,  s_92_16,  s_92_17;
wire  s_92_18,   s_93_0,   s_93_1,   s_93_2,   s_93_3,   s_93_4;
wire   s_93_5,   s_93_6,   s_93_7,   s_93_8,   s_93_9,  s_93_10;
wire  s_93_11,  s_93_12,  s_93_13,  s_93_14,  s_93_15,  s_93_16;
wire  s_93_17,  s_93_18,   s_94_0,   s_94_1,   s_94_2,   s_94_3;
wire   s_94_4,   s_94_5,   s_94_6,   s_94_7,   s_94_8,   s_94_9;
wire  s_94_10,  s_94_11,  s_94_12,  s_94_13,  s_94_14,  s_94_15;
wire  s_94_16,  s_94_17,   s_95_0,   s_95_1,   s_95_2,   s_95_3;
wire   s_95_4,   s_95_5,   s_95_6,   s_95_7,   s_95_8,   s_95_9;
wire  s_95_10,  s_95_11,  s_95_12,  s_95_13,  s_95_14,  s_95_15;
wire  s_95_16,  s_95_17,   s_96_0,   s_96_1,   s_96_2,   s_96_3;
wire   s_96_4,   s_96_5,   s_96_6,   s_96_7,   s_96_8,   s_96_9;
wire  s_96_10,  s_96_11,  s_96_12,  s_96_13,  s_96_14,  s_96_15;
wire  s_96_16,   s_97_0,   s_97_1,   s_97_2,   s_97_3,   s_97_4;
wire   s_97_5,   s_97_6,   s_97_7,   s_97_8,   s_97_9,  s_97_10;
wire  s_97_11,  s_97_12,  s_97_13,  s_97_14,  s_97_15,  s_97_16;
wire   s_98_0,   s_98_1,   s_98_2,   s_98_3,   s_98_4,   s_98_5;
wire   s_98_6,   s_98_7,   s_98_8,   s_98_9,  s_98_10,  s_98_11;
wire  s_98_12,  s_98_13,  s_98_14,  s_98_15,   s_99_0,   s_99_1;
wire   s_99_2,   s_99_3,   s_99_4,   s_99_5,   s_99_6,   s_99_7;
wire   s_99_8,   s_99_9,  s_99_10,  s_99_11,  s_99_12,  s_99_13;
wire  s_99_14,  s_99_15,  s_100_0,  s_100_1,  s_100_2,  s_100_3;
wire  s_100_4,  s_100_5,  s_100_6,  s_100_7,  s_100_8,  s_100_9;
wire s_100_10, s_100_11, s_100_12, s_100_13, s_100_14,  s_101_0;
wire  s_101_1,  s_101_2,  s_101_3,  s_101_4,  s_101_5,  s_101_6;
wire  s_101_7,  s_101_8,  s_101_9, s_101_10, s_101_11, s_101_12;
wire s_101_13, s_101_14,  s_102_0,  s_102_1,  s_102_2,  s_102_3;
wire  s_102_4,  s_102_5,  s_102_6,  s_102_7,  s_102_8,  s_102_9;
wire s_102_10, s_102_11, s_102_12, s_102_13,  s_103_0,  s_103_1;
wire  s_103_2,  s_103_3,  s_103_4,  s_103_5,  s_103_6,  s_103_7;
wire  s_103_8,  s_103_9, s_103_10, s_103_11, s_103_12, s_103_13;
wire  s_104_0,  s_104_1,  s_104_2,  s_104_3,  s_104_4,  s_104_5;
wire  s_104_6,  s_104_7,  s_104_8,  s_104_9, s_104_10, s_104_11;
wire s_104_12,  s_105_0,  s_105_1,  s_105_2,  s_105_3,  s_105_4;
wire  s_105_5,  s_105_6,  s_105_7,  s_105_8,  s_105_9, s_105_10;
wire s_105_11, s_105_12,  s_106_0,  s_106_1,  s_106_2,  s_106_3;
wire  s_106_4,  s_106_5,  s_106_6,  s_106_7,  s_106_8,  s_106_9;
wire s_106_10, s_106_11,  s_107_0,  s_107_1,  s_107_2,  s_107_3;
wire  s_107_4,  s_107_5,  s_107_6,  s_107_7,  s_107_8,  s_107_9;
wire s_107_10, s_107_11,  s_108_0,  s_108_1,  s_108_2,  s_108_3;
wire  s_108_4,  s_108_5,  s_108_6,  s_108_7,  s_108_8,  s_108_9;
wire s_108_10,  s_109_0,  s_109_1,  s_109_2,  s_109_3,  s_109_4;
wire  s_109_5,  s_109_6,  s_109_7,  s_109_8,  s_109_9, s_109_10;
wire  s_110_0,  s_110_1,  s_110_2,  s_110_3,  s_110_4,  s_110_5;
wire  s_110_6,  s_110_7,  s_110_8,  s_110_9,  s_111_0,  s_111_1;
wire  s_111_2,  s_111_3,  s_111_4,  s_111_5,  s_111_6,  s_111_7;
wire  s_111_8,  s_111_9,  s_112_0,  s_112_1,  s_112_2,  s_112_3;
wire  s_112_4,  s_112_5,  s_112_6,  s_112_7,  s_112_8,  s_113_0;
wire  s_113_1,  s_113_2,  s_113_3,  s_113_4,  s_113_5,  s_113_6;
wire  s_113_7,  s_113_8,  s_114_0,  s_114_1,  s_114_2,  s_114_3;
wire  s_114_4,  s_114_5,  s_114_6,  s_114_7,  s_115_0,  s_115_1;
wire  s_115_2,  s_115_3,  s_115_4,  s_115_5,  s_115_6,  s_115_7;
wire  s_116_0,  s_116_1,  s_116_2,  s_116_3,  s_116_4,  s_116_5;
wire  s_116_6,  s_117_0,  s_117_1,  s_117_2,  s_117_3,  s_117_4;
wire  s_117_5,  s_117_6,  s_118_0,  s_118_1,  s_118_2,  s_118_3;
wire  s_118_4,  s_118_5,  s_119_0,  s_119_1,  s_119_2,  s_119_3;
wire  s_119_4,  s_119_5,  s_120_0,  s_120_1,  s_120_2,  s_120_3;
wire  s_120_4,  s_121_0,  s_121_1,  s_121_2,  s_121_3,  s_121_4;
wire  s_122_0,  s_122_1,  s_122_2,  s_122_3,  s_123_0,  s_123_1;
wire  s_123_2,  s_123_3,  s_124_0,  s_124_1,  s_124_2,  s_125_0;
wire  s_125_1,  s_125_2,  s_126_0,  s_126_1,  s_127_0,  s_127_1;

assign {
 s_62_32,  s_60_31,  s_58_30,  s_56_29,  s_54_28,  s_52_27, 
 s_50_26,  s_48_25,  s_46_24,  s_44_23,  s_42_22,  s_40_21, 
 s_38_20,  s_36_19,  s_34_18,  s_32_17,  s_30_16,  s_28_15, 
 s_26_14,  s_24_13,  s_22_12,  s_20_11,  s_18_10,   s_16_9, 
  s_14_8,   s_12_7,   s_10_6,    s_8_5,    s_6_4,    s_4_3, 
   s_2_2,    s_0_1
} = carry;

assign {
  s_65_0,   s_64_0,   s_63_0,   s_62_0,   s_61_0,   s_60_0, 
  s_59_0,   s_58_0,   s_57_0,   s_56_0,   s_55_0,   s_54_0, 
  s_53_0,   s_52_0,   s_51_0,   s_50_0,   s_49_0,   s_48_0, 
  s_47_0,   s_46_0,   s_45_0,   s_44_0,   s_43_0,   s_42_0, 
  s_41_0,   s_40_0,   s_39_0,   s_38_0,   s_37_0,   s_36_0, 
  s_35_0,   s_34_0,   s_33_0,   s_32_0,   s_31_0,   s_30_0, 
  s_29_0,   s_28_0,   s_27_0,   s_26_0,   s_25_0,   s_24_0, 
  s_23_0,   s_22_0,   s_21_0,   s_20_0,   s_19_0,   s_18_0, 
  s_17_0,   s_16_0,   s_15_0,   s_14_0,   s_13_0,   s_12_0, 
  s_11_0,   s_10_0,    s_9_0,    s_8_0,    s_7_0,    s_6_0, 
   s_5_0,    s_4_0,    s_3_0,    s_2_0,    s_1_0,    s_0_0
} = partial_products[(width+2)*(0+1)-1:(width+2)*0];

assign {
  s_67_0,   s_66_0,   s_65_1,   s_64_1,   s_63_1,   s_62_1, 
  s_61_1,   s_60_1,   s_59_1,   s_58_1,   s_57_1,   s_56_1, 
  s_55_1,   s_54_1,   s_53_1,   s_52_1,   s_51_1,   s_50_1, 
  s_49_1,   s_48_1,   s_47_1,   s_46_1,   s_45_1,   s_44_1, 
  s_43_1,   s_42_1,   s_41_1,   s_40_1,   s_39_1,   s_38_1, 
  s_37_1,   s_36_1,   s_35_1,   s_34_1,   s_33_1,   s_32_1, 
  s_31_1,   s_30_1,   s_29_1,   s_28_1,   s_27_1,   s_26_1, 
  s_25_1,   s_24_1,   s_23_1,   s_22_1,   s_21_1,   s_20_1, 
  s_19_1,   s_18_1,   s_17_1,   s_16_1,   s_15_1,   s_14_1, 
  s_13_1,   s_12_1,   s_11_1,   s_10_1,    s_9_1,    s_8_1, 
   s_7_1,    s_6_1,    s_5_1,    s_4_1,    s_3_1,    s_2_1
} = partial_products[(width+2)*(1+1)-1:(width+2)*1];

assign {
  s_69_0,   s_68_0,   s_67_1,   s_66_1,   s_65_2,   s_64_2, 
  s_63_2,   s_62_2,   s_61_2,   s_60_2,   s_59_2,   s_58_2, 
  s_57_2,   s_56_2,   s_55_2,   s_54_2,   s_53_2,   s_52_2, 
  s_51_2,   s_50_2,   s_49_2,   s_48_2,   s_47_2,   s_46_2, 
  s_45_2,   s_44_2,   s_43_2,   s_42_2,   s_41_2,   s_40_2, 
  s_39_2,   s_38_2,   s_37_2,   s_36_2,   s_35_2,   s_34_2, 
  s_33_2,   s_32_2,   s_31_2,   s_30_2,   s_29_2,   s_28_2, 
  s_27_2,   s_26_2,   s_25_2,   s_24_2,   s_23_2,   s_22_2, 
  s_21_2,   s_20_2,   s_19_2,   s_18_2,   s_17_2,   s_16_2, 
  s_15_2,   s_14_2,   s_13_2,   s_12_2,   s_11_2,   s_10_2, 
   s_9_2,    s_8_2,    s_7_2,    s_6_2,    s_5_2,    s_4_2
} = partial_products[(width+2)*(2+1)-1:(width+2)*2];

assign {
  s_71_0,   s_70_0,   s_69_1,   s_68_1,   s_67_2,   s_66_2, 
  s_65_3,   s_64_3,   s_63_3,   s_62_3,   s_61_3,   s_60_3, 
  s_59_3,   s_58_3,   s_57_3,   s_56_3,   s_55_3,   s_54_3, 
  s_53_3,   s_52_3,   s_51_3,   s_50_3,   s_49_3,   s_48_3, 
  s_47_3,   s_46_3,   s_45_3,   s_44_3,   s_43_3,   s_42_3, 
  s_41_3,   s_40_3,   s_39_3,   s_38_3,   s_37_3,   s_36_3, 
  s_35_3,   s_34_3,   s_33_3,   s_32_3,   s_31_3,   s_30_3, 
  s_29_3,   s_28_3,   s_27_3,   s_26_3,   s_25_3,   s_24_3, 
  s_23_3,   s_22_3,   s_21_3,   s_20_3,   s_19_3,   s_18_3, 
  s_17_3,   s_16_3,   s_15_3,   s_14_3,   s_13_3,   s_12_3, 
  s_11_3,   s_10_3,    s_9_3,    s_8_3,    s_7_3,    s_6_3
} = partial_products[(width+2)*(3+1)-1:(width+2)*3];

assign {
  s_73_0,   s_72_0,   s_71_1,   s_70_1,   s_69_2,   s_68_2, 
  s_67_3,   s_66_3,   s_65_4,   s_64_4,   s_63_4,   s_62_4, 
  s_61_4,   s_60_4,   s_59_4,   s_58_4,   s_57_4,   s_56_4, 
  s_55_4,   s_54_4,   s_53_4,   s_52_4,   s_51_4,   s_50_4, 
  s_49_4,   s_48_4,   s_47_4,   s_46_4,   s_45_4,   s_44_4, 
  s_43_4,   s_42_4,   s_41_4,   s_40_4,   s_39_4,   s_38_4, 
  s_37_4,   s_36_4,   s_35_4,   s_34_4,   s_33_4,   s_32_4, 
  s_31_4,   s_30_4,   s_29_4,   s_28_4,   s_27_4,   s_26_4, 
  s_25_4,   s_24_4,   s_23_4,   s_22_4,   s_21_4,   s_20_4, 
  s_19_4,   s_18_4,   s_17_4,   s_16_4,   s_15_4,   s_14_4, 
  s_13_4,   s_12_4,   s_11_4,   s_10_4,    s_9_4,    s_8_4
} = partial_products[(width+2)*(4+1)-1:(width+2)*4];

assign {
  s_75_0,   s_74_0,   s_73_1,   s_72_1,   s_71_2,   s_70_2, 
  s_69_3,   s_68_3,   s_67_4,   s_66_4,   s_65_5,   s_64_5, 
  s_63_5,   s_62_5,   s_61_5,   s_60_5,   s_59_5,   s_58_5, 
  s_57_5,   s_56_5,   s_55_5,   s_54_5,   s_53_5,   s_52_5, 
  s_51_5,   s_50_5,   s_49_5,   s_48_5,   s_47_5,   s_46_5, 
  s_45_5,   s_44_5,   s_43_5,   s_42_5,   s_41_5,   s_40_5, 
  s_39_5,   s_38_5,   s_37_5,   s_36_5,   s_35_5,   s_34_5, 
  s_33_5,   s_32_5,   s_31_5,   s_30_5,   s_29_5,   s_28_5, 
  s_27_5,   s_26_5,   s_25_5,   s_24_5,   s_23_5,   s_22_5, 
  s_21_5,   s_20_5,   s_19_5,   s_18_5,   s_17_5,   s_16_5, 
  s_15_5,   s_14_5,   s_13_5,   s_12_5,   s_11_5,   s_10_5
} = partial_products[(width+2)*(5+1)-1:(width+2)*5];

assign {
  s_77_0,   s_76_0,   s_75_1,   s_74_1,   s_73_2,   s_72_2, 
  s_71_3,   s_70_3,   s_69_4,   s_68_4,   s_67_5,   s_66_5, 
  s_65_6,   s_64_6,   s_63_6,   s_62_6,   s_61_6,   s_60_6, 
  s_59_6,   s_58_6,   s_57_6,   s_56_6,   s_55_6,   s_54_6, 
  s_53_6,   s_52_6,   s_51_6,   s_50_6,   s_49_6,   s_48_6, 
  s_47_6,   s_46_6,   s_45_6,   s_44_6,   s_43_6,   s_42_6, 
  s_41_6,   s_40_6,   s_39_6,   s_38_6,   s_37_6,   s_36_6, 
  s_35_6,   s_34_6,   s_33_6,   s_32_6,   s_31_6,   s_30_6, 
  s_29_6,   s_28_6,   s_27_6,   s_26_6,   s_25_6,   s_24_6, 
  s_23_6,   s_22_6,   s_21_6,   s_20_6,   s_19_6,   s_18_6, 
  s_17_6,   s_16_6,   s_15_6,   s_14_6,   s_13_6,   s_12_6
} = partial_products[(width+2)*(6+1)-1:(width+2)*6];

assign {
  s_79_0,   s_78_0,   s_77_1,   s_76_1,   s_75_2,   s_74_2, 
  s_73_3,   s_72_3,   s_71_4,   s_70_4,   s_69_5,   s_68_5, 
  s_67_6,   s_66_6,   s_65_7,   s_64_7,   s_63_7,   s_62_7, 
  s_61_7,   s_60_7,   s_59_7,   s_58_7,   s_57_7,   s_56_7, 
  s_55_7,   s_54_7,   s_53_7,   s_52_7,   s_51_7,   s_50_7, 
  s_49_7,   s_48_7,   s_47_7,   s_46_7,   s_45_7,   s_44_7, 
  s_43_7,   s_42_7,   s_41_7,   s_40_7,   s_39_7,   s_38_7, 
  s_37_7,   s_36_7,   s_35_7,   s_34_7,   s_33_7,   s_32_7, 
  s_31_7,   s_30_7,   s_29_7,   s_28_7,   s_27_7,   s_26_7, 
  s_25_7,   s_24_7,   s_23_7,   s_22_7,   s_21_7,   s_20_7, 
  s_19_7,   s_18_7,   s_17_7,   s_16_7,   s_15_7,   s_14_7
} = partial_products[(width+2)*(7+1)-1:(width+2)*7];

assign {
  s_81_0,   s_80_0,   s_79_1,   s_78_1,   s_77_2,   s_76_2, 
  s_75_3,   s_74_3,   s_73_4,   s_72_4,   s_71_5,   s_70_5, 
  s_69_6,   s_68_6,   s_67_7,   s_66_7,   s_65_8,   s_64_8, 
  s_63_8,   s_62_8,   s_61_8,   s_60_8,   s_59_8,   s_58_8, 
  s_57_8,   s_56_8,   s_55_8,   s_54_8,   s_53_8,   s_52_8, 
  s_51_8,   s_50_8,   s_49_8,   s_48_8,   s_47_8,   s_46_8, 
  s_45_8,   s_44_8,   s_43_8,   s_42_8,   s_41_8,   s_40_8, 
  s_39_8,   s_38_8,   s_37_8,   s_36_8,   s_35_8,   s_34_8, 
  s_33_8,   s_32_8,   s_31_8,   s_30_8,   s_29_8,   s_28_8, 
  s_27_8,   s_26_8,   s_25_8,   s_24_8,   s_23_8,   s_22_8, 
  s_21_8,   s_20_8,   s_19_8,   s_18_8,   s_17_8,   s_16_8
} = partial_products[(width+2)*(8+1)-1:(width+2)*8];

assign {
  s_83_0,   s_82_0,   s_81_1,   s_80_1,   s_79_2,   s_78_2, 
  s_77_3,   s_76_3,   s_75_4,   s_74_4,   s_73_5,   s_72_5, 
  s_71_6,   s_70_6,   s_69_7,   s_68_7,   s_67_8,   s_66_8, 
  s_65_9,   s_64_9,   s_63_9,   s_62_9,   s_61_9,   s_60_9, 
  s_59_9,   s_58_9,   s_57_9,   s_56_9,   s_55_9,   s_54_9, 
  s_53_9,   s_52_9,   s_51_9,   s_50_9,   s_49_9,   s_48_9, 
  s_47_9,   s_46_9,   s_45_9,   s_44_9,   s_43_9,   s_42_9, 
  s_41_9,   s_40_9,   s_39_9,   s_38_9,   s_37_9,   s_36_9, 
  s_35_9,   s_34_9,   s_33_9,   s_32_9,   s_31_9,   s_30_9, 
  s_29_9,   s_28_9,   s_27_9,   s_26_9,   s_25_9,   s_24_9, 
  s_23_9,   s_22_9,   s_21_9,   s_20_9,   s_19_9,   s_18_9
} = partial_products[(width+2)*(9+1)-1:(width+2)*9];

assign {
  s_85_0,   s_84_0,   s_83_1,   s_82_1,   s_81_2,   s_80_2, 
  s_79_3,   s_78_3,   s_77_4,   s_76_4,   s_75_5,   s_74_5, 
  s_73_6,   s_72_6,   s_71_7,   s_70_7,   s_69_8,   s_68_8, 
  s_67_9,   s_66_9,  s_65_10,  s_64_10,  s_63_10,  s_62_10, 
 s_61_10,  s_60_10,  s_59_10,  s_58_10,  s_57_10,  s_56_10, 
 s_55_10,  s_54_10,  s_53_10,  s_52_10,  s_51_10,  s_50_10, 
 s_49_10,  s_48_10,  s_47_10,  s_46_10,  s_45_10,  s_44_10, 
 s_43_10,  s_42_10,  s_41_10,  s_40_10,  s_39_10,  s_38_10, 
 s_37_10,  s_36_10,  s_35_10,  s_34_10,  s_33_10,  s_32_10, 
 s_31_10,  s_30_10,  s_29_10,  s_28_10,  s_27_10,  s_26_10, 
 s_25_10,  s_24_10,  s_23_10,  s_22_10,  s_21_10,  s_20_10
} = partial_products[(width+2)*(10+1)-1:(width+2)*10];

assign {
  s_87_0,   s_86_0,   s_85_1,   s_84_1,   s_83_2,   s_82_2, 
  s_81_3,   s_80_3,   s_79_4,   s_78_4,   s_77_5,   s_76_5, 
  s_75_6,   s_74_6,   s_73_7,   s_72_7,   s_71_8,   s_70_8, 
  s_69_9,   s_68_9,  s_67_10,  s_66_10,  s_65_11,  s_64_11, 
 s_63_11,  s_62_11,  s_61_11,  s_60_11,  s_59_11,  s_58_11, 
 s_57_11,  s_56_11,  s_55_11,  s_54_11,  s_53_11,  s_52_11, 
 s_51_11,  s_50_11,  s_49_11,  s_48_11,  s_47_11,  s_46_11, 
 s_45_11,  s_44_11,  s_43_11,  s_42_11,  s_41_11,  s_40_11, 
 s_39_11,  s_38_11,  s_37_11,  s_36_11,  s_35_11,  s_34_11, 
 s_33_11,  s_32_11,  s_31_11,  s_30_11,  s_29_11,  s_28_11, 
 s_27_11,  s_26_11,  s_25_11,  s_24_11,  s_23_11,  s_22_11
} = partial_products[(width+2)*(11+1)-1:(width+2)*11];

assign {
  s_89_0,   s_88_0,   s_87_1,   s_86_1,   s_85_2,   s_84_2, 
  s_83_3,   s_82_3,   s_81_4,   s_80_4,   s_79_5,   s_78_5, 
  s_77_6,   s_76_6,   s_75_7,   s_74_7,   s_73_8,   s_72_8, 
  s_71_9,   s_70_9,  s_69_10,  s_68_10,  s_67_11,  s_66_11, 
 s_65_12,  s_64_12,  s_63_12,  s_62_12,  s_61_12,  s_60_12, 
 s_59_12,  s_58_12,  s_57_12,  s_56_12,  s_55_12,  s_54_12, 
 s_53_12,  s_52_12,  s_51_12,  s_50_12,  s_49_12,  s_48_12, 
 s_47_12,  s_46_12,  s_45_12,  s_44_12,  s_43_12,  s_42_12, 
 s_41_12,  s_40_12,  s_39_12,  s_38_12,  s_37_12,  s_36_12, 
 s_35_12,  s_34_12,  s_33_12,  s_32_12,  s_31_12,  s_30_12, 
 s_29_12,  s_28_12,  s_27_12,  s_26_12,  s_25_12,  s_24_12
} = partial_products[(width+2)*(12+1)-1:(width+2)*12];

assign {
  s_91_0,   s_90_0,   s_89_1,   s_88_1,   s_87_2,   s_86_2, 
  s_85_3,   s_84_3,   s_83_4,   s_82_4,   s_81_5,   s_80_5, 
  s_79_6,   s_78_6,   s_77_7,   s_76_7,   s_75_8,   s_74_8, 
  s_73_9,   s_72_9,  s_71_10,  s_70_10,  s_69_11,  s_68_11, 
 s_67_12,  s_66_12,  s_65_13,  s_64_13,  s_63_13,  s_62_13, 
 s_61_13,  s_60_13,  s_59_13,  s_58_13,  s_57_13,  s_56_13, 
 s_55_13,  s_54_13,  s_53_13,  s_52_13,  s_51_13,  s_50_13, 
 s_49_13,  s_48_13,  s_47_13,  s_46_13,  s_45_13,  s_44_13, 
 s_43_13,  s_42_13,  s_41_13,  s_40_13,  s_39_13,  s_38_13, 
 s_37_13,  s_36_13,  s_35_13,  s_34_13,  s_33_13,  s_32_13, 
 s_31_13,  s_30_13,  s_29_13,  s_28_13,  s_27_13,  s_26_13
} = partial_products[(width+2)*(13+1)-1:(width+2)*13];

assign {
  s_93_0,   s_92_0,   s_91_1,   s_90_1,   s_89_2,   s_88_2, 
  s_87_3,   s_86_3,   s_85_4,   s_84_4,   s_83_5,   s_82_5, 
  s_81_6,   s_80_6,   s_79_7,   s_78_7,   s_77_8,   s_76_8, 
  s_75_9,   s_74_9,  s_73_10,  s_72_10,  s_71_11,  s_70_11, 
 s_69_12,  s_68_12,  s_67_13,  s_66_13,  s_65_14,  s_64_14, 
 s_63_14,  s_62_14,  s_61_14,  s_60_14,  s_59_14,  s_58_14, 
 s_57_14,  s_56_14,  s_55_14,  s_54_14,  s_53_14,  s_52_14, 
 s_51_14,  s_50_14,  s_49_14,  s_48_14,  s_47_14,  s_46_14, 
 s_45_14,  s_44_14,  s_43_14,  s_42_14,  s_41_14,  s_40_14, 
 s_39_14,  s_38_14,  s_37_14,  s_36_14,  s_35_14,  s_34_14, 
 s_33_14,  s_32_14,  s_31_14,  s_30_14,  s_29_14,  s_28_14
} = partial_products[(width+2)*(14+1)-1:(width+2)*14];

assign {
  s_95_0,   s_94_0,   s_93_1,   s_92_1,   s_91_2,   s_90_2, 
  s_89_3,   s_88_3,   s_87_4,   s_86_4,   s_85_5,   s_84_5, 
  s_83_6,   s_82_6,   s_81_7,   s_80_7,   s_79_8,   s_78_8, 
  s_77_9,   s_76_9,  s_75_10,  s_74_10,  s_73_11,  s_72_11, 
 s_71_12,  s_70_12,  s_69_13,  s_68_13,  s_67_14,  s_66_14, 
 s_65_15,  s_64_15,  s_63_15,  s_62_15,  s_61_15,  s_60_15, 
 s_59_15,  s_58_15,  s_57_15,  s_56_15,  s_55_15,  s_54_15, 
 s_53_15,  s_52_15,  s_51_15,  s_50_15,  s_49_15,  s_48_15, 
 s_47_15,  s_46_15,  s_45_15,  s_44_15,  s_43_15,  s_42_15, 
 s_41_15,  s_40_15,  s_39_15,  s_38_15,  s_37_15,  s_36_15, 
 s_35_15,  s_34_15,  s_33_15,  s_32_15,  s_31_15,  s_30_15
} = partial_products[(width+2)*(15+1)-1:(width+2)*15];

assign {
  s_97_0,   s_96_0,   s_95_1,   s_94_1,   s_93_2,   s_92_2, 
  s_91_3,   s_90_3,   s_89_4,   s_88_4,   s_87_5,   s_86_5, 
  s_85_6,   s_84_6,   s_83_7,   s_82_7,   s_81_8,   s_80_8, 
  s_79_9,   s_78_9,  s_77_10,  s_76_10,  s_75_11,  s_74_11, 
 s_73_12,  s_72_12,  s_71_13,  s_70_13,  s_69_14,  s_68_14, 
 s_67_15,  s_66_15,  s_65_16,  s_64_16,  s_63_16,  s_62_16, 
 s_61_16,  s_60_16,  s_59_16,  s_58_16,  s_57_16,  s_56_16, 
 s_55_16,  s_54_16,  s_53_16,  s_52_16,  s_51_16,  s_50_16, 
 s_49_16,  s_48_16,  s_47_16,  s_46_16,  s_45_16,  s_44_16, 
 s_43_16,  s_42_16,  s_41_16,  s_40_16,  s_39_16,  s_38_16, 
 s_37_16,  s_36_16,  s_35_16,  s_34_16,  s_33_16,  s_32_16
} = partial_products[(width+2)*(16+1)-1:(width+2)*16];

assign {
  s_99_0,   s_98_0,   s_97_1,   s_96_1,   s_95_2,   s_94_2, 
  s_93_3,   s_92_3,   s_91_4,   s_90_4,   s_89_5,   s_88_5, 
  s_87_6,   s_86_6,   s_85_7,   s_84_7,   s_83_8,   s_82_8, 
  s_81_9,   s_80_9,  s_79_10,  s_78_10,  s_77_11,  s_76_11, 
 s_75_12,  s_74_12,  s_73_13,  s_72_13,  s_71_14,  s_70_14, 
 s_69_15,  s_68_15,  s_67_16,  s_66_16,  s_65_17,  s_64_17, 
 s_63_17,  s_62_17,  s_61_17,  s_60_17,  s_59_17,  s_58_17, 
 s_57_17,  s_56_17,  s_55_17,  s_54_17,  s_53_17,  s_52_17, 
 s_51_17,  s_50_17,  s_49_17,  s_48_17,  s_47_17,  s_46_17, 
 s_45_17,  s_44_17,  s_43_17,  s_42_17,  s_41_17,  s_40_17, 
 s_39_17,  s_38_17,  s_37_17,  s_36_17,  s_35_17,  s_34_17
} = partial_products[(width+2)*(17+1)-1:(width+2)*17];

assign {
 s_101_0,  s_100_0,   s_99_1,   s_98_1,   s_97_2,   s_96_2, 
  s_95_3,   s_94_3,   s_93_4,   s_92_4,   s_91_5,   s_90_5, 
  s_89_6,   s_88_6,   s_87_7,   s_86_7,   s_85_8,   s_84_8, 
  s_83_9,   s_82_9,  s_81_10,  s_80_10,  s_79_11,  s_78_11, 
 s_77_12,  s_76_12,  s_75_13,  s_74_13,  s_73_14,  s_72_14, 
 s_71_15,  s_70_15,  s_69_16,  s_68_16,  s_67_17,  s_66_17, 
 s_65_18,  s_64_18,  s_63_18,  s_62_18,  s_61_18,  s_60_18, 
 s_59_18,  s_58_18,  s_57_18,  s_56_18,  s_55_18,  s_54_18, 
 s_53_18,  s_52_18,  s_51_18,  s_50_18,  s_49_18,  s_48_18, 
 s_47_18,  s_46_18,  s_45_18,  s_44_18,  s_43_18,  s_42_18, 
 s_41_18,  s_40_18,  s_39_18,  s_38_18,  s_37_18,  s_36_18
} = partial_products[(width+2)*(18+1)-1:(width+2)*18];

assign {
 s_103_0,  s_102_0,  s_101_1,  s_100_1,   s_99_2,   s_98_2, 
  s_97_3,   s_96_3,   s_95_4,   s_94_4,   s_93_5,   s_92_5, 
  s_91_6,   s_90_6,   s_89_7,   s_88_7,   s_87_8,   s_86_8, 
  s_85_9,   s_84_9,  s_83_10,  s_82_10,  s_81_11,  s_80_11, 
 s_79_12,  s_78_12,  s_77_13,  s_76_13,  s_75_14,  s_74_14, 
 s_73_15,  s_72_15,  s_71_16,  s_70_16,  s_69_17,  s_68_17, 
 s_67_18,  s_66_18,  s_65_19,  s_64_19,  s_63_19,  s_62_19, 
 s_61_19,  s_60_19,  s_59_19,  s_58_19,  s_57_19,  s_56_19, 
 s_55_19,  s_54_19,  s_53_19,  s_52_19,  s_51_19,  s_50_19, 
 s_49_19,  s_48_19,  s_47_19,  s_46_19,  s_45_19,  s_44_19, 
 s_43_19,  s_42_19,  s_41_19,  s_40_19,  s_39_19,  s_38_19
} = partial_products[(width+2)*(19+1)-1:(width+2)*19];

assign {
 s_105_0,  s_104_0,  s_103_1,  s_102_1,  s_101_2,  s_100_2, 
  s_99_3,   s_98_3,   s_97_4,   s_96_4,   s_95_5,   s_94_5, 
  s_93_6,   s_92_6,   s_91_7,   s_90_7,   s_89_8,   s_88_8, 
  s_87_9,   s_86_9,  s_85_10,  s_84_10,  s_83_11,  s_82_11, 
 s_81_12,  s_80_12,  s_79_13,  s_78_13,  s_77_14,  s_76_14, 
 s_75_15,  s_74_15,  s_73_16,  s_72_16,  s_71_17,  s_70_17, 
 s_69_18,  s_68_18,  s_67_19,  s_66_19,  s_65_20,  s_64_20, 
 s_63_20,  s_62_20,  s_61_20,  s_60_20,  s_59_20,  s_58_20, 
 s_57_20,  s_56_20,  s_55_20,  s_54_20,  s_53_20,  s_52_20, 
 s_51_20,  s_50_20,  s_49_20,  s_48_20,  s_47_20,  s_46_20, 
 s_45_20,  s_44_20,  s_43_20,  s_42_20,  s_41_20,  s_40_20
} = partial_products[(width+2)*(20+1)-1:(width+2)*20];

assign {
 s_107_0,  s_106_0,  s_105_1,  s_104_1,  s_103_2,  s_102_2, 
 s_101_3,  s_100_3,   s_99_4,   s_98_4,   s_97_5,   s_96_5, 
  s_95_6,   s_94_6,   s_93_7,   s_92_7,   s_91_8,   s_90_8, 
  s_89_9,   s_88_9,  s_87_10,  s_86_10,  s_85_11,  s_84_11, 
 s_83_12,  s_82_12,  s_81_13,  s_80_13,  s_79_14,  s_78_14, 
 s_77_15,  s_76_15,  s_75_16,  s_74_16,  s_73_17,  s_72_17, 
 s_71_18,  s_70_18,  s_69_19,  s_68_19,  s_67_20,  s_66_20, 
 s_65_21,  s_64_21,  s_63_21,  s_62_21,  s_61_21,  s_60_21, 
 s_59_21,  s_58_21,  s_57_21,  s_56_21,  s_55_21,  s_54_21, 
 s_53_21,  s_52_21,  s_51_21,  s_50_21,  s_49_21,  s_48_21, 
 s_47_21,  s_46_21,  s_45_21,  s_44_21,  s_43_21,  s_42_21
} = partial_products[(width+2)*(21+1)-1:(width+2)*21];

assign {
 s_109_0,  s_108_0,  s_107_1,  s_106_1,  s_105_2,  s_104_2, 
 s_103_3,  s_102_3,  s_101_4,  s_100_4,   s_99_5,   s_98_5, 
  s_97_6,   s_96_6,   s_95_7,   s_94_7,   s_93_8,   s_92_8, 
  s_91_9,   s_90_9,  s_89_10,  s_88_10,  s_87_11,  s_86_11, 
 s_85_12,  s_84_12,  s_83_13,  s_82_13,  s_81_14,  s_80_14, 
 s_79_15,  s_78_15,  s_77_16,  s_76_16,  s_75_17,  s_74_17, 
 s_73_18,  s_72_18,  s_71_19,  s_70_19,  s_69_20,  s_68_20, 
 s_67_21,  s_66_21,  s_65_22,  s_64_22,  s_63_22,  s_62_22, 
 s_61_22,  s_60_22,  s_59_22,  s_58_22,  s_57_22,  s_56_22, 
 s_55_22,  s_54_22,  s_53_22,  s_52_22,  s_51_22,  s_50_22, 
 s_49_22,  s_48_22,  s_47_22,  s_46_22,  s_45_22,  s_44_22
} = partial_products[(width+2)*(22+1)-1:(width+2)*22];

assign {
 s_111_0,  s_110_0,  s_109_1,  s_108_1,  s_107_2,  s_106_2, 
 s_105_3,  s_104_3,  s_103_4,  s_102_4,  s_101_5,  s_100_5, 
  s_99_6,   s_98_6,   s_97_7,   s_96_7,   s_95_8,   s_94_8, 
  s_93_9,   s_92_9,  s_91_10,  s_90_10,  s_89_11,  s_88_11, 
 s_87_12,  s_86_12,  s_85_13,  s_84_13,  s_83_14,  s_82_14, 
 s_81_15,  s_80_15,  s_79_16,  s_78_16,  s_77_17,  s_76_17, 
 s_75_18,  s_74_18,  s_73_19,  s_72_19,  s_71_20,  s_70_20, 
 s_69_21,  s_68_21,  s_67_22,  s_66_22,  s_65_23,  s_64_23, 
 s_63_23,  s_62_23,  s_61_23,  s_60_23,  s_59_23,  s_58_23, 
 s_57_23,  s_56_23,  s_55_23,  s_54_23,  s_53_23,  s_52_23, 
 s_51_23,  s_50_23,  s_49_23,  s_48_23,  s_47_23,  s_46_23
} = partial_products[(width+2)*(23+1)-1:(width+2)*23];

assign {
 s_113_0,  s_112_0,  s_111_1,  s_110_1,  s_109_2,  s_108_2, 
 s_107_3,  s_106_3,  s_105_4,  s_104_4,  s_103_5,  s_102_5, 
 s_101_6,  s_100_6,   s_99_7,   s_98_7,   s_97_8,   s_96_8, 
  s_95_9,   s_94_9,  s_93_10,  s_92_10,  s_91_11,  s_90_11, 
 s_89_12,  s_88_12,  s_87_13,  s_86_13,  s_85_14,  s_84_14, 
 s_83_15,  s_82_15,  s_81_16,  s_80_16,  s_79_17,  s_78_17, 
 s_77_18,  s_76_18,  s_75_19,  s_74_19,  s_73_20,  s_72_20, 
 s_71_21,  s_70_21,  s_69_22,  s_68_22,  s_67_23,  s_66_23, 
 s_65_24,  s_64_24,  s_63_24,  s_62_24,  s_61_24,  s_60_24, 
 s_59_24,  s_58_24,  s_57_24,  s_56_24,  s_55_24,  s_54_24, 
 s_53_24,  s_52_24,  s_51_24,  s_50_24,  s_49_24,  s_48_24
} = partial_products[(width+2)*(24+1)-1:(width+2)*24];

assign {
 s_115_0,  s_114_0,  s_113_1,  s_112_1,  s_111_2,  s_110_2, 
 s_109_3,  s_108_3,  s_107_4,  s_106_4,  s_105_5,  s_104_5, 
 s_103_6,  s_102_6,  s_101_7,  s_100_7,   s_99_8,   s_98_8, 
  s_97_9,   s_96_9,  s_95_10,  s_94_10,  s_93_11,  s_92_11, 
 s_91_12,  s_90_12,  s_89_13,  s_88_13,  s_87_14,  s_86_14, 
 s_85_15,  s_84_15,  s_83_16,  s_82_16,  s_81_17,  s_80_17, 
 s_79_18,  s_78_18,  s_77_19,  s_76_19,  s_75_20,  s_74_20, 
 s_73_21,  s_72_21,  s_71_22,  s_70_22,  s_69_23,  s_68_23, 
 s_67_24,  s_66_24,  s_65_25,  s_64_25,  s_63_25,  s_62_25, 
 s_61_25,  s_60_25,  s_59_25,  s_58_25,  s_57_25,  s_56_25, 
 s_55_25,  s_54_25,  s_53_25,  s_52_25,  s_51_25,  s_50_25
} = partial_products[(width+2)*(25+1)-1:(width+2)*25];

assign {
 s_117_0,  s_116_0,  s_115_1,  s_114_1,  s_113_2,  s_112_2, 
 s_111_3,  s_110_3,  s_109_4,  s_108_4,  s_107_5,  s_106_5, 
 s_105_6,  s_104_6,  s_103_7,  s_102_7,  s_101_8,  s_100_8, 
  s_99_9,   s_98_9,  s_97_10,  s_96_10,  s_95_11,  s_94_11, 
 s_93_12,  s_92_12,  s_91_13,  s_90_13,  s_89_14,  s_88_14, 
 s_87_15,  s_86_15,  s_85_16,  s_84_16,  s_83_17,  s_82_17, 
 s_81_18,  s_80_18,  s_79_19,  s_78_19,  s_77_20,  s_76_20, 
 s_75_21,  s_74_21,  s_73_22,  s_72_22,  s_71_23,  s_70_23, 
 s_69_24,  s_68_24,  s_67_25,  s_66_25,  s_65_26,  s_64_26, 
 s_63_26,  s_62_26,  s_61_26,  s_60_26,  s_59_26,  s_58_26, 
 s_57_26,  s_56_26,  s_55_26,  s_54_26,  s_53_26,  s_52_26
} = partial_products[(width+2)*(26+1)-1:(width+2)*26];

assign {
 s_119_0,  s_118_0,  s_117_1,  s_116_1,  s_115_2,  s_114_2, 
 s_113_3,  s_112_3,  s_111_4,  s_110_4,  s_109_5,  s_108_5, 
 s_107_6,  s_106_6,  s_105_7,  s_104_7,  s_103_8,  s_102_8, 
 s_101_9,  s_100_9,  s_99_10,  s_98_10,  s_97_11,  s_96_11, 
 s_95_12,  s_94_12,  s_93_13,  s_92_13,  s_91_14,  s_90_14, 
 s_89_15,  s_88_15,  s_87_16,  s_86_16,  s_85_17,  s_84_17, 
 s_83_18,  s_82_18,  s_81_19,  s_80_19,  s_79_20,  s_78_20, 
 s_77_21,  s_76_21,  s_75_22,  s_74_22,  s_73_23,  s_72_23, 
 s_71_24,  s_70_24,  s_69_25,  s_68_25,  s_67_26,  s_66_26, 
 s_65_27,  s_64_27,  s_63_27,  s_62_27,  s_61_27,  s_60_27, 
 s_59_27,  s_58_27,  s_57_27,  s_56_27,  s_55_27,  s_54_27
} = partial_products[(width+2)*(27+1)-1:(width+2)*27];

assign {
 s_121_0,  s_120_0,  s_119_1,  s_118_1,  s_117_2,  s_116_2, 
 s_115_3,  s_114_3,  s_113_4,  s_112_4,  s_111_5,  s_110_5, 
 s_109_6,  s_108_6,  s_107_7,  s_106_7,  s_105_8,  s_104_8, 
 s_103_9,  s_102_9, s_101_10, s_100_10,  s_99_11,  s_98_11, 
 s_97_12,  s_96_12,  s_95_13,  s_94_13,  s_93_14,  s_92_14, 
 s_91_15,  s_90_15,  s_89_16,  s_88_16,  s_87_17,  s_86_17, 
 s_85_18,  s_84_18,  s_83_19,  s_82_19,  s_81_20,  s_80_20, 
 s_79_21,  s_78_21,  s_77_22,  s_76_22,  s_75_23,  s_74_23, 
 s_73_24,  s_72_24,  s_71_25,  s_70_25,  s_69_26,  s_68_26, 
 s_67_27,  s_66_27,  s_65_28,  s_64_28,  s_63_28,  s_62_28, 
 s_61_28,  s_60_28,  s_59_28,  s_58_28,  s_57_28,  s_56_28
} = partial_products[(width+2)*(28+1)-1:(width+2)*28];

assign {
 s_123_0,  s_122_0,  s_121_1,  s_120_1,  s_119_2,  s_118_2, 
 s_117_3,  s_116_3,  s_115_4,  s_114_4,  s_113_5,  s_112_5, 
 s_111_6,  s_110_6,  s_109_7,  s_108_7,  s_107_8,  s_106_8, 
 s_105_9,  s_104_9, s_103_10, s_102_10, s_101_11, s_100_11, 
 s_99_12,  s_98_12,  s_97_13,  s_96_13,  s_95_14,  s_94_14, 
 s_93_15,  s_92_15,  s_91_16,  s_90_16,  s_89_17,  s_88_17, 
 s_87_18,  s_86_18,  s_85_19,  s_84_19,  s_83_20,  s_82_20, 
 s_81_21,  s_80_21,  s_79_22,  s_78_22,  s_77_23,  s_76_23, 
 s_75_24,  s_74_24,  s_73_25,  s_72_25,  s_71_26,  s_70_26, 
 s_69_27,  s_68_27,  s_67_28,  s_66_28,  s_65_29,  s_64_29, 
 s_63_29,  s_62_29,  s_61_29,  s_60_29,  s_59_29,  s_58_29
} = partial_products[(width+2)*(29+1)-1:(width+2)*29];

assign {
 s_125_0,  s_124_0,  s_123_1,  s_122_1,  s_121_2,  s_120_2, 
 s_119_3,  s_118_3,  s_117_4,  s_116_4,  s_115_5,  s_114_5, 
 s_113_6,  s_112_6,  s_111_7,  s_110_7,  s_109_8,  s_108_8, 
 s_107_9,  s_106_9, s_105_10, s_104_10, s_103_11, s_102_11, 
s_101_12, s_100_12,  s_99_13,  s_98_13,  s_97_14,  s_96_14, 
 s_95_15,  s_94_15,  s_93_16,  s_92_16,  s_91_17,  s_90_17, 
 s_89_18,  s_88_18,  s_87_19,  s_86_19,  s_85_20,  s_84_20, 
 s_83_21,  s_82_21,  s_81_22,  s_80_22,  s_79_23,  s_78_23, 
 s_77_24,  s_76_24,  s_75_25,  s_74_25,  s_73_26,  s_72_26, 
 s_71_27,  s_70_27,  s_69_28,  s_68_28,  s_67_29,  s_66_29, 
 s_65_30,  s_64_30,  s_63_30,  s_62_30,  s_61_30,  s_60_30
} = partial_products[(width+2)*(30+1)-1:(width+2)*30];

assign {
 s_127_0,  s_126_0,  s_125_1,  s_124_1,  s_123_2,  s_122_2, 
 s_121_3,  s_120_3,  s_119_4,  s_118_4,  s_117_5,  s_116_5, 
 s_115_6,  s_114_6,  s_113_7,  s_112_7,  s_111_8,  s_110_8, 
 s_109_9,  s_108_9, s_107_10, s_106_10, s_105_11, s_104_11, 
s_103_12, s_102_12, s_101_13, s_100_13,  s_99_14,  s_98_14, 
 s_97_15,  s_96_15,  s_95_16,  s_94_16,  s_93_17,  s_92_17, 
 s_91_18,  s_90_18,  s_89_19,  s_88_19,  s_87_20,  s_86_20, 
 s_85_21,  s_84_21,  s_83_22,  s_82_22,  s_81_23,  s_80_23, 
 s_79_24,  s_78_24,  s_77_25,  s_76_25,  s_75_26,  s_74_26, 
 s_73_27,  s_72_27,  s_71_28,  s_70_28,  s_69_29,  s_68_29, 
 s_67_30,  s_66_30,  s_65_31,  s_64_31,  s_63_31,  s_62_31
} = partial_products[(width+2)*(31+1)-1:(width+2)*31];

assign {
 s_127_1,  s_126_1,  s_125_2,  s_124_2,  s_123_3,  s_122_3, 
 s_121_4,  s_120_4,  s_119_5,  s_118_5,  s_117_6,  s_116_6, 
 s_115_7,  s_114_7,  s_113_8,  s_112_8,  s_111_9,  s_110_9, 
s_109_10, s_108_10, s_107_11, s_106_11, s_105_12, s_104_12, 
s_103_13, s_102_13, s_101_14, s_100_14,  s_99_15,  s_98_15, 
 s_97_16,  s_96_16,  s_95_17,  s_94_17,  s_93_18,  s_92_18, 
 s_91_19,  s_90_19,  s_89_20,  s_88_20,  s_87_21,  s_86_21, 
 s_85_22,  s_84_22,  s_83_23,  s_82_23,  s_81_24,  s_80_24, 
 s_79_25,  s_78_25,  s_77_26,  s_76_26,  s_75_27,  s_74_27, 
 s_73_28,  s_72_28,  s_71_29,  s_70_29,  s_69_30,  s_68_30, 
 s_67_31,  s_66_31,  s_65_32,  s_64_32
} = partial_products[(width+2)*(width/2+1)-1:(width+2)*width/2+2];

/* u0_1 Output nets */
wire t_0,      t_1;
/* u1_2 Output nets */
wire t_2,      t_3;
/* u0_3 Output nets */
wire t_4,      t_5;
/* u1_4 Output nets */
wire t_6,      t_7;
/* u1_5 Output nets */
wire t_8,      t_9;
/* u2_6 Output nets */
wire t_10,     t_11,     t_12;
/* u2_7 Output nets */
wire t_13,     t_14,     t_15;
/* u2_8 Output nets */
wire t_16,     t_17,     t_18;
/* u0_9 Output nets */
wire t_19,     t_20;
/* u2_10 Output nets */
wire t_21,     t_22,     t_23;
/* u2_11 Output nets */
wire t_24,     t_25,     t_26;
/* u1_12 Output nets */
wire t_27,     t_28;
/* u2_13 Output nets */
wire t_29,     t_30,     t_31;
/* u0_14 Output nets */
wire t_32,     t_33;
/* u2_15 Output nets */
wire t_34,     t_35,     t_36;
/* u1_16 Output nets */
wire t_37,     t_38;
/* u2_17 Output nets */
wire t_39,     t_40,     t_41;
/* u1_18 Output nets */
wire t_42,     t_43;
/* u2_19 Output nets */
wire t_44,     t_45,     t_46;
/* u2_20 Output nets */
wire t_47,     t_48,     t_49;
/* u2_21 Output nets */
wire t_50,     t_51,     t_52;
/* u2_22 Output nets */
wire t_53,     t_54,     t_55;
/* u2_23 Output nets */
wire t_56,     t_57,     t_58;
/* u2_24 Output nets */
wire t_59,     t_60,     t_61;
/* u0_25 Output nets */
wire t_62,     t_63;
/* u2_26 Output nets */
wire t_64,     t_65,     t_66;
/* u2_27 Output nets */
wire t_67,     t_68,     t_69;
/* u2_28 Output nets */
wire t_70,     t_71,     t_72;
/* u2_29 Output nets */
wire t_73,     t_74,     t_75;
/* u1_30 Output nets */
wire t_76,     t_77;
/* u2_31 Output nets */
wire t_78,     t_79,     t_80;
/* u2_32 Output nets */
wire t_81,     t_82,     t_83;
/* u0_33 Output nets */
wire t_84,     t_85;
/* u2_34 Output nets */
wire t_86,     t_87,     t_88;
/* u2_35 Output nets */
wire t_89,     t_90,     t_91;
/* u1_36 Output nets */
wire t_92,     t_93;
/* u2_37 Output nets */
wire t_94,     t_95,     t_96;
/* u2_38 Output nets */
wire t_97,     t_98,     t_99;
/* u1_39 Output nets */
wire t_100,    t_101;
/* u2_40 Output nets */
wire t_102,    t_103,    t_104;
/* u2_41 Output nets */
wire t_105,    t_106,    t_107;
/* u2_42 Output nets */
wire t_108,    t_109,    t_110;
/* u2_43 Output nets */
wire t_111,    t_112,    t_113;
/* u2_44 Output nets */
wire t_114,    t_115,    t_116;
/* u2_45 Output nets */
wire t_117,    t_118,    t_119;
/* u2_46 Output nets */
wire t_120,    t_121,    t_122;
/* u2_47 Output nets */
wire t_123,    t_124,    t_125;
/* u2_48 Output nets */
wire t_126,    t_127,    t_128;
/* u0_49 Output nets */
wire t_129,    t_130;
/* u2_50 Output nets */
wire t_131,    t_132,    t_133;
/* u2_51 Output nets */
wire t_134,    t_135,    t_136;
/* u2_52 Output nets */
wire t_137,    t_138,    t_139;
/* u2_53 Output nets */
wire t_140,    t_141,    t_142;
/* u2_54 Output nets */
wire t_143,    t_144,    t_145;
/* u2_55 Output nets */
wire t_146,    t_147,    t_148;
/* u1_56 Output nets */
wire t_149,    t_150;
/* u2_57 Output nets */
wire t_151,    t_152,    t_153;
/* u2_58 Output nets */
wire t_154,    t_155,    t_156;
/* u2_59 Output nets */
wire t_157,    t_158,    t_159;
/* u0_60 Output nets */
wire t_160,    t_161;
/* u2_61 Output nets */
wire t_162,    t_163,    t_164;
/* u2_62 Output nets */
wire t_165,    t_166,    t_167;
/* u2_63 Output nets */
wire t_168,    t_169,    t_170;
/* u1_64 Output nets */
wire t_171,    t_172;
/* u2_65 Output nets */
wire t_173,    t_174,    t_175;
/* u2_66 Output nets */
wire t_176,    t_177,    t_178;
/* u2_67 Output nets */
wire t_179,    t_180,    t_181;
/* u1_68 Output nets */
wire t_182,    t_183;
/* u2_69 Output nets */
wire t_184,    t_185,    t_186;
/* u2_70 Output nets */
wire t_187,    t_188,    t_189;
/* u2_71 Output nets */
wire t_190,    t_191,    t_192;
/* u2_72 Output nets */
wire t_193,    t_194,    t_195;
/* u2_73 Output nets */
wire t_196,    t_197,    t_198;
/* u2_74 Output nets */
wire t_199,    t_200,    t_201;
/* u2_75 Output nets */
wire t_202,    t_203,    t_204;
/* u2_76 Output nets */
wire t_205,    t_206,    t_207;
/* u2_77 Output nets */
wire t_208,    t_209,    t_210;
/* u2_78 Output nets */
wire t_211,    t_212,    t_213;
/* u2_79 Output nets */
wire t_214,    t_215,    t_216;
/* u2_80 Output nets */
wire t_217,    t_218,    t_219;
/* u0_81 Output nets */
wire t_220,    t_221;
/* u2_82 Output nets */
wire t_222,    t_223,    t_224;
/* u2_83 Output nets */
wire t_225,    t_226,    t_227;
/* u2_84 Output nets */
wire t_228,    t_229,    t_230;
/* u2_85 Output nets */
wire t_231,    t_232,    t_233;
/* u2_86 Output nets */
wire t_234,    t_235,    t_236;
/* u2_87 Output nets */
wire t_237,    t_238,    t_239;
/* u2_88 Output nets */
wire t_240,    t_241,    t_242;
/* u2_89 Output nets */
wire t_243,    t_244,    t_245;
/* u1_90 Output nets */
wire t_246,    t_247;
/* u2_91 Output nets */
wire t_248,    t_249,    t_250;
/* u2_92 Output nets */
wire t_251,    t_252,    t_253;
/* u2_93 Output nets */
wire t_254,    t_255,    t_256;
/* u2_94 Output nets */
wire t_257,    t_258,    t_259;
/* u0_95 Output nets */
wire t_260,    t_261;
/* u2_96 Output nets */
wire t_262,    t_263,    t_264;
/* u2_97 Output nets */
wire t_265,    t_266,    t_267;
/* u2_98 Output nets */
wire t_268,    t_269,    t_270;
/* u2_99 Output nets */
wire t_271,    t_272,    t_273;
/* u1_100 Output nets */
wire t_274,    t_275;
/* u2_101 Output nets */
wire t_276,    t_277,    t_278;
/* u2_102 Output nets */
wire t_279,    t_280,    t_281;
/* u2_103 Output nets */
wire t_282,    t_283,    t_284;
/* u2_104 Output nets */
wire t_285,    t_286,    t_287;
/* u1_105 Output nets */
wire t_288,    t_289;
/* u2_106 Output nets */
wire t_290,    t_291,    t_292;
/* u2_107 Output nets */
wire t_293,    t_294,    t_295;
/* u2_108 Output nets */
wire t_296,    t_297,    t_298;
/* u2_109 Output nets */
wire t_299,    t_300,    t_301;
/* u2_110 Output nets */
wire t_302,    t_303,    t_304;
/* u2_111 Output nets */
wire t_305,    t_306,    t_307;
/* u2_112 Output nets */
wire t_308,    t_309,    t_310;
/* u2_113 Output nets */
wire t_311,    t_312,    t_313;
/* u2_114 Output nets */
wire t_314,    t_315,    t_316;
/* u2_115 Output nets */
wire t_317,    t_318,    t_319;
/* u2_116 Output nets */
wire t_320,    t_321,    t_322;
/* u2_117 Output nets */
wire t_323,    t_324,    t_325;
/* u2_118 Output nets */
wire t_326,    t_327,    t_328;
/* u2_119 Output nets */
wire t_329,    t_330,    t_331;
/* u2_120 Output nets */
wire t_332,    t_333,    t_334;
/* u0_121 Output nets */
wire t_335,    t_336;
/* u2_122 Output nets */
wire t_337,    t_338,    t_339;
/* u2_123 Output nets */
wire t_340,    t_341,    t_342;
/* u2_124 Output nets */
wire t_343,    t_344,    t_345;
/* u2_125 Output nets */
wire t_346,    t_347,    t_348;
/* u2_126 Output nets */
wire t_349,    t_350,    t_351;
/* u2_127 Output nets */
wire t_352,    t_353,    t_354;
/* u2_128 Output nets */
wire t_355,    t_356,    t_357;
/* u2_129 Output nets */
wire t_358,    t_359,    t_360;
/* u2_130 Output nets */
wire t_361,    t_362,    t_363;
/* u2_131 Output nets */
wire t_364,    t_365,    t_366;
/* u1_132 Output nets */
wire t_367,    t_368;
/* u2_133 Output nets */
wire t_369,    t_370,    t_371;
/* u2_134 Output nets */
wire t_372,    t_373,    t_374;
/* u2_135 Output nets */
wire t_375,    t_376,    t_377;
/* u2_136 Output nets */
wire t_378,    t_379,    t_380;
/* u2_137 Output nets */
wire t_381,    t_382,    t_383;
/* u0_138 Output nets */
wire t_384,    t_385;
/* u2_139 Output nets */
wire t_386,    t_387,    t_388;
/* u2_140 Output nets */
wire t_389,    t_390,    t_391;
/* u2_141 Output nets */
wire t_392,    t_393,    t_394;
/* u2_142 Output nets */
wire t_395,    t_396,    t_397;
/* u2_143 Output nets */
wire t_398,    t_399,    t_400;
/* u1_144 Output nets */
wire t_401,    t_402;
/* u2_145 Output nets */
wire t_403,    t_404,    t_405;
/* u2_146 Output nets */
wire t_406,    t_407,    t_408;
/* u2_147 Output nets */
wire t_409,    t_410,    t_411;
/* u2_148 Output nets */
wire t_412,    t_413,    t_414;
/* u2_149 Output nets */
wire t_415,    t_416,    t_417;
/* u1_150 Output nets */
wire t_418,    t_419;
/* u2_151 Output nets */
wire t_420,    t_421,    t_422;
/* u2_152 Output nets */
wire t_423,    t_424,    t_425;
/* u2_153 Output nets */
wire t_426,    t_427,    t_428;
/* u2_154 Output nets */
wire t_429,    t_430,    t_431;
/* u2_155 Output nets */
wire t_432,    t_433,    t_434;
/* u2_156 Output nets */
wire t_435,    t_436,    t_437;
/* u2_157 Output nets */
wire t_438,    t_439,    t_440;
/* u2_158 Output nets */
wire t_441,    t_442,    t_443;
/* u2_159 Output nets */
wire t_444,    t_445,    t_446;
/* u2_160 Output nets */
wire t_447,    t_448,    t_449;
/* u2_161 Output nets */
wire t_450,    t_451,    t_452;
/* u2_162 Output nets */
wire t_453,    t_454,    t_455;
/* u2_163 Output nets */
wire t_456,    t_457,    t_458;
/* u2_164 Output nets */
wire t_459,    t_460,    t_461;
/* u2_165 Output nets */
wire t_462,    t_463,    t_464;
/* u2_166 Output nets */
wire t_465,    t_466,    t_467;
/* u2_167 Output nets */
wire t_468,    t_469,    t_470;
/* u2_168 Output nets */
wire t_471,    t_472,    t_473;
/* u0_169 Output nets */
wire t_474,    t_475;
/* u2_170 Output nets */
wire t_476,    t_477,    t_478;
/* u2_171 Output nets */
wire t_479,    t_480,    t_481;
/* u2_172 Output nets */
wire t_482,    t_483,    t_484;
/* u2_173 Output nets */
wire t_485,    t_486,    t_487;
/* u2_174 Output nets */
wire t_488,    t_489,    t_490;
/* u2_175 Output nets */
wire t_491,    t_492,    t_493;
/* u2_176 Output nets */
wire t_494,    t_495,    t_496;
/* u2_177 Output nets */
wire t_497,    t_498,    t_499;
/* u2_178 Output nets */
wire t_500,    t_501,    t_502;
/* u2_179 Output nets */
wire t_503,    t_504,    t_505;
/* u2_180 Output nets */
wire t_506,    t_507,    t_508;
/* u2_181 Output nets */
wire t_509,    t_510,    t_511;
/* u1_182 Output nets */
wire t_512,    t_513;
/* u2_183 Output nets */
wire t_514,    t_515,    t_516;
/* u2_184 Output nets */
wire t_517,    t_518,    t_519;
/* u2_185 Output nets */
wire t_520,    t_521,    t_522;
/* u2_186 Output nets */
wire t_523,    t_524,    t_525;
/* u2_187 Output nets */
wire t_526,    t_527,    t_528;
/* u2_188 Output nets */
wire t_529,    t_530,    t_531;
/* u0_189 Output nets */
wire t_532,    t_533;
/* u2_190 Output nets */
wire t_534,    t_535,    t_536;
/* u2_191 Output nets */
wire t_537,    t_538,    t_539;
/* u2_192 Output nets */
wire t_540,    t_541,    t_542;
/* u2_193 Output nets */
wire t_543,    t_544,    t_545;
/* u2_194 Output nets */
wire t_546,    t_547,    t_548;
/* u2_195 Output nets */
wire t_549,    t_550,    t_551;
/* u1_196 Output nets */
wire t_552,    t_553;
/* u2_197 Output nets */
wire t_554,    t_555,    t_556;
/* u2_198 Output nets */
wire t_557,    t_558,    t_559;
/* u2_199 Output nets */
wire t_560,    t_561,    t_562;
/* u2_200 Output nets */
wire t_563,    t_564,    t_565;
/* u2_201 Output nets */
wire t_566,    t_567,    t_568;
/* u2_202 Output nets */
wire t_569,    t_570,    t_571;
/* u1_203 Output nets */
wire t_572,    t_573;
/* u2_204 Output nets */
wire t_574,    t_575,    t_576;
/* u2_205 Output nets */
wire t_577,    t_578,    t_579;
/* u2_206 Output nets */
wire t_580,    t_581,    t_582;
/* u2_207 Output nets */
wire t_583,    t_584,    t_585;
/* u2_208 Output nets */
wire t_586,    t_587,    t_588;
/* u2_209 Output nets */
wire t_589,    t_590,    t_591;
/* u2_210 Output nets */
wire t_592,    t_593,    t_594;
/* u2_211 Output nets */
wire t_595,    t_596,    t_597;
/* u2_212 Output nets */
wire t_598,    t_599,    t_600;
/* u2_213 Output nets */
wire t_601,    t_602,    t_603;
/* u2_214 Output nets */
wire t_604,    t_605,    t_606;
/* u2_215 Output nets */
wire t_607,    t_608,    t_609;
/* u2_216 Output nets */
wire t_610,    t_611,    t_612;
/* u2_217 Output nets */
wire t_613,    t_614,    t_615;
/* u2_218 Output nets */
wire t_616,    t_617,    t_618;
/* u2_219 Output nets */
wire t_619,    t_620,    t_621;
/* u2_220 Output nets */
wire t_622,    t_623,    t_624;
/* u2_221 Output nets */
wire t_625,    t_626,    t_627;
/* u2_222 Output nets */
wire t_628,    t_629,    t_630;
/* u2_223 Output nets */
wire t_631,    t_632,    t_633;
/* u2_224 Output nets */
wire t_634,    t_635,    t_636;
/* u0_225 Output nets */
wire t_637,    t_638;
/* u2_226 Output nets */
wire t_639,    t_640,    t_641;
/* u2_227 Output nets */
wire t_642,    t_643,    t_644;
/* u2_228 Output nets */
wire t_645,    t_646,    t_647;
/* u2_229 Output nets */
wire t_648,    t_649,    t_650;
/* u2_230 Output nets */
wire t_651,    t_652,    t_653;
/* u2_231 Output nets */
wire t_654,    t_655,    t_656;
/* u2_232 Output nets */
wire t_657,    t_658,    t_659;
/* u2_233 Output nets */
wire t_660,    t_661,    t_662;
/* u2_234 Output nets */
wire t_663,    t_664,    t_665;
/* u2_235 Output nets */
wire t_666,    t_667,    t_668;
/* u2_236 Output nets */
wire t_669,    t_670,    t_671;
/* u2_237 Output nets */
wire t_672,    t_673,    t_674;
/* u2_238 Output nets */
wire t_675,    t_676,    t_677;
/* u2_239 Output nets */
wire t_678,    t_679,    t_680;
/* u1_240 Output nets */
wire t_681,    t_682;
/* u2_241 Output nets */
wire t_683,    t_684,    t_685;
/* u2_242 Output nets */
wire t_686,    t_687,    t_688;
/* u2_243 Output nets */
wire t_689,    t_690,    t_691;
/* u2_244 Output nets */
wire t_692,    t_693,    t_694;
/* u2_245 Output nets */
wire t_695,    t_696,    t_697;
/* u2_246 Output nets */
wire t_698,    t_699,    t_700;
/* u2_247 Output nets */
wire t_701,    t_702,    t_703;
/* u0_248 Output nets */
wire t_704,    t_705;
/* u2_249 Output nets */
wire t_706,    t_707,    t_708;
/* u2_250 Output nets */
wire t_709,    t_710,    t_711;
/* u2_251 Output nets */
wire t_712,    t_713,    t_714;
/* u2_252 Output nets */
wire t_715,    t_716,    t_717;
/* u2_253 Output nets */
wire t_718,    t_719,    t_720;
/* u2_254 Output nets */
wire t_721,    t_722,    t_723;
/* u2_255 Output nets */
wire t_724,    t_725,    t_726;
/* u1_256 Output nets */
wire t_727,    t_728;
/* u2_257 Output nets */
wire t_729,    t_730,    t_731;
/* u2_258 Output nets */
wire t_732,    t_733,    t_734;
/* u2_259 Output nets */
wire t_735,    t_736,    t_737;
/* u2_260 Output nets */
wire t_738,    t_739,    t_740;
/* u2_261 Output nets */
wire t_741,    t_742,    t_743;
/* u2_262 Output nets */
wire t_744,    t_745,    t_746;
/* u2_263 Output nets */
wire t_747,    t_748,    t_749;
/* u1_264 Output nets */
wire t_750,    t_751;
/* u2_265 Output nets */
wire t_752,    t_753,    t_754;
/* u2_266 Output nets */
wire t_755,    t_756,    t_757;
/* u2_267 Output nets */
wire t_758,    t_759,    t_760;
/* u2_268 Output nets */
wire t_761,    t_762,    t_763;
/* u2_269 Output nets */
wire t_764,    t_765,    t_766;
/* u2_270 Output nets */
wire t_767,    t_768,    t_769;
/* u2_271 Output nets */
wire t_770,    t_771,    t_772;
/* u2_272 Output nets */
wire t_773,    t_774,    t_775;
/* u2_273 Output nets */
wire t_776,    t_777,    t_778;
/* u2_274 Output nets */
wire t_779,    t_780,    t_781;
/* u2_275 Output nets */
wire t_782,    t_783,    t_784;
/* u2_276 Output nets */
wire t_785,    t_786,    t_787;
/* u2_277 Output nets */
wire t_788,    t_789,    t_790;
/* u2_278 Output nets */
wire t_791,    t_792,    t_793;
/* u2_279 Output nets */
wire t_794,    t_795,    t_796;
/* u2_280 Output nets */
wire t_797,    t_798,    t_799;
/* u2_281 Output nets */
wire t_800,    t_801,    t_802;
/* u2_282 Output nets */
wire t_803,    t_804,    t_805;
/* u2_283 Output nets */
wire t_806,    t_807,    t_808;
/* u2_284 Output nets */
wire t_809,    t_810,    t_811;
/* u2_285 Output nets */
wire t_812,    t_813,    t_814;
/* u2_286 Output nets */
wire t_815,    t_816,    t_817;
/* u2_287 Output nets */
wire t_818,    t_819,    t_820;
/* u2_288 Output nets */
wire t_821,    t_822,    t_823;
/* u2_289 Output nets */
wire t_824,    t_825,    t_826;
/* u2_290 Output nets */
wire t_827,    t_828,    t_829;
/* u2_291 Output nets */
wire t_830,    t_831,    t_832;
/* u2_292 Output nets */
wire t_833,    t_834,    t_835;
/* u2_293 Output nets */
wire t_836,    t_837,    t_838;
/* u2_294 Output nets */
wire t_839,    t_840,    t_841;
/* u2_295 Output nets */
wire t_842,    t_843,    t_844;
/* u2_296 Output nets */
wire t_845,    t_846,    t_847;
/* u2_297 Output nets */
wire t_848,    t_849,    t_850;
/* u2_298 Output nets */
wire t_851,    t_852,    t_853;
/* u2_299 Output nets */
wire t_854,    t_855,    t_856;
/* u2_300 Output nets */
wire t_857,    t_858,    t_859;
/* u2_301 Output nets */
wire t_860,    t_861,    t_862;
/* u2_302 Output nets */
wire t_863,    t_864,    t_865;
/* u2_303 Output nets */
wire t_866,    t_867,    t_868;
/* u2_304 Output nets */
wire t_869,    t_870,    t_871;
/* u2_305 Output nets */
wire t_872,    t_873,    t_874;
/* u2_306 Output nets */
wire t_875,    t_876,    t_877;
/* u2_307 Output nets */
wire t_878,    t_879,    t_880;
/* u2_308 Output nets */
wire t_881,    t_882,    t_883;
/* u2_309 Output nets */
wire t_884,    t_885,    t_886;
/* u2_310 Output nets */
wire t_887,    t_888,    t_889;
/* u2_311 Output nets */
wire t_890,    t_891,    t_892;
/* u2_312 Output nets */
wire t_893,    t_894,    t_895;
/* u2_313 Output nets */
wire t_896,    t_897,    t_898;
/* u2_314 Output nets */
wire t_899,    t_900,    t_901;
/* u2_315 Output nets */
wire t_902,    t_903,    t_904;
/* u2_316 Output nets */
wire t_905,    t_906,    t_907;
/* u2_317 Output nets */
wire t_908,    t_909,    t_910;
/* u2_318 Output nets */
wire t_911,    t_912,    t_913;
/* u2_319 Output nets */
wire t_914,    t_915,    t_916;
/* u1_320 Output nets */
wire t_917,    t_918;
/* u2_321 Output nets */
wire t_919,    t_920,    t_921;
/* u2_322 Output nets */
wire t_922,    t_923,    t_924;
/* u2_323 Output nets */
wire t_925,    t_926,    t_927;
/* u2_324 Output nets */
wire t_928,    t_929,    t_930;
/* u2_325 Output nets */
wire t_931,    t_932,    t_933;
/* u2_326 Output nets */
wire t_934,    t_935,    t_936;
/* u2_327 Output nets */
wire t_937,    t_938,    t_939;
/* u1_328 Output nets */
wire t_940,    t_941;
/* u2_329 Output nets */
wire t_942,    t_943,    t_944;
/* u2_330 Output nets */
wire t_945,    t_946,    t_947;
/* u2_331 Output nets */
wire t_948,    t_949,    t_950;
/* u2_332 Output nets */
wire t_951,    t_952,    t_953;
/* u2_333 Output nets */
wire t_954,    t_955,    t_956;
/* u2_334 Output nets */
wire t_957,    t_958,    t_959;
/* u2_335 Output nets */
wire t_960,    t_961,    t_962;
/* u0_336 Output nets */
wire t_963,    t_964;
/* u2_337 Output nets */
wire t_965,    t_966,    t_967;
/* u2_338 Output nets */
wire t_968,    t_969,    t_970;
/* u2_339 Output nets */
wire t_971,    t_972,    t_973;
/* u2_340 Output nets */
wire t_974,    t_975,    t_976;
/* u2_341 Output nets */
wire t_977,    t_978,    t_979;
/* u2_342 Output nets */
wire t_980,    t_981,    t_982;
/* u2_343 Output nets */
wire t_983,    t_984,    t_985;
/* u0_344 Output nets */
wire t_986,    t_987;
/* u2_345 Output nets */
wire t_988,    t_989,    t_990;
/* u2_346 Output nets */
wire t_991,    t_992,    t_993;
/* u2_347 Output nets */
wire t_994,    t_995,    t_996;
/* u2_348 Output nets */
wire t_997,    t_998,    t_999;
/* u2_349 Output nets */
wire t_1000,   t_1001,   t_1002;
/* u2_350 Output nets */
wire t_1003,   t_1004,   t_1005;
/* u2_351 Output nets */
wire t_1006,   t_1007,   t_1008;
/* u2_352 Output nets */
wire t_1009,   t_1010,   t_1011;
/* u2_353 Output nets */
wire t_1012,   t_1013,   t_1014;
/* u2_354 Output nets */
wire t_1015,   t_1016,   t_1017;
/* u2_355 Output nets */
wire t_1018,   t_1019,   t_1020;
/* u2_356 Output nets */
wire t_1021,   t_1022,   t_1023;
/* u2_357 Output nets */
wire t_1024,   t_1025,   t_1026;
/* u2_358 Output nets */
wire t_1027,   t_1028,   t_1029;
/* u2_359 Output nets */
wire t_1030,   t_1031,   t_1032;
/* u2_360 Output nets */
wire t_1033,   t_1034,   t_1035;
/* u2_361 Output nets */
wire t_1036,   t_1037,   t_1038;
/* u2_362 Output nets */
wire t_1039,   t_1040,   t_1041;
/* u2_363 Output nets */
wire t_1042,   t_1043,   t_1044;
/* u2_364 Output nets */
wire t_1045,   t_1046,   t_1047;
/* u2_365 Output nets */
wire t_1048,   t_1049,   t_1050;
/* u2_366 Output nets */
wire t_1051,   t_1052,   t_1053;
/* u2_367 Output nets */
wire t_1054,   t_1055,   t_1056;
/* u2_368 Output nets */
wire t_1057,   t_1058,   t_1059;
/* u2_369 Output nets */
wire t_1060,   t_1061,   t_1062;
/* u2_370 Output nets */
wire t_1063,   t_1064,   t_1065;
/* u2_371 Output nets */
wire t_1066,   t_1067,   t_1068;
/* u2_372 Output nets */
wire t_1069,   t_1070,   t_1071;
/* u2_373 Output nets */
wire t_1072,   t_1073,   t_1074;
/* u2_374 Output nets */
wire t_1075,   t_1076,   t_1077;
/* u2_375 Output nets */
wire t_1078,   t_1079,   t_1080;
/* u2_376 Output nets */
wire t_1081,   t_1082,   t_1083;
/* u2_377 Output nets */
wire t_1084,   t_1085,   t_1086;
/* u2_378 Output nets */
wire t_1087,   t_1088,   t_1089;
/* u1_379 Output nets */
wire t_1090,   t_1091;
/* u2_380 Output nets */
wire t_1092,   t_1093,   t_1094;
/* u2_381 Output nets */
wire t_1095,   t_1096,   t_1097;
/* u2_382 Output nets */
wire t_1098,   t_1099,   t_1100;
/* u2_383 Output nets */
wire t_1101,   t_1102,   t_1103;
/* u2_384 Output nets */
wire t_1104,   t_1105,   t_1106;
/* u2_385 Output nets */
wire t_1107,   t_1108,   t_1109;
/* u1_386 Output nets */
wire t_1110,   t_1111;
/* u2_387 Output nets */
wire t_1112,   t_1113,   t_1114;
/* u2_388 Output nets */
wire t_1115,   t_1116,   t_1117;
/* u2_389 Output nets */
wire t_1118,   t_1119,   t_1120;
/* u2_390 Output nets */
wire t_1121,   t_1122,   t_1123;
/* u2_391 Output nets */
wire t_1124,   t_1125,   t_1126;
/* u2_392 Output nets */
wire t_1127,   t_1128,   t_1129;
/* u0_393 Output nets */
wire t_1130,   t_1131;
/* u2_394 Output nets */
wire t_1132,   t_1133,   t_1134;
/* u2_395 Output nets */
wire t_1135,   t_1136,   t_1137;
/* u2_396 Output nets */
wire t_1138,   t_1139,   t_1140;
/* u2_397 Output nets */
wire t_1141,   t_1142,   t_1143;
/* u2_398 Output nets */
wire t_1144,   t_1145,   t_1146;
/* u2_399 Output nets */
wire t_1147,   t_1148,   t_1149;
/* u0_400 Output nets */
wire t_1150,   t_1151;
/* u2_401 Output nets */
wire t_1152,   t_1153,   t_1154;
/* u2_402 Output nets */
wire t_1155,   t_1156,   t_1157;
/* u2_403 Output nets */
wire t_1158,   t_1159,   t_1160;
/* u2_404 Output nets */
wire t_1161,   t_1162,   t_1163;
/* u2_405 Output nets */
wire t_1164,   t_1165,   t_1166;
/* u2_406 Output nets */
wire t_1167,   t_1168,   t_1169;
/* u2_407 Output nets */
wire t_1170,   t_1171,   t_1172;
/* u2_408 Output nets */
wire t_1173,   t_1174,   t_1175;
/* u2_409 Output nets */
wire t_1176,   t_1177,   t_1178;
/* u2_410 Output nets */
wire t_1179,   t_1180,   t_1181;
/* u2_411 Output nets */
wire t_1182,   t_1183,   t_1184;
/* u2_412 Output nets */
wire t_1185,   t_1186,   t_1187;
/* u2_413 Output nets */
wire t_1188,   t_1189,   t_1190;
/* u2_414 Output nets */
wire t_1191,   t_1192,   t_1193;
/* u2_415 Output nets */
wire t_1194,   t_1195,   t_1196;
/* u2_416 Output nets */
wire t_1197,   t_1198,   t_1199;
/* u2_417 Output nets */
wire t_1200,   t_1201,   t_1202;
/* u2_418 Output nets */
wire t_1203,   t_1204,   t_1205;
/* u2_419 Output nets */
wire t_1206,   t_1207,   t_1208;
/* u2_420 Output nets */
wire t_1209,   t_1210,   t_1211;
/* u2_421 Output nets */
wire t_1212,   t_1213,   t_1214;
/* u2_422 Output nets */
wire t_1215,   t_1216,   t_1217;
/* u2_423 Output nets */
wire t_1218,   t_1219,   t_1220;
/* u2_424 Output nets */
wire t_1221,   t_1222,   t_1223;
/* u2_425 Output nets */
wire t_1224,   t_1225,   t_1226;
/* u2_426 Output nets */
wire t_1227,   t_1228,   t_1229;
/* u2_427 Output nets */
wire t_1230,   t_1231,   t_1232;
/* u2_428 Output nets */
wire t_1233,   t_1234,   t_1235;
/* u2_429 Output nets */
wire t_1236,   t_1237,   t_1238;
/* u1_430 Output nets */
wire t_1239,   t_1240;
/* u2_431 Output nets */
wire t_1241,   t_1242,   t_1243;
/* u2_432 Output nets */
wire t_1244,   t_1245,   t_1246;
/* u2_433 Output nets */
wire t_1247,   t_1248,   t_1249;
/* u2_434 Output nets */
wire t_1250,   t_1251,   t_1252;
/* u2_435 Output nets */
wire t_1253,   t_1254,   t_1255;
/* u1_436 Output nets */
wire t_1256,   t_1257;
/* u2_437 Output nets */
wire t_1258,   t_1259,   t_1260;
/* u2_438 Output nets */
wire t_1261,   t_1262,   t_1263;
/* u2_439 Output nets */
wire t_1264,   t_1265,   t_1266;
/* u2_440 Output nets */
wire t_1267,   t_1268,   t_1269;
/* u2_441 Output nets */
wire t_1270,   t_1271,   t_1272;
/* u0_442 Output nets */
wire t_1273,   t_1274;
/* u2_443 Output nets */
wire t_1275,   t_1276,   t_1277;
/* u2_444 Output nets */
wire t_1278,   t_1279,   t_1280;
/* u2_445 Output nets */
wire t_1281,   t_1282,   t_1283;
/* u2_446 Output nets */
wire t_1284,   t_1285,   t_1286;
/* u2_447 Output nets */
wire t_1287,   t_1288,   t_1289;
/* u0_448 Output nets */
wire t_1290,   t_1291;
/* u2_449 Output nets */
wire t_1292,   t_1293,   t_1294;
/* u2_450 Output nets */
wire t_1295,   t_1296,   t_1297;
/* u2_451 Output nets */
wire t_1298,   t_1299,   t_1300;
/* u2_452 Output nets */
wire t_1301,   t_1302,   t_1303;
/* u2_453 Output nets */
wire t_1304,   t_1305,   t_1306;
/* u2_454 Output nets */
wire t_1307,   t_1308,   t_1309;
/* u2_455 Output nets */
wire t_1310,   t_1311,   t_1312;
/* u2_456 Output nets */
wire t_1313,   t_1314,   t_1315;
/* u2_457 Output nets */
wire t_1316,   t_1317,   t_1318;
/* u2_458 Output nets */
wire t_1319,   t_1320,   t_1321;
/* u2_459 Output nets */
wire t_1322,   t_1323,   t_1324;
/* u2_460 Output nets */
wire t_1325,   t_1326,   t_1327;
/* u2_461 Output nets */
wire t_1328,   t_1329,   t_1330;
/* u2_462 Output nets */
wire t_1331,   t_1332,   t_1333;
/* u2_463 Output nets */
wire t_1334,   t_1335,   t_1336;
/* u2_464 Output nets */
wire t_1337,   t_1338,   t_1339;
/* u2_465 Output nets */
wire t_1340,   t_1341,   t_1342;
/* u2_466 Output nets */
wire t_1343,   t_1344,   t_1345;
/* u2_467 Output nets */
wire t_1346,   t_1347,   t_1348;
/* u2_468 Output nets */
wire t_1349,   t_1350,   t_1351;
/* u2_469 Output nets */
wire t_1352,   t_1353,   t_1354;
/* u2_470 Output nets */
wire t_1355,   t_1356,   t_1357;
/* u2_471 Output nets */
wire t_1358,   t_1359,   t_1360;
/* u2_472 Output nets */
wire t_1361,   t_1362,   t_1363;
/* u1_473 Output nets */
wire t_1364,   t_1365;
/* u2_474 Output nets */
wire t_1366,   t_1367,   t_1368;
/* u2_475 Output nets */
wire t_1369,   t_1370,   t_1371;
/* u2_476 Output nets */
wire t_1372,   t_1373,   t_1374;
/* u2_477 Output nets */
wire t_1375,   t_1376,   t_1377;
/* u1_478 Output nets */
wire t_1378,   t_1379;
/* u2_479 Output nets */
wire t_1380,   t_1381,   t_1382;
/* u2_480 Output nets */
wire t_1383,   t_1384,   t_1385;
/* u2_481 Output nets */
wire t_1386,   t_1387,   t_1388;
/* u2_482 Output nets */
wire t_1389,   t_1390,   t_1391;
/* u0_483 Output nets */
wire t_1392,   t_1393;
/* u2_484 Output nets */
wire t_1394,   t_1395,   t_1396;
/* u2_485 Output nets */
wire t_1397,   t_1398,   t_1399;
/* u2_486 Output nets */
wire t_1400,   t_1401,   t_1402;
/* u2_487 Output nets */
wire t_1403,   t_1404,   t_1405;
/* u0_488 Output nets */
wire t_1406,   t_1407;
/* u2_489 Output nets */
wire t_1408,   t_1409,   t_1410;
/* u2_490 Output nets */
wire t_1411,   t_1412,   t_1413;
/* u2_491 Output nets */
wire t_1414,   t_1415,   t_1416;
/* u2_492 Output nets */
wire t_1417,   t_1418,   t_1419;
/* u2_493 Output nets */
wire t_1420,   t_1421,   t_1422;
/* u2_494 Output nets */
wire t_1423,   t_1424,   t_1425;
/* u2_495 Output nets */
wire t_1426,   t_1427,   t_1428;
/* u2_496 Output nets */
wire t_1429,   t_1430,   t_1431;
/* u2_497 Output nets */
wire t_1432,   t_1433,   t_1434;
/* u2_498 Output nets */
wire t_1435,   t_1436,   t_1437;
/* u2_499 Output nets */
wire t_1438,   t_1439,   t_1440;
/* u2_500 Output nets */
wire t_1441,   t_1442,   t_1443;
/* u2_501 Output nets */
wire t_1444,   t_1445,   t_1446;
/* u2_502 Output nets */
wire t_1447,   t_1448,   t_1449;
/* u2_503 Output nets */
wire t_1450,   t_1451,   t_1452;
/* u2_504 Output nets */
wire t_1453,   t_1454,   t_1455;
/* u2_505 Output nets */
wire t_1456,   t_1457,   t_1458;
/* u2_506 Output nets */
wire t_1459,   t_1460,   t_1461;
/* u2_507 Output nets */
wire t_1462,   t_1463,   t_1464;
/* u1_508 Output nets */
wire t_1465,   t_1466;
/* u2_509 Output nets */
wire t_1467,   t_1468,   t_1469;
/* u2_510 Output nets */
wire t_1470,   t_1471,   t_1472;
/* u2_511 Output nets */
wire t_1473,   t_1474,   t_1475;
/* u1_512 Output nets */
wire t_1476,   t_1477;
/* u2_513 Output nets */
wire t_1478,   t_1479,   t_1480;
/* u2_514 Output nets */
wire t_1481,   t_1482,   t_1483;
/* u2_515 Output nets */
wire t_1484,   t_1485,   t_1486;
/* u0_516 Output nets */
wire t_1487,   t_1488;
/* u2_517 Output nets */
wire t_1489,   t_1490,   t_1491;
/* u2_518 Output nets */
wire t_1492,   t_1493,   t_1494;
/* u2_519 Output nets */
wire t_1495,   t_1496,   t_1497;
/* u0_520 Output nets */
wire t_1498,   t_1499;
/* u2_521 Output nets */
wire t_1500,   t_1501,   t_1502;
/* u2_522 Output nets */
wire t_1503,   t_1504,   t_1505;
/* u2_523 Output nets */
wire t_1506,   t_1507,   t_1508;
/* u2_524 Output nets */
wire t_1509,   t_1510,   t_1511;
/* u2_525 Output nets */
wire t_1512,   t_1513,   t_1514;
/* u2_526 Output nets */
wire t_1515,   t_1516,   t_1517;
/* u2_527 Output nets */
wire t_1518,   t_1519,   t_1520;
/* u2_528 Output nets */
wire t_1521,   t_1522,   t_1523;
/* u2_529 Output nets */
wire t_1524,   t_1525,   t_1526;
/* u2_530 Output nets */
wire t_1527,   t_1528,   t_1529;
/* u2_531 Output nets */
wire t_1530,   t_1531,   t_1532;
/* u2_532 Output nets */
wire t_1533,   t_1534,   t_1535;
/* u2_533 Output nets */
wire t_1536,   t_1537,   t_1538;
/* u2_534 Output nets */
wire t_1539,   t_1540,   t_1541;
/* u1_535 Output nets */
wire t_1542,   t_1543;
/* u2_536 Output nets */
wire t_1544,   t_1545,   t_1546;
/* u2_537 Output nets */
wire t_1547,   t_1548,   t_1549;
/* u1_538 Output nets */
wire t_1550,   t_1551;
/* u2_539 Output nets */
wire t_1552,   t_1553,   t_1554;
/* u2_540 Output nets */
wire t_1555,   t_1556,   t_1557;
/* u0_541 Output nets */
wire t_1558,   t_1559;
/* u2_542 Output nets */
wire t_1560,   t_1561,   t_1562;
/* u2_543 Output nets */
wire t_1563,   t_1564,   t_1565;
/* u0_544 Output nets */
wire t_1566,   t_1567;
/* u2_545 Output nets */
wire t_1568,   t_1569,   t_1570;
/* u2_546 Output nets */
wire t_1571,   t_1572,   t_1573;
/* u2_547 Output nets */
wire t_1574,   t_1575,   t_1576;
/* u2_548 Output nets */
wire t_1577,   t_1578,   t_1579;
/* u2_549 Output nets */
wire t_1580,   t_1581,   t_1582;
/* u2_550 Output nets */
wire t_1583,   t_1584,   t_1585;
/* u2_551 Output nets */
wire t_1586,   t_1587,   t_1588;
/* u2_552 Output nets */
wire t_1589,   t_1590,   t_1591;
/* u2_553 Output nets */
wire t_1592,   t_1593,   t_1594;
/* u1_554 Output nets */
wire t_1595,   t_1596;
/* u2_555 Output nets */
wire t_1597,   t_1598,   t_1599;
/* u1_556 Output nets */
wire t_1600,   t_1601;
/* u2_557 Output nets */
wire t_1602,   t_1603,   t_1604;
/* u0_558 Output nets */
wire t_1605,   t_1606;
/* u2_559 Output nets */
wire t_1607,   t_1608,   t_1609;
/* u0_560 Output nets */
wire t_1610,   t_1611;
/* u2_561 Output nets */
wire t_1612,   t_1613,   t_1614;
/* u2_562 Output nets */
wire t_1615,   t_1616,   t_1617;
/* u2_563 Output nets */
wire t_1618,   t_1619,   t_1620;
/* u2_564 Output nets */
wire t_1621,   t_1622,   t_1623;
/* u1_565 Output nets */
wire t_1624,   t_1625;
/* u1_566 Output nets */
wire t_1626,   t_1627;
/* u0_567 Output nets */
wire t_1628,   t_1629;
/* u0_568 Output nets */
wire t_1630;

/* compress stage 1 */
half_adder u0_1(.a(s_0_1), .b(s_0_0), .o(t_0), .cout(t_1));
compressor_3_2 u1_2(.a(s_2_2), .b(s_2_1), .cin(s_2_0), .o(t_2), .cout(t_3));
half_adder u0_3(.a(s_3_1), .b(s_3_0), .o(t_4), .cout(t_5));
compressor_3_2 u1_4(.a(s_4_2), .b(s_4_1), .cin(s_4_0), .o(t_6), .cout(t_7));
compressor_3_2 u1_5(.a(s_5_2), .b(s_5_1), .cin(s_5_0), .o(t_8), .cout(t_9));
compressor_4_2 u2_6(.a(s_6_4), .b(s_6_3), .c(s_6_2), .d(s_6_1), .cin(s_6_0), .o(t_10), .co(t_11), .cout(t_12));
compressor_4_2 u2_7(.a(s_7_3), .b(s_7_2), .c(s_7_1), .d(s_7_0), .cin(t_12), .o(t_13), .co(t_14), .cout(t_15));
compressor_4_2 u2_8(.a(s_8_3), .b(s_8_2), .c(s_8_1), .d(s_8_0), .cin(t_15), .o(t_16), .co(t_17), .cout(t_18));
half_adder u0_9(.a(s_8_5), .b(s_8_4), .o(t_19), .cout(t_20));
compressor_4_2 u2_10(.a(s_9_3), .b(s_9_2), .c(s_9_1), .d(s_9_0), .cin(t_18), .o(t_21), .co(t_22), .cout(t_23));
compressor_4_2 u2_11(.a(s_10_3), .b(s_10_2), .c(s_10_1), .d(s_10_0), .cin(t_23), .o(t_24), .co(t_25), .cout(t_26));
compressor_3_2 u1_12(.a(s_10_6), .b(s_10_5), .cin(s_10_4), .o(t_27), .cout(t_28));
compressor_4_2 u2_13(.a(s_11_3), .b(s_11_2), .c(s_11_1), .d(s_11_0), .cin(t_26), .o(t_29), .co(t_30), .cout(t_31));
half_adder u0_14(.a(s_11_5), .b(s_11_4), .o(t_32), .cout(t_33));
compressor_4_2 u2_15(.a(s_12_3), .b(s_12_2), .c(s_12_1), .d(s_12_0), .cin(t_31), .o(t_34), .co(t_35), .cout(t_36));
compressor_3_2 u1_16(.a(s_12_6), .b(s_12_5), .cin(s_12_4), .o(t_37), .cout(t_38));
compressor_4_2 u2_17(.a(s_13_3), .b(s_13_2), .c(s_13_1), .d(s_13_0), .cin(t_36), .o(t_39), .co(t_40), .cout(t_41));
compressor_3_2 u1_18(.a(s_13_6), .b(s_13_5), .cin(s_13_4), .o(t_42), .cout(t_43));
compressor_4_2 u2_19(.a(s_14_3), .b(s_14_2), .c(s_14_1), .d(s_14_0), .cin(t_41), .o(t_44), .co(t_45), .cout(t_46));
compressor_4_2 u2_20(.a(s_14_8), .b(s_14_7), .c(s_14_6), .d(s_14_5), .cin(s_14_4), .o(t_47), .co(t_48), .cout(t_49));
compressor_4_2 u2_21(.a(s_15_3), .b(s_15_2), .c(s_15_1), .d(s_15_0), .cin(t_46), .o(t_50), .co(t_51), .cout(t_52));
compressor_4_2 u2_22(.a(s_15_7), .b(s_15_6), .c(s_15_5), .d(s_15_4), .cin(t_49), .o(t_53), .co(t_54), .cout(t_55));
compressor_4_2 u2_23(.a(s_16_3), .b(s_16_2), .c(s_16_1), .d(s_16_0), .cin(t_52), .o(t_56), .co(t_57), .cout(t_58));
compressor_4_2 u2_24(.a(s_16_7), .b(s_16_6), .c(s_16_5), .d(s_16_4), .cin(t_55), .o(t_59), .co(t_60), .cout(t_61));
half_adder u0_25(.a(s_16_9), .b(s_16_8), .o(t_62), .cout(t_63));
compressor_4_2 u2_26(.a(s_17_3), .b(s_17_2), .c(s_17_1), .d(s_17_0), .cin(t_58), .o(t_64), .co(t_65), .cout(t_66));
compressor_4_2 u2_27(.a(s_17_7), .b(s_17_6), .c(s_17_5), .d(s_17_4), .cin(t_61), .o(t_67), .co(t_68), .cout(t_69));
compressor_4_2 u2_28(.a(s_18_3), .b(s_18_2), .c(s_18_1), .d(s_18_0), .cin(t_66), .o(t_70), .co(t_71), .cout(t_72));
compressor_4_2 u2_29(.a(s_18_7), .b(s_18_6), .c(s_18_5), .d(s_18_4), .cin(t_69), .o(t_73), .co(t_74), .cout(t_75));
compressor_3_2 u1_30(.a(s_18_10), .b(s_18_9), .cin(s_18_8), .o(t_76), .cout(t_77));
compressor_4_2 u2_31(.a(s_19_3), .b(s_19_2), .c(s_19_1), .d(s_19_0), .cin(t_72), .o(t_78), .co(t_79), .cout(t_80));
compressor_4_2 u2_32(.a(s_19_7), .b(s_19_6), .c(s_19_5), .d(s_19_4), .cin(t_75), .o(t_81), .co(t_82), .cout(t_83));
half_adder u0_33(.a(s_19_9), .b(s_19_8), .o(t_84), .cout(t_85));
compressor_4_2 u2_34(.a(s_20_3), .b(s_20_2), .c(s_20_1), .d(s_20_0), .cin(t_80), .o(t_86), .co(t_87), .cout(t_88));
compressor_4_2 u2_35(.a(s_20_7), .b(s_20_6), .c(s_20_5), .d(s_20_4), .cin(t_83), .o(t_89), .co(t_90), .cout(t_91));
compressor_3_2 u1_36(.a(s_20_10), .b(s_20_9), .cin(s_20_8), .o(t_92), .cout(t_93));
compressor_4_2 u2_37(.a(s_21_3), .b(s_21_2), .c(s_21_1), .d(s_21_0), .cin(t_88), .o(t_94), .co(t_95), .cout(t_96));
compressor_4_2 u2_38(.a(s_21_7), .b(s_21_6), .c(s_21_5), .d(s_21_4), .cin(t_91), .o(t_97), .co(t_98), .cout(t_99));
compressor_3_2 u1_39(.a(s_21_10), .b(s_21_9), .cin(s_21_8), .o(t_100), .cout(t_101));
compressor_4_2 u2_40(.a(s_22_3), .b(s_22_2), .c(s_22_1), .d(s_22_0), .cin(t_96), .o(t_102), .co(t_103), .cout(t_104));
compressor_4_2 u2_41(.a(s_22_7), .b(s_22_6), .c(s_22_5), .d(s_22_4), .cin(t_99), .o(t_105), .co(t_106), .cout(t_107));
compressor_4_2 u2_42(.a(s_22_12), .b(s_22_11), .c(s_22_10), .d(s_22_9), .cin(s_22_8), .o(t_108), .co(t_109), .cout(t_110));
compressor_4_2 u2_43(.a(s_23_3), .b(s_23_2), .c(s_23_1), .d(s_23_0), .cin(t_104), .o(t_111), .co(t_112), .cout(t_113));
compressor_4_2 u2_44(.a(s_23_7), .b(s_23_6), .c(s_23_5), .d(s_23_4), .cin(t_107), .o(t_114), .co(t_115), .cout(t_116));
compressor_4_2 u2_45(.a(s_23_11), .b(s_23_10), .c(s_23_9), .d(s_23_8), .cin(t_110), .o(t_117), .co(t_118), .cout(t_119));
compressor_4_2 u2_46(.a(s_24_3), .b(s_24_2), .c(s_24_1), .d(s_24_0), .cin(t_113), .o(t_120), .co(t_121), .cout(t_122));
compressor_4_2 u2_47(.a(s_24_7), .b(s_24_6), .c(s_24_5), .d(s_24_4), .cin(t_116), .o(t_123), .co(t_124), .cout(t_125));
compressor_4_2 u2_48(.a(s_24_11), .b(s_24_10), .c(s_24_9), .d(s_24_8), .cin(t_119), .o(t_126), .co(t_127), .cout(t_128));
half_adder u0_49(.a(s_24_13), .b(s_24_12), .o(t_129), .cout(t_130));
compressor_4_2 u2_50(.a(s_25_3), .b(s_25_2), .c(s_25_1), .d(s_25_0), .cin(t_122), .o(t_131), .co(t_132), .cout(t_133));
compressor_4_2 u2_51(.a(s_25_7), .b(s_25_6), .c(s_25_5), .d(s_25_4), .cin(t_125), .o(t_134), .co(t_135), .cout(t_136));
compressor_4_2 u2_52(.a(s_25_11), .b(s_25_10), .c(s_25_9), .d(s_25_8), .cin(t_128), .o(t_137), .co(t_138), .cout(t_139));
compressor_4_2 u2_53(.a(s_26_3), .b(s_26_2), .c(s_26_1), .d(s_26_0), .cin(t_133), .o(t_140), .co(t_141), .cout(t_142));
compressor_4_2 u2_54(.a(s_26_7), .b(s_26_6), .c(s_26_5), .d(s_26_4), .cin(t_136), .o(t_143), .co(t_144), .cout(t_145));
compressor_4_2 u2_55(.a(s_26_11), .b(s_26_10), .c(s_26_9), .d(s_26_8), .cin(t_139), .o(t_146), .co(t_147), .cout(t_148));
compressor_3_2 u1_56(.a(s_26_14), .b(s_26_13), .cin(s_26_12), .o(t_149), .cout(t_150));
compressor_4_2 u2_57(.a(s_27_3), .b(s_27_2), .c(s_27_1), .d(s_27_0), .cin(t_142), .o(t_151), .co(t_152), .cout(t_153));
compressor_4_2 u2_58(.a(s_27_7), .b(s_27_6), .c(s_27_5), .d(s_27_4), .cin(t_145), .o(t_154), .co(t_155), .cout(t_156));
compressor_4_2 u2_59(.a(s_27_11), .b(s_27_10), .c(s_27_9), .d(s_27_8), .cin(t_148), .o(t_157), .co(t_158), .cout(t_159));
half_adder u0_60(.a(s_27_13), .b(s_27_12), .o(t_160), .cout(t_161));
compressor_4_2 u2_61(.a(s_28_3), .b(s_28_2), .c(s_28_1), .d(s_28_0), .cin(t_153), .o(t_162), .co(t_163), .cout(t_164));
compressor_4_2 u2_62(.a(s_28_7), .b(s_28_6), .c(s_28_5), .d(s_28_4), .cin(t_156), .o(t_165), .co(t_166), .cout(t_167));
compressor_4_2 u2_63(.a(s_28_11), .b(s_28_10), .c(s_28_9), .d(s_28_8), .cin(t_159), .o(t_168), .co(t_169), .cout(t_170));
compressor_3_2 u1_64(.a(s_28_14), .b(s_28_13), .cin(s_28_12), .o(t_171), .cout(t_172));
compressor_4_2 u2_65(.a(s_29_3), .b(s_29_2), .c(s_29_1), .d(s_29_0), .cin(t_164), .o(t_173), .co(t_174), .cout(t_175));
compressor_4_2 u2_66(.a(s_29_7), .b(s_29_6), .c(s_29_5), .d(s_29_4), .cin(t_167), .o(t_176), .co(t_177), .cout(t_178));
compressor_4_2 u2_67(.a(s_29_11), .b(s_29_10), .c(s_29_9), .d(s_29_8), .cin(t_170), .o(t_179), .co(t_180), .cout(t_181));
compressor_3_2 u1_68(.a(s_29_14), .b(s_29_13), .cin(s_29_12), .o(t_182), .cout(t_183));
compressor_4_2 u2_69(.a(s_30_3), .b(s_30_2), .c(s_30_1), .d(s_30_0), .cin(t_175), .o(t_184), .co(t_185), .cout(t_186));
compressor_4_2 u2_70(.a(s_30_7), .b(s_30_6), .c(s_30_5), .d(s_30_4), .cin(t_178), .o(t_187), .co(t_188), .cout(t_189));
compressor_4_2 u2_71(.a(s_30_11), .b(s_30_10), .c(s_30_9), .d(s_30_8), .cin(t_181), .o(t_190), .co(t_191), .cout(t_192));
compressor_4_2 u2_72(.a(s_30_16), .b(s_30_15), .c(s_30_14), .d(s_30_13), .cin(s_30_12), .o(t_193), .co(t_194), .cout(t_195));
compressor_4_2 u2_73(.a(s_31_3), .b(s_31_2), .c(s_31_1), .d(s_31_0), .cin(t_186), .o(t_196), .co(t_197), .cout(t_198));
compressor_4_2 u2_74(.a(s_31_7), .b(s_31_6), .c(s_31_5), .d(s_31_4), .cin(t_189), .o(t_199), .co(t_200), .cout(t_201));
compressor_4_2 u2_75(.a(s_31_11), .b(s_31_10), .c(s_31_9), .d(s_31_8), .cin(t_192), .o(t_202), .co(t_203), .cout(t_204));
compressor_4_2 u2_76(.a(s_31_15), .b(s_31_14), .c(s_31_13), .d(s_31_12), .cin(t_195), .o(t_205), .co(t_206), .cout(t_207));
compressor_4_2 u2_77(.a(s_32_3), .b(s_32_2), .c(s_32_1), .d(s_32_0), .cin(t_198), .o(t_208), .co(t_209), .cout(t_210));
compressor_4_2 u2_78(.a(s_32_7), .b(s_32_6), .c(s_32_5), .d(s_32_4), .cin(t_201), .o(t_211), .co(t_212), .cout(t_213));
compressor_4_2 u2_79(.a(s_32_11), .b(s_32_10), .c(s_32_9), .d(s_32_8), .cin(t_204), .o(t_214), .co(t_215), .cout(t_216));
compressor_4_2 u2_80(.a(s_32_15), .b(s_32_14), .c(s_32_13), .d(s_32_12), .cin(t_207), .o(t_217), .co(t_218), .cout(t_219));
half_adder u0_81(.a(s_32_17), .b(s_32_16), .o(t_220), .cout(t_221));
compressor_4_2 u2_82(.a(s_33_3), .b(s_33_2), .c(s_33_1), .d(s_33_0), .cin(t_210), .o(t_222), .co(t_223), .cout(t_224));
compressor_4_2 u2_83(.a(s_33_7), .b(s_33_6), .c(s_33_5), .d(s_33_4), .cin(t_213), .o(t_225), .co(t_226), .cout(t_227));
compressor_4_2 u2_84(.a(s_33_11), .b(s_33_10), .c(s_33_9), .d(s_33_8), .cin(t_216), .o(t_228), .co(t_229), .cout(t_230));
compressor_4_2 u2_85(.a(s_33_15), .b(s_33_14), .c(s_33_13), .d(s_33_12), .cin(t_219), .o(t_231), .co(t_232), .cout(t_233));
compressor_4_2 u2_86(.a(s_34_3), .b(s_34_2), .c(s_34_1), .d(s_34_0), .cin(t_224), .o(t_234), .co(t_235), .cout(t_236));
compressor_4_2 u2_87(.a(s_34_7), .b(s_34_6), .c(s_34_5), .d(s_34_4), .cin(t_227), .o(t_237), .co(t_238), .cout(t_239));
compressor_4_2 u2_88(.a(s_34_11), .b(s_34_10), .c(s_34_9), .d(s_34_8), .cin(t_230), .o(t_240), .co(t_241), .cout(t_242));
compressor_4_2 u2_89(.a(s_34_15), .b(s_34_14), .c(s_34_13), .d(s_34_12), .cin(t_233), .o(t_243), .co(t_244), .cout(t_245));
compressor_3_2 u1_90(.a(s_34_18), .b(s_34_17), .cin(s_34_16), .o(t_246), .cout(t_247));
compressor_4_2 u2_91(.a(s_35_3), .b(s_35_2), .c(s_35_1), .d(s_35_0), .cin(t_236), .o(t_248), .co(t_249), .cout(t_250));
compressor_4_2 u2_92(.a(s_35_7), .b(s_35_6), .c(s_35_5), .d(s_35_4), .cin(t_239), .o(t_251), .co(t_252), .cout(t_253));
compressor_4_2 u2_93(.a(s_35_11), .b(s_35_10), .c(s_35_9), .d(s_35_8), .cin(t_242), .o(t_254), .co(t_255), .cout(t_256));
compressor_4_2 u2_94(.a(s_35_15), .b(s_35_14), .c(s_35_13), .d(s_35_12), .cin(t_245), .o(t_257), .co(t_258), .cout(t_259));
half_adder u0_95(.a(s_35_17), .b(s_35_16), .o(t_260), .cout(t_261));
compressor_4_2 u2_96(.a(s_36_3), .b(s_36_2), .c(s_36_1), .d(s_36_0), .cin(t_250), .o(t_262), .co(t_263), .cout(t_264));
compressor_4_2 u2_97(.a(s_36_7), .b(s_36_6), .c(s_36_5), .d(s_36_4), .cin(t_253), .o(t_265), .co(t_266), .cout(t_267));
compressor_4_2 u2_98(.a(s_36_11), .b(s_36_10), .c(s_36_9), .d(s_36_8), .cin(t_256), .o(t_268), .co(t_269), .cout(t_270));
compressor_4_2 u2_99(.a(s_36_15), .b(s_36_14), .c(s_36_13), .d(s_36_12), .cin(t_259), .o(t_271), .co(t_272), .cout(t_273));
compressor_3_2 u1_100(.a(s_36_18), .b(s_36_17), .cin(s_36_16), .o(t_274), .cout(t_275));
compressor_4_2 u2_101(.a(s_37_3), .b(s_37_2), .c(s_37_1), .d(s_37_0), .cin(t_264), .o(t_276), .co(t_277), .cout(t_278));
compressor_4_2 u2_102(.a(s_37_7), .b(s_37_6), .c(s_37_5), .d(s_37_4), .cin(t_267), .o(t_279), .co(t_280), .cout(t_281));
compressor_4_2 u2_103(.a(s_37_11), .b(s_37_10), .c(s_37_9), .d(s_37_8), .cin(t_270), .o(t_282), .co(t_283), .cout(t_284));
compressor_4_2 u2_104(.a(s_37_15), .b(s_37_14), .c(s_37_13), .d(s_37_12), .cin(t_273), .o(t_285), .co(t_286), .cout(t_287));
compressor_3_2 u1_105(.a(s_37_18), .b(s_37_17), .cin(s_37_16), .o(t_288), .cout(t_289));
compressor_4_2 u2_106(.a(s_38_3), .b(s_38_2), .c(s_38_1), .d(s_38_0), .cin(t_278), .o(t_290), .co(t_291), .cout(t_292));
compressor_4_2 u2_107(.a(s_38_7), .b(s_38_6), .c(s_38_5), .d(s_38_4), .cin(t_281), .o(t_293), .co(t_294), .cout(t_295));
compressor_4_2 u2_108(.a(s_38_11), .b(s_38_10), .c(s_38_9), .d(s_38_8), .cin(t_284), .o(t_296), .co(t_297), .cout(t_298));
compressor_4_2 u2_109(.a(s_38_15), .b(s_38_14), .c(s_38_13), .d(s_38_12), .cin(t_287), .o(t_299), .co(t_300), .cout(t_301));
compressor_4_2 u2_110(.a(s_38_20), .b(s_38_19), .c(s_38_18), .d(s_38_17), .cin(s_38_16), .o(t_302), .co(t_303), .cout(t_304));
compressor_4_2 u2_111(.a(s_39_3), .b(s_39_2), .c(s_39_1), .d(s_39_0), .cin(t_292), .o(t_305), .co(t_306), .cout(t_307));
compressor_4_2 u2_112(.a(s_39_7), .b(s_39_6), .c(s_39_5), .d(s_39_4), .cin(t_295), .o(t_308), .co(t_309), .cout(t_310));
compressor_4_2 u2_113(.a(s_39_11), .b(s_39_10), .c(s_39_9), .d(s_39_8), .cin(t_298), .o(t_311), .co(t_312), .cout(t_313));
compressor_4_2 u2_114(.a(s_39_15), .b(s_39_14), .c(s_39_13), .d(s_39_12), .cin(t_301), .o(t_314), .co(t_315), .cout(t_316));
compressor_4_2 u2_115(.a(s_39_19), .b(s_39_18), .c(s_39_17), .d(s_39_16), .cin(t_304), .o(t_317), .co(t_318), .cout(t_319));
compressor_4_2 u2_116(.a(s_40_3), .b(s_40_2), .c(s_40_1), .d(s_40_0), .cin(t_307), .o(t_320), .co(t_321), .cout(t_322));
compressor_4_2 u2_117(.a(s_40_7), .b(s_40_6), .c(s_40_5), .d(s_40_4), .cin(t_310), .o(t_323), .co(t_324), .cout(t_325));
compressor_4_2 u2_118(.a(s_40_11), .b(s_40_10), .c(s_40_9), .d(s_40_8), .cin(t_313), .o(t_326), .co(t_327), .cout(t_328));
compressor_4_2 u2_119(.a(s_40_15), .b(s_40_14), .c(s_40_13), .d(s_40_12), .cin(t_316), .o(t_329), .co(t_330), .cout(t_331));
compressor_4_2 u2_120(.a(s_40_19), .b(s_40_18), .c(s_40_17), .d(s_40_16), .cin(t_319), .o(t_332), .co(t_333), .cout(t_334));
half_adder u0_121(.a(s_40_21), .b(s_40_20), .o(t_335), .cout(t_336));
compressor_4_2 u2_122(.a(s_41_3), .b(s_41_2), .c(s_41_1), .d(s_41_0), .cin(t_322), .o(t_337), .co(t_338), .cout(t_339));
compressor_4_2 u2_123(.a(s_41_7), .b(s_41_6), .c(s_41_5), .d(s_41_4), .cin(t_325), .o(t_340), .co(t_341), .cout(t_342));
compressor_4_2 u2_124(.a(s_41_11), .b(s_41_10), .c(s_41_9), .d(s_41_8), .cin(t_328), .o(t_343), .co(t_344), .cout(t_345));
compressor_4_2 u2_125(.a(s_41_15), .b(s_41_14), .c(s_41_13), .d(s_41_12), .cin(t_331), .o(t_346), .co(t_347), .cout(t_348));
compressor_4_2 u2_126(.a(s_41_19), .b(s_41_18), .c(s_41_17), .d(s_41_16), .cin(t_334), .o(t_349), .co(t_350), .cout(t_351));
compressor_4_2 u2_127(.a(s_42_3), .b(s_42_2), .c(s_42_1), .d(s_42_0), .cin(t_339), .o(t_352), .co(t_353), .cout(t_354));
compressor_4_2 u2_128(.a(s_42_7), .b(s_42_6), .c(s_42_5), .d(s_42_4), .cin(t_342), .o(t_355), .co(t_356), .cout(t_357));
compressor_4_2 u2_129(.a(s_42_11), .b(s_42_10), .c(s_42_9), .d(s_42_8), .cin(t_345), .o(t_358), .co(t_359), .cout(t_360));
compressor_4_2 u2_130(.a(s_42_15), .b(s_42_14), .c(s_42_13), .d(s_42_12), .cin(t_348), .o(t_361), .co(t_362), .cout(t_363));
compressor_4_2 u2_131(.a(s_42_19), .b(s_42_18), .c(s_42_17), .d(s_42_16), .cin(t_351), .o(t_364), .co(t_365), .cout(t_366));
compressor_3_2 u1_132(.a(s_42_22), .b(s_42_21), .cin(s_42_20), .o(t_367), .cout(t_368));
compressor_4_2 u2_133(.a(s_43_3), .b(s_43_2), .c(s_43_1), .d(s_43_0), .cin(t_354), .o(t_369), .co(t_370), .cout(t_371));
compressor_4_2 u2_134(.a(s_43_7), .b(s_43_6), .c(s_43_5), .d(s_43_4), .cin(t_357), .o(t_372), .co(t_373), .cout(t_374));
compressor_4_2 u2_135(.a(s_43_11), .b(s_43_10), .c(s_43_9), .d(s_43_8), .cin(t_360), .o(t_375), .co(t_376), .cout(t_377));
compressor_4_2 u2_136(.a(s_43_15), .b(s_43_14), .c(s_43_13), .d(s_43_12), .cin(t_363), .o(t_378), .co(t_379), .cout(t_380));
compressor_4_2 u2_137(.a(s_43_19), .b(s_43_18), .c(s_43_17), .d(s_43_16), .cin(t_366), .o(t_381), .co(t_382), .cout(t_383));
half_adder u0_138(.a(s_43_21), .b(s_43_20), .o(t_384), .cout(t_385));
compressor_4_2 u2_139(.a(s_44_3), .b(s_44_2), .c(s_44_1), .d(s_44_0), .cin(t_371), .o(t_386), .co(t_387), .cout(t_388));
compressor_4_2 u2_140(.a(s_44_7), .b(s_44_6), .c(s_44_5), .d(s_44_4), .cin(t_374), .o(t_389), .co(t_390), .cout(t_391));
compressor_4_2 u2_141(.a(s_44_11), .b(s_44_10), .c(s_44_9), .d(s_44_8), .cin(t_377), .o(t_392), .co(t_393), .cout(t_394));
compressor_4_2 u2_142(.a(s_44_15), .b(s_44_14), .c(s_44_13), .d(s_44_12), .cin(t_380), .o(t_395), .co(t_396), .cout(t_397));
compressor_4_2 u2_143(.a(s_44_19), .b(s_44_18), .c(s_44_17), .d(s_44_16), .cin(t_383), .o(t_398), .co(t_399), .cout(t_400));
compressor_3_2 u1_144(.a(s_44_22), .b(s_44_21), .cin(s_44_20), .o(t_401), .cout(t_402));
compressor_4_2 u2_145(.a(s_45_3), .b(s_45_2), .c(s_45_1), .d(s_45_0), .cin(t_388), .o(t_403), .co(t_404), .cout(t_405));
compressor_4_2 u2_146(.a(s_45_7), .b(s_45_6), .c(s_45_5), .d(s_45_4), .cin(t_391), .o(t_406), .co(t_407), .cout(t_408));
compressor_4_2 u2_147(.a(s_45_11), .b(s_45_10), .c(s_45_9), .d(s_45_8), .cin(t_394), .o(t_409), .co(t_410), .cout(t_411));
compressor_4_2 u2_148(.a(s_45_15), .b(s_45_14), .c(s_45_13), .d(s_45_12), .cin(t_397), .o(t_412), .co(t_413), .cout(t_414));
compressor_4_2 u2_149(.a(s_45_19), .b(s_45_18), .c(s_45_17), .d(s_45_16), .cin(t_400), .o(t_415), .co(t_416), .cout(t_417));
compressor_3_2 u1_150(.a(s_45_22), .b(s_45_21), .cin(s_45_20), .o(t_418), .cout(t_419));
compressor_4_2 u2_151(.a(s_46_3), .b(s_46_2), .c(s_46_1), .d(s_46_0), .cin(t_405), .o(t_420), .co(t_421), .cout(t_422));
compressor_4_2 u2_152(.a(s_46_7), .b(s_46_6), .c(s_46_5), .d(s_46_4), .cin(t_408), .o(t_423), .co(t_424), .cout(t_425));
compressor_4_2 u2_153(.a(s_46_11), .b(s_46_10), .c(s_46_9), .d(s_46_8), .cin(t_411), .o(t_426), .co(t_427), .cout(t_428));
compressor_4_2 u2_154(.a(s_46_15), .b(s_46_14), .c(s_46_13), .d(s_46_12), .cin(t_414), .o(t_429), .co(t_430), .cout(t_431));
compressor_4_2 u2_155(.a(s_46_19), .b(s_46_18), .c(s_46_17), .d(s_46_16), .cin(t_417), .o(t_432), .co(t_433), .cout(t_434));
compressor_4_2 u2_156(.a(s_46_24), .b(s_46_23), .c(s_46_22), .d(s_46_21), .cin(s_46_20), .o(t_435), .co(t_436), .cout(t_437));
compressor_4_2 u2_157(.a(s_47_3), .b(s_47_2), .c(s_47_1), .d(s_47_0), .cin(t_422), .o(t_438), .co(t_439), .cout(t_440));
compressor_4_2 u2_158(.a(s_47_7), .b(s_47_6), .c(s_47_5), .d(s_47_4), .cin(t_425), .o(t_441), .co(t_442), .cout(t_443));
compressor_4_2 u2_159(.a(s_47_11), .b(s_47_10), .c(s_47_9), .d(s_47_8), .cin(t_428), .o(t_444), .co(t_445), .cout(t_446));
compressor_4_2 u2_160(.a(s_47_15), .b(s_47_14), .c(s_47_13), .d(s_47_12), .cin(t_431), .o(t_447), .co(t_448), .cout(t_449));
compressor_4_2 u2_161(.a(s_47_19), .b(s_47_18), .c(s_47_17), .d(s_47_16), .cin(t_434), .o(t_450), .co(t_451), .cout(t_452));
compressor_4_2 u2_162(.a(s_47_23), .b(s_47_22), .c(s_47_21), .d(s_47_20), .cin(t_437), .o(t_453), .co(t_454), .cout(t_455));
compressor_4_2 u2_163(.a(s_48_3), .b(s_48_2), .c(s_48_1), .d(s_48_0), .cin(t_440), .o(t_456), .co(t_457), .cout(t_458));
compressor_4_2 u2_164(.a(s_48_7), .b(s_48_6), .c(s_48_5), .d(s_48_4), .cin(t_443), .o(t_459), .co(t_460), .cout(t_461));
compressor_4_2 u2_165(.a(s_48_11), .b(s_48_10), .c(s_48_9), .d(s_48_8), .cin(t_446), .o(t_462), .co(t_463), .cout(t_464));
compressor_4_2 u2_166(.a(s_48_15), .b(s_48_14), .c(s_48_13), .d(s_48_12), .cin(t_449), .o(t_465), .co(t_466), .cout(t_467));
compressor_4_2 u2_167(.a(s_48_19), .b(s_48_18), .c(s_48_17), .d(s_48_16), .cin(t_452), .o(t_468), .co(t_469), .cout(t_470));
compressor_4_2 u2_168(.a(s_48_23), .b(s_48_22), .c(s_48_21), .d(s_48_20), .cin(t_455), .o(t_471), .co(t_472), .cout(t_473));
half_adder u0_169(.a(s_48_25), .b(s_48_24), .o(t_474), .cout(t_475));
compressor_4_2 u2_170(.a(s_49_3), .b(s_49_2), .c(s_49_1), .d(s_49_0), .cin(t_458), .o(t_476), .co(t_477), .cout(t_478));
compressor_4_2 u2_171(.a(s_49_7), .b(s_49_6), .c(s_49_5), .d(s_49_4), .cin(t_461), .o(t_479), .co(t_480), .cout(t_481));
compressor_4_2 u2_172(.a(s_49_11), .b(s_49_10), .c(s_49_9), .d(s_49_8), .cin(t_464), .o(t_482), .co(t_483), .cout(t_484));
compressor_4_2 u2_173(.a(s_49_15), .b(s_49_14), .c(s_49_13), .d(s_49_12), .cin(t_467), .o(t_485), .co(t_486), .cout(t_487));
compressor_4_2 u2_174(.a(s_49_19), .b(s_49_18), .c(s_49_17), .d(s_49_16), .cin(t_470), .o(t_488), .co(t_489), .cout(t_490));
compressor_4_2 u2_175(.a(s_49_23), .b(s_49_22), .c(s_49_21), .d(s_49_20), .cin(t_473), .o(t_491), .co(t_492), .cout(t_493));
compressor_4_2 u2_176(.a(s_50_3), .b(s_50_2), .c(s_50_1), .d(s_50_0), .cin(t_478), .o(t_494), .co(t_495), .cout(t_496));
compressor_4_2 u2_177(.a(s_50_7), .b(s_50_6), .c(s_50_5), .d(s_50_4), .cin(t_481), .o(t_497), .co(t_498), .cout(t_499));
compressor_4_2 u2_178(.a(s_50_11), .b(s_50_10), .c(s_50_9), .d(s_50_8), .cin(t_484), .o(t_500), .co(t_501), .cout(t_502));
compressor_4_2 u2_179(.a(s_50_15), .b(s_50_14), .c(s_50_13), .d(s_50_12), .cin(t_487), .o(t_503), .co(t_504), .cout(t_505));
compressor_4_2 u2_180(.a(s_50_19), .b(s_50_18), .c(s_50_17), .d(s_50_16), .cin(t_490), .o(t_506), .co(t_507), .cout(t_508));
compressor_4_2 u2_181(.a(s_50_23), .b(s_50_22), .c(s_50_21), .d(s_50_20), .cin(t_493), .o(t_509), .co(t_510), .cout(t_511));
compressor_3_2 u1_182(.a(s_50_26), .b(s_50_25), .cin(s_50_24), .o(t_512), .cout(t_513));
compressor_4_2 u2_183(.a(s_51_3), .b(s_51_2), .c(s_51_1), .d(s_51_0), .cin(t_496), .o(t_514), .co(t_515), .cout(t_516));
compressor_4_2 u2_184(.a(s_51_7), .b(s_51_6), .c(s_51_5), .d(s_51_4), .cin(t_499), .o(t_517), .co(t_518), .cout(t_519));
compressor_4_2 u2_185(.a(s_51_11), .b(s_51_10), .c(s_51_9), .d(s_51_8), .cin(t_502), .o(t_520), .co(t_521), .cout(t_522));
compressor_4_2 u2_186(.a(s_51_15), .b(s_51_14), .c(s_51_13), .d(s_51_12), .cin(t_505), .o(t_523), .co(t_524), .cout(t_525));
compressor_4_2 u2_187(.a(s_51_19), .b(s_51_18), .c(s_51_17), .d(s_51_16), .cin(t_508), .o(t_526), .co(t_527), .cout(t_528));
compressor_4_2 u2_188(.a(s_51_23), .b(s_51_22), .c(s_51_21), .d(s_51_20), .cin(t_511), .o(t_529), .co(t_530), .cout(t_531));
half_adder u0_189(.a(s_51_25), .b(s_51_24), .o(t_532), .cout(t_533));
compressor_4_2 u2_190(.a(s_52_3), .b(s_52_2), .c(s_52_1), .d(s_52_0), .cin(t_516), .o(t_534), .co(t_535), .cout(t_536));
compressor_4_2 u2_191(.a(s_52_7), .b(s_52_6), .c(s_52_5), .d(s_52_4), .cin(t_519), .o(t_537), .co(t_538), .cout(t_539));
compressor_4_2 u2_192(.a(s_52_11), .b(s_52_10), .c(s_52_9), .d(s_52_8), .cin(t_522), .o(t_540), .co(t_541), .cout(t_542));
compressor_4_2 u2_193(.a(s_52_15), .b(s_52_14), .c(s_52_13), .d(s_52_12), .cin(t_525), .o(t_543), .co(t_544), .cout(t_545));
compressor_4_2 u2_194(.a(s_52_19), .b(s_52_18), .c(s_52_17), .d(s_52_16), .cin(t_528), .o(t_546), .co(t_547), .cout(t_548));
compressor_4_2 u2_195(.a(s_52_23), .b(s_52_22), .c(s_52_21), .d(s_52_20), .cin(t_531), .o(t_549), .co(t_550), .cout(t_551));
compressor_3_2 u1_196(.a(s_52_26), .b(s_52_25), .cin(s_52_24), .o(t_552), .cout(t_553));
compressor_4_2 u2_197(.a(s_53_3), .b(s_53_2), .c(s_53_1), .d(s_53_0), .cin(t_536), .o(t_554), .co(t_555), .cout(t_556));
compressor_4_2 u2_198(.a(s_53_7), .b(s_53_6), .c(s_53_5), .d(s_53_4), .cin(t_539), .o(t_557), .co(t_558), .cout(t_559));
compressor_4_2 u2_199(.a(s_53_11), .b(s_53_10), .c(s_53_9), .d(s_53_8), .cin(t_542), .o(t_560), .co(t_561), .cout(t_562));
compressor_4_2 u2_200(.a(s_53_15), .b(s_53_14), .c(s_53_13), .d(s_53_12), .cin(t_545), .o(t_563), .co(t_564), .cout(t_565));
compressor_4_2 u2_201(.a(s_53_19), .b(s_53_18), .c(s_53_17), .d(s_53_16), .cin(t_548), .o(t_566), .co(t_567), .cout(t_568));
compressor_4_2 u2_202(.a(s_53_23), .b(s_53_22), .c(s_53_21), .d(s_53_20), .cin(t_551), .o(t_569), .co(t_570), .cout(t_571));
compressor_3_2 u1_203(.a(s_53_26), .b(s_53_25), .cin(s_53_24), .o(t_572), .cout(t_573));
compressor_4_2 u2_204(.a(s_54_3), .b(s_54_2), .c(s_54_1), .d(s_54_0), .cin(t_556), .o(t_574), .co(t_575), .cout(t_576));
compressor_4_2 u2_205(.a(s_54_7), .b(s_54_6), .c(s_54_5), .d(s_54_4), .cin(t_559), .o(t_577), .co(t_578), .cout(t_579));
compressor_4_2 u2_206(.a(s_54_11), .b(s_54_10), .c(s_54_9), .d(s_54_8), .cin(t_562), .o(t_580), .co(t_581), .cout(t_582));
compressor_4_2 u2_207(.a(s_54_15), .b(s_54_14), .c(s_54_13), .d(s_54_12), .cin(t_565), .o(t_583), .co(t_584), .cout(t_585));
compressor_4_2 u2_208(.a(s_54_19), .b(s_54_18), .c(s_54_17), .d(s_54_16), .cin(t_568), .o(t_586), .co(t_587), .cout(t_588));
compressor_4_2 u2_209(.a(s_54_23), .b(s_54_22), .c(s_54_21), .d(s_54_20), .cin(t_571), .o(t_589), .co(t_590), .cout(t_591));
compressor_4_2 u2_210(.a(s_54_28), .b(s_54_27), .c(s_54_26), .d(s_54_25), .cin(s_54_24), .o(t_592), .co(t_593), .cout(t_594));
compressor_4_2 u2_211(.a(s_55_3), .b(s_55_2), .c(s_55_1), .d(s_55_0), .cin(t_576), .o(t_595), .co(t_596), .cout(t_597));
compressor_4_2 u2_212(.a(s_55_7), .b(s_55_6), .c(s_55_5), .d(s_55_4), .cin(t_579), .o(t_598), .co(t_599), .cout(t_600));
compressor_4_2 u2_213(.a(s_55_11), .b(s_55_10), .c(s_55_9), .d(s_55_8), .cin(t_582), .o(t_601), .co(t_602), .cout(t_603));
compressor_4_2 u2_214(.a(s_55_15), .b(s_55_14), .c(s_55_13), .d(s_55_12), .cin(t_585), .o(t_604), .co(t_605), .cout(t_606));
compressor_4_2 u2_215(.a(s_55_19), .b(s_55_18), .c(s_55_17), .d(s_55_16), .cin(t_588), .o(t_607), .co(t_608), .cout(t_609));
compressor_4_2 u2_216(.a(s_55_23), .b(s_55_22), .c(s_55_21), .d(s_55_20), .cin(t_591), .o(t_610), .co(t_611), .cout(t_612));
compressor_4_2 u2_217(.a(s_55_27), .b(s_55_26), .c(s_55_25), .d(s_55_24), .cin(t_594), .o(t_613), .co(t_614), .cout(t_615));
compressor_4_2 u2_218(.a(s_56_3), .b(s_56_2), .c(s_56_1), .d(s_56_0), .cin(t_597), .o(t_616), .co(t_617), .cout(t_618));
compressor_4_2 u2_219(.a(s_56_7), .b(s_56_6), .c(s_56_5), .d(s_56_4), .cin(t_600), .o(t_619), .co(t_620), .cout(t_621));
compressor_4_2 u2_220(.a(s_56_11), .b(s_56_10), .c(s_56_9), .d(s_56_8), .cin(t_603), .o(t_622), .co(t_623), .cout(t_624));
compressor_4_2 u2_221(.a(s_56_15), .b(s_56_14), .c(s_56_13), .d(s_56_12), .cin(t_606), .o(t_625), .co(t_626), .cout(t_627));
compressor_4_2 u2_222(.a(s_56_19), .b(s_56_18), .c(s_56_17), .d(s_56_16), .cin(t_609), .o(t_628), .co(t_629), .cout(t_630));
compressor_4_2 u2_223(.a(s_56_23), .b(s_56_22), .c(s_56_21), .d(s_56_20), .cin(t_612), .o(t_631), .co(t_632), .cout(t_633));
compressor_4_2 u2_224(.a(s_56_27), .b(s_56_26), .c(s_56_25), .d(s_56_24), .cin(t_615), .o(t_634), .co(t_635), .cout(t_636));
half_adder u0_225(.a(s_56_29), .b(s_56_28), .o(t_637), .cout(t_638));
compressor_4_2 u2_226(.a(s_57_3), .b(s_57_2), .c(s_57_1), .d(s_57_0), .cin(t_618), .o(t_639), .co(t_640), .cout(t_641));
compressor_4_2 u2_227(.a(s_57_7), .b(s_57_6), .c(s_57_5), .d(s_57_4), .cin(t_621), .o(t_642), .co(t_643), .cout(t_644));
compressor_4_2 u2_228(.a(s_57_11), .b(s_57_10), .c(s_57_9), .d(s_57_8), .cin(t_624), .o(t_645), .co(t_646), .cout(t_647));
compressor_4_2 u2_229(.a(s_57_15), .b(s_57_14), .c(s_57_13), .d(s_57_12), .cin(t_627), .o(t_648), .co(t_649), .cout(t_650));
compressor_4_2 u2_230(.a(s_57_19), .b(s_57_18), .c(s_57_17), .d(s_57_16), .cin(t_630), .o(t_651), .co(t_652), .cout(t_653));
compressor_4_2 u2_231(.a(s_57_23), .b(s_57_22), .c(s_57_21), .d(s_57_20), .cin(t_633), .o(t_654), .co(t_655), .cout(t_656));
compressor_4_2 u2_232(.a(s_57_27), .b(s_57_26), .c(s_57_25), .d(s_57_24), .cin(t_636), .o(t_657), .co(t_658), .cout(t_659));
compressor_4_2 u2_233(.a(s_58_3), .b(s_58_2), .c(s_58_1), .d(s_58_0), .cin(t_641), .o(t_660), .co(t_661), .cout(t_662));
compressor_4_2 u2_234(.a(s_58_7), .b(s_58_6), .c(s_58_5), .d(s_58_4), .cin(t_644), .o(t_663), .co(t_664), .cout(t_665));
compressor_4_2 u2_235(.a(s_58_11), .b(s_58_10), .c(s_58_9), .d(s_58_8), .cin(t_647), .o(t_666), .co(t_667), .cout(t_668));
compressor_4_2 u2_236(.a(s_58_15), .b(s_58_14), .c(s_58_13), .d(s_58_12), .cin(t_650), .o(t_669), .co(t_670), .cout(t_671));
compressor_4_2 u2_237(.a(s_58_19), .b(s_58_18), .c(s_58_17), .d(s_58_16), .cin(t_653), .o(t_672), .co(t_673), .cout(t_674));
compressor_4_2 u2_238(.a(s_58_23), .b(s_58_22), .c(s_58_21), .d(s_58_20), .cin(t_656), .o(t_675), .co(t_676), .cout(t_677));
compressor_4_2 u2_239(.a(s_58_27), .b(s_58_26), .c(s_58_25), .d(s_58_24), .cin(t_659), .o(t_678), .co(t_679), .cout(t_680));
compressor_3_2 u1_240(.a(s_58_30), .b(s_58_29), .cin(s_58_28), .o(t_681), .cout(t_682));
compressor_4_2 u2_241(.a(s_59_3), .b(s_59_2), .c(s_59_1), .d(s_59_0), .cin(t_662), .o(t_683), .co(t_684), .cout(t_685));
compressor_4_2 u2_242(.a(s_59_7), .b(s_59_6), .c(s_59_5), .d(s_59_4), .cin(t_665), .o(t_686), .co(t_687), .cout(t_688));
compressor_4_2 u2_243(.a(s_59_11), .b(s_59_10), .c(s_59_9), .d(s_59_8), .cin(t_668), .o(t_689), .co(t_690), .cout(t_691));
compressor_4_2 u2_244(.a(s_59_15), .b(s_59_14), .c(s_59_13), .d(s_59_12), .cin(t_671), .o(t_692), .co(t_693), .cout(t_694));
compressor_4_2 u2_245(.a(s_59_19), .b(s_59_18), .c(s_59_17), .d(s_59_16), .cin(t_674), .o(t_695), .co(t_696), .cout(t_697));
compressor_4_2 u2_246(.a(s_59_23), .b(s_59_22), .c(s_59_21), .d(s_59_20), .cin(t_677), .o(t_698), .co(t_699), .cout(t_700));
compressor_4_2 u2_247(.a(s_59_27), .b(s_59_26), .c(s_59_25), .d(s_59_24), .cin(t_680), .o(t_701), .co(t_702), .cout(t_703));
half_adder u0_248(.a(s_59_29), .b(s_59_28), .o(t_704), .cout(t_705));
compressor_4_2 u2_249(.a(s_60_3), .b(s_60_2), .c(s_60_1), .d(s_60_0), .cin(t_685), .o(t_706), .co(t_707), .cout(t_708));
compressor_4_2 u2_250(.a(s_60_7), .b(s_60_6), .c(s_60_5), .d(s_60_4), .cin(t_688), .o(t_709), .co(t_710), .cout(t_711));
compressor_4_2 u2_251(.a(s_60_11), .b(s_60_10), .c(s_60_9), .d(s_60_8), .cin(t_691), .o(t_712), .co(t_713), .cout(t_714));
compressor_4_2 u2_252(.a(s_60_15), .b(s_60_14), .c(s_60_13), .d(s_60_12), .cin(t_694), .o(t_715), .co(t_716), .cout(t_717));
compressor_4_2 u2_253(.a(s_60_19), .b(s_60_18), .c(s_60_17), .d(s_60_16), .cin(t_697), .o(t_718), .co(t_719), .cout(t_720));
compressor_4_2 u2_254(.a(s_60_23), .b(s_60_22), .c(s_60_21), .d(s_60_20), .cin(t_700), .o(t_721), .co(t_722), .cout(t_723));
compressor_4_2 u2_255(.a(s_60_27), .b(s_60_26), .c(s_60_25), .d(s_60_24), .cin(t_703), .o(t_724), .co(t_725), .cout(t_726));
compressor_3_2 u1_256(.a(s_60_30), .b(s_60_29), .cin(s_60_28), .o(t_727), .cout(t_728));
compressor_4_2 u2_257(.a(s_61_3), .b(s_61_2), .c(s_61_1), .d(s_61_0), .cin(t_708), .o(t_729), .co(t_730), .cout(t_731));
compressor_4_2 u2_258(.a(s_61_7), .b(s_61_6), .c(s_61_5), .d(s_61_4), .cin(t_711), .o(t_732), .co(t_733), .cout(t_734));
compressor_4_2 u2_259(.a(s_61_11), .b(s_61_10), .c(s_61_9), .d(s_61_8), .cin(t_714), .o(t_735), .co(t_736), .cout(t_737));
compressor_4_2 u2_260(.a(s_61_15), .b(s_61_14), .c(s_61_13), .d(s_61_12), .cin(t_717), .o(t_738), .co(t_739), .cout(t_740));
compressor_4_2 u2_261(.a(s_61_19), .b(s_61_18), .c(s_61_17), .d(s_61_16), .cin(t_720), .o(t_741), .co(t_742), .cout(t_743));
compressor_4_2 u2_262(.a(s_61_23), .b(s_61_22), .c(s_61_21), .d(s_61_20), .cin(t_723), .o(t_744), .co(t_745), .cout(t_746));
compressor_4_2 u2_263(.a(s_61_27), .b(s_61_26), .c(s_61_25), .d(s_61_24), .cin(t_726), .o(t_747), .co(t_748), .cout(t_749));
compressor_3_2 u1_264(.a(s_61_30), .b(s_61_29), .cin(s_61_28), .o(t_750), .cout(t_751));
compressor_4_2 u2_265(.a(s_62_3), .b(s_62_2), .c(s_62_1), .d(s_62_0), .cin(t_731), .o(t_752), .co(t_753), .cout(t_754));
compressor_4_2 u2_266(.a(s_62_7), .b(s_62_6), .c(s_62_5), .d(s_62_4), .cin(t_734), .o(t_755), .co(t_756), .cout(t_757));
compressor_4_2 u2_267(.a(s_62_11), .b(s_62_10), .c(s_62_9), .d(s_62_8), .cin(t_737), .o(t_758), .co(t_759), .cout(t_760));
compressor_4_2 u2_268(.a(s_62_15), .b(s_62_14), .c(s_62_13), .d(s_62_12), .cin(t_740), .o(t_761), .co(t_762), .cout(t_763));
compressor_4_2 u2_269(.a(s_62_19), .b(s_62_18), .c(s_62_17), .d(s_62_16), .cin(t_743), .o(t_764), .co(t_765), .cout(t_766));
compressor_4_2 u2_270(.a(s_62_23), .b(s_62_22), .c(s_62_21), .d(s_62_20), .cin(t_746), .o(t_767), .co(t_768), .cout(t_769));
compressor_4_2 u2_271(.a(s_62_27), .b(s_62_26), .c(s_62_25), .d(s_62_24), .cin(t_749), .o(t_770), .co(t_771), .cout(t_772));
compressor_4_2 u2_272(.a(s_62_32), .b(s_62_31), .c(s_62_30), .d(s_62_29), .cin(s_62_28), .o(t_773), .co(t_774), .cout(t_775));
compressor_4_2 u2_273(.a(s_63_3), .b(s_63_2), .c(s_63_1), .d(s_63_0), .cin(t_754), .o(t_776), .co(t_777), .cout(t_778));
compressor_4_2 u2_274(.a(s_63_7), .b(s_63_6), .c(s_63_5), .d(s_63_4), .cin(t_757), .o(t_779), .co(t_780), .cout(t_781));
compressor_4_2 u2_275(.a(s_63_11), .b(s_63_10), .c(s_63_9), .d(s_63_8), .cin(t_760), .o(t_782), .co(t_783), .cout(t_784));
compressor_4_2 u2_276(.a(s_63_15), .b(s_63_14), .c(s_63_13), .d(s_63_12), .cin(t_763), .o(t_785), .co(t_786), .cout(t_787));
compressor_4_2 u2_277(.a(s_63_19), .b(s_63_18), .c(s_63_17), .d(s_63_16), .cin(t_766), .o(t_788), .co(t_789), .cout(t_790));
compressor_4_2 u2_278(.a(s_63_23), .b(s_63_22), .c(s_63_21), .d(s_63_20), .cin(t_769), .o(t_791), .co(t_792), .cout(t_793));
compressor_4_2 u2_279(.a(s_63_27), .b(s_63_26), .c(s_63_25), .d(s_63_24), .cin(t_772), .o(t_794), .co(t_795), .cout(t_796));
compressor_4_2 u2_280(.a(s_63_31), .b(s_63_30), .c(s_63_29), .d(s_63_28), .cin(t_775), .o(t_797), .co(t_798), .cout(t_799));
compressor_4_2 u2_281(.a(s_64_3), .b(s_64_2), .c(s_64_1), .d(s_64_0), .cin(t_778), .o(t_800), .co(t_801), .cout(t_802));
compressor_4_2 u2_282(.a(s_64_7), .b(s_64_6), .c(s_64_5), .d(s_64_4), .cin(t_781), .o(t_803), .co(t_804), .cout(t_805));
compressor_4_2 u2_283(.a(s_64_11), .b(s_64_10), .c(s_64_9), .d(s_64_8), .cin(t_784), .o(t_806), .co(t_807), .cout(t_808));
compressor_4_2 u2_284(.a(s_64_15), .b(s_64_14), .c(s_64_13), .d(s_64_12), .cin(t_787), .o(t_809), .co(t_810), .cout(t_811));
compressor_4_2 u2_285(.a(s_64_19), .b(s_64_18), .c(s_64_17), .d(s_64_16), .cin(t_790), .o(t_812), .co(t_813), .cout(t_814));
compressor_4_2 u2_286(.a(s_64_23), .b(s_64_22), .c(s_64_21), .d(s_64_20), .cin(t_793), .o(t_815), .co(t_816), .cout(t_817));
compressor_4_2 u2_287(.a(s_64_27), .b(s_64_26), .c(s_64_25), .d(s_64_24), .cin(t_796), .o(t_818), .co(t_819), .cout(t_820));
compressor_4_2 u2_288(.a(s_64_31), .b(s_64_30), .c(s_64_29), .d(s_64_28), .cin(t_799), .o(t_821), .co(t_822), .cout(t_823));
compressor_4_2 u2_289(.a(s_65_3), .b(s_65_2), .c(s_65_1), .d(s_65_0), .cin(t_802), .o(t_824), .co(t_825), .cout(t_826));
compressor_4_2 u2_290(.a(s_65_7), .b(s_65_6), .c(s_65_5), .d(s_65_4), .cin(t_805), .o(t_827), .co(t_828), .cout(t_829));
compressor_4_2 u2_291(.a(s_65_11), .b(s_65_10), .c(s_65_9), .d(s_65_8), .cin(t_808), .o(t_830), .co(t_831), .cout(t_832));
compressor_4_2 u2_292(.a(s_65_15), .b(s_65_14), .c(s_65_13), .d(s_65_12), .cin(t_811), .o(t_833), .co(t_834), .cout(t_835));
compressor_4_2 u2_293(.a(s_65_19), .b(s_65_18), .c(s_65_17), .d(s_65_16), .cin(t_814), .o(t_836), .co(t_837), .cout(t_838));
compressor_4_2 u2_294(.a(s_65_23), .b(s_65_22), .c(s_65_21), .d(s_65_20), .cin(t_817), .o(t_839), .co(t_840), .cout(t_841));
compressor_4_2 u2_295(.a(s_65_27), .b(s_65_26), .c(s_65_25), .d(s_65_24), .cin(t_820), .o(t_842), .co(t_843), .cout(t_844));
compressor_4_2 u2_296(.a(s_65_31), .b(s_65_30), .c(s_65_29), .d(s_65_28), .cin(t_823), .o(t_845), .co(t_846), .cout(t_847));
compressor_4_2 u2_297(.a(s_66_3), .b(s_66_2), .c(s_66_1), .d(s_66_0), .cin(t_826), .o(t_848), .co(t_849), .cout(t_850));
compressor_4_2 u2_298(.a(s_66_7), .b(s_66_6), .c(s_66_5), .d(s_66_4), .cin(t_829), .o(t_851), .co(t_852), .cout(t_853));
compressor_4_2 u2_299(.a(s_66_11), .b(s_66_10), .c(s_66_9), .d(s_66_8), .cin(t_832), .o(t_854), .co(t_855), .cout(t_856));
compressor_4_2 u2_300(.a(s_66_15), .b(s_66_14), .c(s_66_13), .d(s_66_12), .cin(t_835), .o(t_857), .co(t_858), .cout(t_859));
compressor_4_2 u2_301(.a(s_66_19), .b(s_66_18), .c(s_66_17), .d(s_66_16), .cin(t_838), .o(t_860), .co(t_861), .cout(t_862));
compressor_4_2 u2_302(.a(s_66_23), .b(s_66_22), .c(s_66_21), .d(s_66_20), .cin(t_841), .o(t_863), .co(t_864), .cout(t_865));
compressor_4_2 u2_303(.a(s_66_27), .b(s_66_26), .c(s_66_25), .d(s_66_24), .cin(t_844), .o(t_866), .co(t_867), .cout(t_868));
compressor_4_2 u2_304(.a(s_66_31), .b(s_66_30), .c(s_66_29), .d(s_66_28), .cin(t_847), .o(t_869), .co(t_870), .cout(t_871));
compressor_4_2 u2_305(.a(s_67_3), .b(s_67_2), .c(s_67_1), .d(s_67_0), .cin(t_850), .o(t_872), .co(t_873), .cout(t_874));
compressor_4_2 u2_306(.a(s_67_7), .b(s_67_6), .c(s_67_5), .d(s_67_4), .cin(t_853), .o(t_875), .co(t_876), .cout(t_877));
compressor_4_2 u2_307(.a(s_67_11), .b(s_67_10), .c(s_67_9), .d(s_67_8), .cin(t_856), .o(t_878), .co(t_879), .cout(t_880));
compressor_4_2 u2_308(.a(s_67_15), .b(s_67_14), .c(s_67_13), .d(s_67_12), .cin(t_859), .o(t_881), .co(t_882), .cout(t_883));
compressor_4_2 u2_309(.a(s_67_19), .b(s_67_18), .c(s_67_17), .d(s_67_16), .cin(t_862), .o(t_884), .co(t_885), .cout(t_886));
compressor_4_2 u2_310(.a(s_67_23), .b(s_67_22), .c(s_67_21), .d(s_67_20), .cin(t_865), .o(t_887), .co(t_888), .cout(t_889));
compressor_4_2 u2_311(.a(s_67_27), .b(s_67_26), .c(s_67_25), .d(s_67_24), .cin(t_868), .o(t_890), .co(t_891), .cout(t_892));
compressor_4_2 u2_312(.a(s_67_31), .b(s_67_30), .c(s_67_29), .d(s_67_28), .cin(t_871), .o(t_893), .co(t_894), .cout(t_895));
compressor_4_2 u2_313(.a(s_68_3), .b(s_68_2), .c(s_68_1), .d(s_68_0), .cin(t_874), .o(t_896), .co(t_897), .cout(t_898));
compressor_4_2 u2_314(.a(s_68_7), .b(s_68_6), .c(s_68_5), .d(s_68_4), .cin(t_877), .o(t_899), .co(t_900), .cout(t_901));
compressor_4_2 u2_315(.a(s_68_11), .b(s_68_10), .c(s_68_9), .d(s_68_8), .cin(t_880), .o(t_902), .co(t_903), .cout(t_904));
compressor_4_2 u2_316(.a(s_68_15), .b(s_68_14), .c(s_68_13), .d(s_68_12), .cin(t_883), .o(t_905), .co(t_906), .cout(t_907));
compressor_4_2 u2_317(.a(s_68_19), .b(s_68_18), .c(s_68_17), .d(s_68_16), .cin(t_886), .o(t_908), .co(t_909), .cout(t_910));
compressor_4_2 u2_318(.a(s_68_23), .b(s_68_22), .c(s_68_21), .d(s_68_20), .cin(t_889), .o(t_911), .co(t_912), .cout(t_913));
compressor_4_2 u2_319(.a(s_68_27), .b(s_68_26), .c(s_68_25), .d(s_68_24), .cin(t_892), .o(t_914), .co(t_915), .cout(t_916));
compressor_3_2 u1_320(.a(s_68_29), .b(s_68_28), .cin(t_895), .o(t_917), .cout(t_918));
compressor_4_2 u2_321(.a(s_69_3), .b(s_69_2), .c(s_69_1), .d(s_69_0), .cin(t_898), .o(t_919), .co(t_920), .cout(t_921));
compressor_4_2 u2_322(.a(s_69_7), .b(s_69_6), .c(s_69_5), .d(s_69_4), .cin(t_901), .o(t_922), .co(t_923), .cout(t_924));
compressor_4_2 u2_323(.a(s_69_11), .b(s_69_10), .c(s_69_9), .d(s_69_8), .cin(t_904), .o(t_925), .co(t_926), .cout(t_927));
compressor_4_2 u2_324(.a(s_69_15), .b(s_69_14), .c(s_69_13), .d(s_69_12), .cin(t_907), .o(t_928), .co(t_929), .cout(t_930));
compressor_4_2 u2_325(.a(s_69_19), .b(s_69_18), .c(s_69_17), .d(s_69_16), .cin(t_910), .o(t_931), .co(t_932), .cout(t_933));
compressor_4_2 u2_326(.a(s_69_23), .b(s_69_22), .c(s_69_21), .d(s_69_20), .cin(t_913), .o(t_934), .co(t_935), .cout(t_936));
compressor_4_2 u2_327(.a(s_69_27), .b(s_69_26), .c(s_69_25), .d(s_69_24), .cin(t_916), .o(t_937), .co(t_938), .cout(t_939));
compressor_3_2 u1_328(.a(s_69_30), .b(s_69_29), .cin(s_69_28), .o(t_940), .cout(t_941));
compressor_4_2 u2_329(.a(s_70_3), .b(s_70_2), .c(s_70_1), .d(s_70_0), .cin(t_921), .o(t_942), .co(t_943), .cout(t_944));
compressor_4_2 u2_330(.a(s_70_7), .b(s_70_6), .c(s_70_5), .d(s_70_4), .cin(t_924), .o(t_945), .co(t_946), .cout(t_947));
compressor_4_2 u2_331(.a(s_70_11), .b(s_70_10), .c(s_70_9), .d(s_70_8), .cin(t_927), .o(t_948), .co(t_949), .cout(t_950));
compressor_4_2 u2_332(.a(s_70_15), .b(s_70_14), .c(s_70_13), .d(s_70_12), .cin(t_930), .o(t_951), .co(t_952), .cout(t_953));
compressor_4_2 u2_333(.a(s_70_19), .b(s_70_18), .c(s_70_17), .d(s_70_16), .cin(t_933), .o(t_954), .co(t_955), .cout(t_956));
compressor_4_2 u2_334(.a(s_70_23), .b(s_70_22), .c(s_70_21), .d(s_70_20), .cin(t_936), .o(t_957), .co(t_958), .cout(t_959));
compressor_4_2 u2_335(.a(s_70_27), .b(s_70_26), .c(s_70_25), .d(s_70_24), .cin(t_939), .o(t_960), .co(t_961), .cout(t_962));
half_adder u0_336(.a(s_70_29), .b(s_70_28), .o(t_963), .cout(t_964));
compressor_4_2 u2_337(.a(s_71_3), .b(s_71_2), .c(s_71_1), .d(s_71_0), .cin(t_944), .o(t_965), .co(t_966), .cout(t_967));
compressor_4_2 u2_338(.a(s_71_7), .b(s_71_6), .c(s_71_5), .d(s_71_4), .cin(t_947), .o(t_968), .co(t_969), .cout(t_970));
compressor_4_2 u2_339(.a(s_71_11), .b(s_71_10), .c(s_71_9), .d(s_71_8), .cin(t_950), .o(t_971), .co(t_972), .cout(t_973));
compressor_4_2 u2_340(.a(s_71_15), .b(s_71_14), .c(s_71_13), .d(s_71_12), .cin(t_953), .o(t_974), .co(t_975), .cout(t_976));
compressor_4_2 u2_341(.a(s_71_19), .b(s_71_18), .c(s_71_17), .d(s_71_16), .cin(t_956), .o(t_977), .co(t_978), .cout(t_979));
compressor_4_2 u2_342(.a(s_71_23), .b(s_71_22), .c(s_71_21), .d(s_71_20), .cin(t_959), .o(t_980), .co(t_981), .cout(t_982));
compressor_4_2 u2_343(.a(s_71_27), .b(s_71_26), .c(s_71_25), .d(s_71_24), .cin(t_962), .o(t_983), .co(t_984), .cout(t_985));
half_adder u0_344(.a(s_71_29), .b(s_71_28), .o(t_986), .cout(t_987));
compressor_4_2 u2_345(.a(s_72_3), .b(s_72_2), .c(s_72_1), .d(s_72_0), .cin(t_967), .o(t_988), .co(t_989), .cout(t_990));
compressor_4_2 u2_346(.a(s_72_7), .b(s_72_6), .c(s_72_5), .d(s_72_4), .cin(t_970), .o(t_991), .co(t_992), .cout(t_993));
compressor_4_2 u2_347(.a(s_72_11), .b(s_72_10), .c(s_72_9), .d(s_72_8), .cin(t_973), .o(t_994), .co(t_995), .cout(t_996));
compressor_4_2 u2_348(.a(s_72_15), .b(s_72_14), .c(s_72_13), .d(s_72_12), .cin(t_976), .o(t_997), .co(t_998), .cout(t_999));
compressor_4_2 u2_349(.a(s_72_19), .b(s_72_18), .c(s_72_17), .d(s_72_16), .cin(t_979), .o(t_1000), .co(t_1001), .cout(t_1002));
compressor_4_2 u2_350(.a(s_72_23), .b(s_72_22), .c(s_72_21), .d(s_72_20), .cin(t_982), .o(t_1003), .co(t_1004), .cout(t_1005));
compressor_4_2 u2_351(.a(s_72_27), .b(s_72_26), .c(s_72_25), .d(s_72_24), .cin(t_985), .o(t_1006), .co(t_1007), .cout(t_1008));
compressor_4_2 u2_352(.a(s_73_3), .b(s_73_2), .c(s_73_1), .d(s_73_0), .cin(t_990), .o(t_1009), .co(t_1010), .cout(t_1011));
compressor_4_2 u2_353(.a(s_73_7), .b(s_73_6), .c(s_73_5), .d(s_73_4), .cin(t_993), .o(t_1012), .co(t_1013), .cout(t_1014));
compressor_4_2 u2_354(.a(s_73_11), .b(s_73_10), .c(s_73_9), .d(s_73_8), .cin(t_996), .o(t_1015), .co(t_1016), .cout(t_1017));
compressor_4_2 u2_355(.a(s_73_15), .b(s_73_14), .c(s_73_13), .d(s_73_12), .cin(t_999), .o(t_1018), .co(t_1019), .cout(t_1020));
compressor_4_2 u2_356(.a(s_73_19), .b(s_73_18), .c(s_73_17), .d(s_73_16), .cin(t_1002), .o(t_1021), .co(t_1022), .cout(t_1023));
compressor_4_2 u2_357(.a(s_73_23), .b(s_73_22), .c(s_73_21), .d(s_73_20), .cin(t_1005), .o(t_1024), .co(t_1025), .cout(t_1026));
compressor_4_2 u2_358(.a(s_73_27), .b(s_73_26), .c(s_73_25), .d(s_73_24), .cin(t_1008), .o(t_1027), .co(t_1028), .cout(t_1029));
compressor_4_2 u2_359(.a(s_74_3), .b(s_74_2), .c(s_74_1), .d(s_74_0), .cin(t_1011), .o(t_1030), .co(t_1031), .cout(t_1032));
compressor_4_2 u2_360(.a(s_74_7), .b(s_74_6), .c(s_74_5), .d(s_74_4), .cin(t_1014), .o(t_1033), .co(t_1034), .cout(t_1035));
compressor_4_2 u2_361(.a(s_74_11), .b(s_74_10), .c(s_74_9), .d(s_74_8), .cin(t_1017), .o(t_1036), .co(t_1037), .cout(t_1038));
compressor_4_2 u2_362(.a(s_74_15), .b(s_74_14), .c(s_74_13), .d(s_74_12), .cin(t_1020), .o(t_1039), .co(t_1040), .cout(t_1041));
compressor_4_2 u2_363(.a(s_74_19), .b(s_74_18), .c(s_74_17), .d(s_74_16), .cin(t_1023), .o(t_1042), .co(t_1043), .cout(t_1044));
compressor_4_2 u2_364(.a(s_74_23), .b(s_74_22), .c(s_74_21), .d(s_74_20), .cin(t_1026), .o(t_1045), .co(t_1046), .cout(t_1047));
compressor_4_2 u2_365(.a(s_74_27), .b(s_74_26), .c(s_74_25), .d(s_74_24), .cin(t_1029), .o(t_1048), .co(t_1049), .cout(t_1050));
compressor_4_2 u2_366(.a(s_75_3), .b(s_75_2), .c(s_75_1), .d(s_75_0), .cin(t_1032), .o(t_1051), .co(t_1052), .cout(t_1053));
compressor_4_2 u2_367(.a(s_75_7), .b(s_75_6), .c(s_75_5), .d(s_75_4), .cin(t_1035), .o(t_1054), .co(t_1055), .cout(t_1056));
compressor_4_2 u2_368(.a(s_75_11), .b(s_75_10), .c(s_75_9), .d(s_75_8), .cin(t_1038), .o(t_1057), .co(t_1058), .cout(t_1059));
compressor_4_2 u2_369(.a(s_75_15), .b(s_75_14), .c(s_75_13), .d(s_75_12), .cin(t_1041), .o(t_1060), .co(t_1061), .cout(t_1062));
compressor_4_2 u2_370(.a(s_75_19), .b(s_75_18), .c(s_75_17), .d(s_75_16), .cin(t_1044), .o(t_1063), .co(t_1064), .cout(t_1065));
compressor_4_2 u2_371(.a(s_75_23), .b(s_75_22), .c(s_75_21), .d(s_75_20), .cin(t_1047), .o(t_1066), .co(t_1067), .cout(t_1068));
compressor_4_2 u2_372(.a(s_75_27), .b(s_75_26), .c(s_75_25), .d(s_75_24), .cin(t_1050), .o(t_1069), .co(t_1070), .cout(t_1071));
compressor_4_2 u2_373(.a(s_76_3), .b(s_76_2), .c(s_76_1), .d(s_76_0), .cin(t_1053), .o(t_1072), .co(t_1073), .cout(t_1074));
compressor_4_2 u2_374(.a(s_76_7), .b(s_76_6), .c(s_76_5), .d(s_76_4), .cin(t_1056), .o(t_1075), .co(t_1076), .cout(t_1077));
compressor_4_2 u2_375(.a(s_76_11), .b(s_76_10), .c(s_76_9), .d(s_76_8), .cin(t_1059), .o(t_1078), .co(t_1079), .cout(t_1080));
compressor_4_2 u2_376(.a(s_76_15), .b(s_76_14), .c(s_76_13), .d(s_76_12), .cin(t_1062), .o(t_1081), .co(t_1082), .cout(t_1083));
compressor_4_2 u2_377(.a(s_76_19), .b(s_76_18), .c(s_76_17), .d(s_76_16), .cin(t_1065), .o(t_1084), .co(t_1085), .cout(t_1086));
compressor_4_2 u2_378(.a(s_76_23), .b(s_76_22), .c(s_76_21), .d(s_76_20), .cin(t_1068), .o(t_1087), .co(t_1088), .cout(t_1089));
compressor_3_2 u1_379(.a(s_76_25), .b(s_76_24), .cin(t_1071), .o(t_1090), .cout(t_1091));
compressor_4_2 u2_380(.a(s_77_3), .b(s_77_2), .c(s_77_1), .d(s_77_0), .cin(t_1074), .o(t_1092), .co(t_1093), .cout(t_1094));
compressor_4_2 u2_381(.a(s_77_7), .b(s_77_6), .c(s_77_5), .d(s_77_4), .cin(t_1077), .o(t_1095), .co(t_1096), .cout(t_1097));
compressor_4_2 u2_382(.a(s_77_11), .b(s_77_10), .c(s_77_9), .d(s_77_8), .cin(t_1080), .o(t_1098), .co(t_1099), .cout(t_1100));
compressor_4_2 u2_383(.a(s_77_15), .b(s_77_14), .c(s_77_13), .d(s_77_12), .cin(t_1083), .o(t_1101), .co(t_1102), .cout(t_1103));
compressor_4_2 u2_384(.a(s_77_19), .b(s_77_18), .c(s_77_17), .d(s_77_16), .cin(t_1086), .o(t_1104), .co(t_1105), .cout(t_1106));
compressor_4_2 u2_385(.a(s_77_23), .b(s_77_22), .c(s_77_21), .d(s_77_20), .cin(t_1089), .o(t_1107), .co(t_1108), .cout(t_1109));
compressor_3_2 u1_386(.a(s_77_26), .b(s_77_25), .cin(s_77_24), .o(t_1110), .cout(t_1111));
compressor_4_2 u2_387(.a(s_78_3), .b(s_78_2), .c(s_78_1), .d(s_78_0), .cin(t_1094), .o(t_1112), .co(t_1113), .cout(t_1114));
compressor_4_2 u2_388(.a(s_78_7), .b(s_78_6), .c(s_78_5), .d(s_78_4), .cin(t_1097), .o(t_1115), .co(t_1116), .cout(t_1117));
compressor_4_2 u2_389(.a(s_78_11), .b(s_78_10), .c(s_78_9), .d(s_78_8), .cin(t_1100), .o(t_1118), .co(t_1119), .cout(t_1120));
compressor_4_2 u2_390(.a(s_78_15), .b(s_78_14), .c(s_78_13), .d(s_78_12), .cin(t_1103), .o(t_1121), .co(t_1122), .cout(t_1123));
compressor_4_2 u2_391(.a(s_78_19), .b(s_78_18), .c(s_78_17), .d(s_78_16), .cin(t_1106), .o(t_1124), .co(t_1125), .cout(t_1126));
compressor_4_2 u2_392(.a(s_78_23), .b(s_78_22), .c(s_78_21), .d(s_78_20), .cin(t_1109), .o(t_1127), .co(t_1128), .cout(t_1129));
half_adder u0_393(.a(s_78_25), .b(s_78_24), .o(t_1130), .cout(t_1131));
compressor_4_2 u2_394(.a(s_79_3), .b(s_79_2), .c(s_79_1), .d(s_79_0), .cin(t_1114), .o(t_1132), .co(t_1133), .cout(t_1134));
compressor_4_2 u2_395(.a(s_79_7), .b(s_79_6), .c(s_79_5), .d(s_79_4), .cin(t_1117), .o(t_1135), .co(t_1136), .cout(t_1137));
compressor_4_2 u2_396(.a(s_79_11), .b(s_79_10), .c(s_79_9), .d(s_79_8), .cin(t_1120), .o(t_1138), .co(t_1139), .cout(t_1140));
compressor_4_2 u2_397(.a(s_79_15), .b(s_79_14), .c(s_79_13), .d(s_79_12), .cin(t_1123), .o(t_1141), .co(t_1142), .cout(t_1143));
compressor_4_2 u2_398(.a(s_79_19), .b(s_79_18), .c(s_79_17), .d(s_79_16), .cin(t_1126), .o(t_1144), .co(t_1145), .cout(t_1146));
compressor_4_2 u2_399(.a(s_79_23), .b(s_79_22), .c(s_79_21), .d(s_79_20), .cin(t_1129), .o(t_1147), .co(t_1148), .cout(t_1149));
half_adder u0_400(.a(s_79_25), .b(s_79_24), .o(t_1150), .cout(t_1151));
compressor_4_2 u2_401(.a(s_80_3), .b(s_80_2), .c(s_80_1), .d(s_80_0), .cin(t_1134), .o(t_1152), .co(t_1153), .cout(t_1154));
compressor_4_2 u2_402(.a(s_80_7), .b(s_80_6), .c(s_80_5), .d(s_80_4), .cin(t_1137), .o(t_1155), .co(t_1156), .cout(t_1157));
compressor_4_2 u2_403(.a(s_80_11), .b(s_80_10), .c(s_80_9), .d(s_80_8), .cin(t_1140), .o(t_1158), .co(t_1159), .cout(t_1160));
compressor_4_2 u2_404(.a(s_80_15), .b(s_80_14), .c(s_80_13), .d(s_80_12), .cin(t_1143), .o(t_1161), .co(t_1162), .cout(t_1163));
compressor_4_2 u2_405(.a(s_80_19), .b(s_80_18), .c(s_80_17), .d(s_80_16), .cin(t_1146), .o(t_1164), .co(t_1165), .cout(t_1166));
compressor_4_2 u2_406(.a(s_80_23), .b(s_80_22), .c(s_80_21), .d(s_80_20), .cin(t_1149), .o(t_1167), .co(t_1168), .cout(t_1169));
compressor_4_2 u2_407(.a(s_81_3), .b(s_81_2), .c(s_81_1), .d(s_81_0), .cin(t_1154), .o(t_1170), .co(t_1171), .cout(t_1172));
compressor_4_2 u2_408(.a(s_81_7), .b(s_81_6), .c(s_81_5), .d(s_81_4), .cin(t_1157), .o(t_1173), .co(t_1174), .cout(t_1175));
compressor_4_2 u2_409(.a(s_81_11), .b(s_81_10), .c(s_81_9), .d(s_81_8), .cin(t_1160), .o(t_1176), .co(t_1177), .cout(t_1178));
compressor_4_2 u2_410(.a(s_81_15), .b(s_81_14), .c(s_81_13), .d(s_81_12), .cin(t_1163), .o(t_1179), .co(t_1180), .cout(t_1181));
compressor_4_2 u2_411(.a(s_81_19), .b(s_81_18), .c(s_81_17), .d(s_81_16), .cin(t_1166), .o(t_1182), .co(t_1183), .cout(t_1184));
compressor_4_2 u2_412(.a(s_81_23), .b(s_81_22), .c(s_81_21), .d(s_81_20), .cin(t_1169), .o(t_1185), .co(t_1186), .cout(t_1187));
compressor_4_2 u2_413(.a(s_82_3), .b(s_82_2), .c(s_82_1), .d(s_82_0), .cin(t_1172), .o(t_1188), .co(t_1189), .cout(t_1190));
compressor_4_2 u2_414(.a(s_82_7), .b(s_82_6), .c(s_82_5), .d(s_82_4), .cin(t_1175), .o(t_1191), .co(t_1192), .cout(t_1193));
compressor_4_2 u2_415(.a(s_82_11), .b(s_82_10), .c(s_82_9), .d(s_82_8), .cin(t_1178), .o(t_1194), .co(t_1195), .cout(t_1196));
compressor_4_2 u2_416(.a(s_82_15), .b(s_82_14), .c(s_82_13), .d(s_82_12), .cin(t_1181), .o(t_1197), .co(t_1198), .cout(t_1199));
compressor_4_2 u2_417(.a(s_82_19), .b(s_82_18), .c(s_82_17), .d(s_82_16), .cin(t_1184), .o(t_1200), .co(t_1201), .cout(t_1202));
compressor_4_2 u2_418(.a(s_82_23), .b(s_82_22), .c(s_82_21), .d(s_82_20), .cin(t_1187), .o(t_1203), .co(t_1204), .cout(t_1205));
compressor_4_2 u2_419(.a(s_83_3), .b(s_83_2), .c(s_83_1), .d(s_83_0), .cin(t_1190), .o(t_1206), .co(t_1207), .cout(t_1208));
compressor_4_2 u2_420(.a(s_83_7), .b(s_83_6), .c(s_83_5), .d(s_83_4), .cin(t_1193), .o(t_1209), .co(t_1210), .cout(t_1211));
compressor_4_2 u2_421(.a(s_83_11), .b(s_83_10), .c(s_83_9), .d(s_83_8), .cin(t_1196), .o(t_1212), .co(t_1213), .cout(t_1214));
compressor_4_2 u2_422(.a(s_83_15), .b(s_83_14), .c(s_83_13), .d(s_83_12), .cin(t_1199), .o(t_1215), .co(t_1216), .cout(t_1217));
compressor_4_2 u2_423(.a(s_83_19), .b(s_83_18), .c(s_83_17), .d(s_83_16), .cin(t_1202), .o(t_1218), .co(t_1219), .cout(t_1220));
compressor_4_2 u2_424(.a(s_83_23), .b(s_83_22), .c(s_83_21), .d(s_83_20), .cin(t_1205), .o(t_1221), .co(t_1222), .cout(t_1223));
compressor_4_2 u2_425(.a(s_84_3), .b(s_84_2), .c(s_84_1), .d(s_84_0), .cin(t_1208), .o(t_1224), .co(t_1225), .cout(t_1226));
compressor_4_2 u2_426(.a(s_84_7), .b(s_84_6), .c(s_84_5), .d(s_84_4), .cin(t_1211), .o(t_1227), .co(t_1228), .cout(t_1229));
compressor_4_2 u2_427(.a(s_84_11), .b(s_84_10), .c(s_84_9), .d(s_84_8), .cin(t_1214), .o(t_1230), .co(t_1231), .cout(t_1232));
compressor_4_2 u2_428(.a(s_84_15), .b(s_84_14), .c(s_84_13), .d(s_84_12), .cin(t_1217), .o(t_1233), .co(t_1234), .cout(t_1235));
compressor_4_2 u2_429(.a(s_84_19), .b(s_84_18), .c(s_84_17), .d(s_84_16), .cin(t_1220), .o(t_1236), .co(t_1237), .cout(t_1238));
compressor_3_2 u1_430(.a(s_84_21), .b(s_84_20), .cin(t_1223), .o(t_1239), .cout(t_1240));
compressor_4_2 u2_431(.a(s_85_3), .b(s_85_2), .c(s_85_1), .d(s_85_0), .cin(t_1226), .o(t_1241), .co(t_1242), .cout(t_1243));
compressor_4_2 u2_432(.a(s_85_7), .b(s_85_6), .c(s_85_5), .d(s_85_4), .cin(t_1229), .o(t_1244), .co(t_1245), .cout(t_1246));
compressor_4_2 u2_433(.a(s_85_11), .b(s_85_10), .c(s_85_9), .d(s_85_8), .cin(t_1232), .o(t_1247), .co(t_1248), .cout(t_1249));
compressor_4_2 u2_434(.a(s_85_15), .b(s_85_14), .c(s_85_13), .d(s_85_12), .cin(t_1235), .o(t_1250), .co(t_1251), .cout(t_1252));
compressor_4_2 u2_435(.a(s_85_19), .b(s_85_18), .c(s_85_17), .d(s_85_16), .cin(t_1238), .o(t_1253), .co(t_1254), .cout(t_1255));
compressor_3_2 u1_436(.a(s_85_22), .b(s_85_21), .cin(s_85_20), .o(t_1256), .cout(t_1257));
compressor_4_2 u2_437(.a(s_86_3), .b(s_86_2), .c(s_86_1), .d(s_86_0), .cin(t_1243), .o(t_1258), .co(t_1259), .cout(t_1260));
compressor_4_2 u2_438(.a(s_86_7), .b(s_86_6), .c(s_86_5), .d(s_86_4), .cin(t_1246), .o(t_1261), .co(t_1262), .cout(t_1263));
compressor_4_2 u2_439(.a(s_86_11), .b(s_86_10), .c(s_86_9), .d(s_86_8), .cin(t_1249), .o(t_1264), .co(t_1265), .cout(t_1266));
compressor_4_2 u2_440(.a(s_86_15), .b(s_86_14), .c(s_86_13), .d(s_86_12), .cin(t_1252), .o(t_1267), .co(t_1268), .cout(t_1269));
compressor_4_2 u2_441(.a(s_86_19), .b(s_86_18), .c(s_86_17), .d(s_86_16), .cin(t_1255), .o(t_1270), .co(t_1271), .cout(t_1272));
half_adder u0_442(.a(s_86_21), .b(s_86_20), .o(t_1273), .cout(t_1274));
compressor_4_2 u2_443(.a(s_87_3), .b(s_87_2), .c(s_87_1), .d(s_87_0), .cin(t_1260), .o(t_1275), .co(t_1276), .cout(t_1277));
compressor_4_2 u2_444(.a(s_87_7), .b(s_87_6), .c(s_87_5), .d(s_87_4), .cin(t_1263), .o(t_1278), .co(t_1279), .cout(t_1280));
compressor_4_2 u2_445(.a(s_87_11), .b(s_87_10), .c(s_87_9), .d(s_87_8), .cin(t_1266), .o(t_1281), .co(t_1282), .cout(t_1283));
compressor_4_2 u2_446(.a(s_87_15), .b(s_87_14), .c(s_87_13), .d(s_87_12), .cin(t_1269), .o(t_1284), .co(t_1285), .cout(t_1286));
compressor_4_2 u2_447(.a(s_87_19), .b(s_87_18), .c(s_87_17), .d(s_87_16), .cin(t_1272), .o(t_1287), .co(t_1288), .cout(t_1289));
half_adder u0_448(.a(s_87_21), .b(s_87_20), .o(t_1290), .cout(t_1291));
compressor_4_2 u2_449(.a(s_88_3), .b(s_88_2), .c(s_88_1), .d(s_88_0), .cin(t_1277), .o(t_1292), .co(t_1293), .cout(t_1294));
compressor_4_2 u2_450(.a(s_88_7), .b(s_88_6), .c(s_88_5), .d(s_88_4), .cin(t_1280), .o(t_1295), .co(t_1296), .cout(t_1297));
compressor_4_2 u2_451(.a(s_88_11), .b(s_88_10), .c(s_88_9), .d(s_88_8), .cin(t_1283), .o(t_1298), .co(t_1299), .cout(t_1300));
compressor_4_2 u2_452(.a(s_88_15), .b(s_88_14), .c(s_88_13), .d(s_88_12), .cin(t_1286), .o(t_1301), .co(t_1302), .cout(t_1303));
compressor_4_2 u2_453(.a(s_88_19), .b(s_88_18), .c(s_88_17), .d(s_88_16), .cin(t_1289), .o(t_1304), .co(t_1305), .cout(t_1306));
compressor_4_2 u2_454(.a(s_89_3), .b(s_89_2), .c(s_89_1), .d(s_89_0), .cin(t_1294), .o(t_1307), .co(t_1308), .cout(t_1309));
compressor_4_2 u2_455(.a(s_89_7), .b(s_89_6), .c(s_89_5), .d(s_89_4), .cin(t_1297), .o(t_1310), .co(t_1311), .cout(t_1312));
compressor_4_2 u2_456(.a(s_89_11), .b(s_89_10), .c(s_89_9), .d(s_89_8), .cin(t_1300), .o(t_1313), .co(t_1314), .cout(t_1315));
compressor_4_2 u2_457(.a(s_89_15), .b(s_89_14), .c(s_89_13), .d(s_89_12), .cin(t_1303), .o(t_1316), .co(t_1317), .cout(t_1318));
compressor_4_2 u2_458(.a(s_89_19), .b(s_89_18), .c(s_89_17), .d(s_89_16), .cin(t_1306), .o(t_1319), .co(t_1320), .cout(t_1321));
compressor_4_2 u2_459(.a(s_90_3), .b(s_90_2), .c(s_90_1), .d(s_90_0), .cin(t_1309), .o(t_1322), .co(t_1323), .cout(t_1324));
compressor_4_2 u2_460(.a(s_90_7), .b(s_90_6), .c(s_90_5), .d(s_90_4), .cin(t_1312), .o(t_1325), .co(t_1326), .cout(t_1327));
compressor_4_2 u2_461(.a(s_90_11), .b(s_90_10), .c(s_90_9), .d(s_90_8), .cin(t_1315), .o(t_1328), .co(t_1329), .cout(t_1330));
compressor_4_2 u2_462(.a(s_90_15), .b(s_90_14), .c(s_90_13), .d(s_90_12), .cin(t_1318), .o(t_1331), .co(t_1332), .cout(t_1333));
compressor_4_2 u2_463(.a(s_90_19), .b(s_90_18), .c(s_90_17), .d(s_90_16), .cin(t_1321), .o(t_1334), .co(t_1335), .cout(t_1336));
compressor_4_2 u2_464(.a(s_91_3), .b(s_91_2), .c(s_91_1), .d(s_91_0), .cin(t_1324), .o(t_1337), .co(t_1338), .cout(t_1339));
compressor_4_2 u2_465(.a(s_91_7), .b(s_91_6), .c(s_91_5), .d(s_91_4), .cin(t_1327), .o(t_1340), .co(t_1341), .cout(t_1342));
compressor_4_2 u2_466(.a(s_91_11), .b(s_91_10), .c(s_91_9), .d(s_91_8), .cin(t_1330), .o(t_1343), .co(t_1344), .cout(t_1345));
compressor_4_2 u2_467(.a(s_91_15), .b(s_91_14), .c(s_91_13), .d(s_91_12), .cin(t_1333), .o(t_1346), .co(t_1347), .cout(t_1348));
compressor_4_2 u2_468(.a(s_91_19), .b(s_91_18), .c(s_91_17), .d(s_91_16), .cin(t_1336), .o(t_1349), .co(t_1350), .cout(t_1351));
compressor_4_2 u2_469(.a(s_92_3), .b(s_92_2), .c(s_92_1), .d(s_92_0), .cin(t_1339), .o(t_1352), .co(t_1353), .cout(t_1354));
compressor_4_2 u2_470(.a(s_92_7), .b(s_92_6), .c(s_92_5), .d(s_92_4), .cin(t_1342), .o(t_1355), .co(t_1356), .cout(t_1357));
compressor_4_2 u2_471(.a(s_92_11), .b(s_92_10), .c(s_92_9), .d(s_92_8), .cin(t_1345), .o(t_1358), .co(t_1359), .cout(t_1360));
compressor_4_2 u2_472(.a(s_92_15), .b(s_92_14), .c(s_92_13), .d(s_92_12), .cin(t_1348), .o(t_1361), .co(t_1362), .cout(t_1363));
compressor_3_2 u1_473(.a(s_92_17), .b(s_92_16), .cin(t_1351), .o(t_1364), .cout(t_1365));
compressor_4_2 u2_474(.a(s_93_3), .b(s_93_2), .c(s_93_1), .d(s_93_0), .cin(t_1354), .o(t_1366), .co(t_1367), .cout(t_1368));
compressor_4_2 u2_475(.a(s_93_7), .b(s_93_6), .c(s_93_5), .d(s_93_4), .cin(t_1357), .o(t_1369), .co(t_1370), .cout(t_1371));
compressor_4_2 u2_476(.a(s_93_11), .b(s_93_10), .c(s_93_9), .d(s_93_8), .cin(t_1360), .o(t_1372), .co(t_1373), .cout(t_1374));
compressor_4_2 u2_477(.a(s_93_15), .b(s_93_14), .c(s_93_13), .d(s_93_12), .cin(t_1363), .o(t_1375), .co(t_1376), .cout(t_1377));
compressor_3_2 u1_478(.a(s_93_18), .b(s_93_17), .cin(s_93_16), .o(t_1378), .cout(t_1379));
compressor_4_2 u2_479(.a(s_94_3), .b(s_94_2), .c(s_94_1), .d(s_94_0), .cin(t_1368), .o(t_1380), .co(t_1381), .cout(t_1382));
compressor_4_2 u2_480(.a(s_94_7), .b(s_94_6), .c(s_94_5), .d(s_94_4), .cin(t_1371), .o(t_1383), .co(t_1384), .cout(t_1385));
compressor_4_2 u2_481(.a(s_94_11), .b(s_94_10), .c(s_94_9), .d(s_94_8), .cin(t_1374), .o(t_1386), .co(t_1387), .cout(t_1388));
compressor_4_2 u2_482(.a(s_94_15), .b(s_94_14), .c(s_94_13), .d(s_94_12), .cin(t_1377), .o(t_1389), .co(t_1390), .cout(t_1391));
half_adder u0_483(.a(s_94_17), .b(s_94_16), .o(t_1392), .cout(t_1393));
compressor_4_2 u2_484(.a(s_95_3), .b(s_95_2), .c(s_95_1), .d(s_95_0), .cin(t_1382), .o(t_1394), .co(t_1395), .cout(t_1396));
compressor_4_2 u2_485(.a(s_95_7), .b(s_95_6), .c(s_95_5), .d(s_95_4), .cin(t_1385), .o(t_1397), .co(t_1398), .cout(t_1399));
compressor_4_2 u2_486(.a(s_95_11), .b(s_95_10), .c(s_95_9), .d(s_95_8), .cin(t_1388), .o(t_1400), .co(t_1401), .cout(t_1402));
compressor_4_2 u2_487(.a(s_95_15), .b(s_95_14), .c(s_95_13), .d(s_95_12), .cin(t_1391), .o(t_1403), .co(t_1404), .cout(t_1405));
half_adder u0_488(.a(s_95_17), .b(s_95_16), .o(t_1406), .cout(t_1407));
compressor_4_2 u2_489(.a(s_96_3), .b(s_96_2), .c(s_96_1), .d(s_96_0), .cin(t_1396), .o(t_1408), .co(t_1409), .cout(t_1410));
compressor_4_2 u2_490(.a(s_96_7), .b(s_96_6), .c(s_96_5), .d(s_96_4), .cin(t_1399), .o(t_1411), .co(t_1412), .cout(t_1413));
compressor_4_2 u2_491(.a(s_96_11), .b(s_96_10), .c(s_96_9), .d(s_96_8), .cin(t_1402), .o(t_1414), .co(t_1415), .cout(t_1416));
compressor_4_2 u2_492(.a(s_96_15), .b(s_96_14), .c(s_96_13), .d(s_96_12), .cin(t_1405), .o(t_1417), .co(t_1418), .cout(t_1419));
compressor_4_2 u2_493(.a(s_97_3), .b(s_97_2), .c(s_97_1), .d(s_97_0), .cin(t_1410), .o(t_1420), .co(t_1421), .cout(t_1422));
compressor_4_2 u2_494(.a(s_97_7), .b(s_97_6), .c(s_97_5), .d(s_97_4), .cin(t_1413), .o(t_1423), .co(t_1424), .cout(t_1425));
compressor_4_2 u2_495(.a(s_97_11), .b(s_97_10), .c(s_97_9), .d(s_97_8), .cin(t_1416), .o(t_1426), .co(t_1427), .cout(t_1428));
compressor_4_2 u2_496(.a(s_97_15), .b(s_97_14), .c(s_97_13), .d(s_97_12), .cin(t_1419), .o(t_1429), .co(t_1430), .cout(t_1431));
compressor_4_2 u2_497(.a(s_98_3), .b(s_98_2), .c(s_98_1), .d(s_98_0), .cin(t_1422), .o(t_1432), .co(t_1433), .cout(t_1434));
compressor_4_2 u2_498(.a(s_98_7), .b(s_98_6), .c(s_98_5), .d(s_98_4), .cin(t_1425), .o(t_1435), .co(t_1436), .cout(t_1437));
compressor_4_2 u2_499(.a(s_98_11), .b(s_98_10), .c(s_98_9), .d(s_98_8), .cin(t_1428), .o(t_1438), .co(t_1439), .cout(t_1440));
compressor_4_2 u2_500(.a(s_98_15), .b(s_98_14), .c(s_98_13), .d(s_98_12), .cin(t_1431), .o(t_1441), .co(t_1442), .cout(t_1443));
compressor_4_2 u2_501(.a(s_99_3), .b(s_99_2), .c(s_99_1), .d(s_99_0), .cin(t_1434), .o(t_1444), .co(t_1445), .cout(t_1446));
compressor_4_2 u2_502(.a(s_99_7), .b(s_99_6), .c(s_99_5), .d(s_99_4), .cin(t_1437), .o(t_1447), .co(t_1448), .cout(t_1449));
compressor_4_2 u2_503(.a(s_99_11), .b(s_99_10), .c(s_99_9), .d(s_99_8), .cin(t_1440), .o(t_1450), .co(t_1451), .cout(t_1452));
compressor_4_2 u2_504(.a(s_99_15), .b(s_99_14), .c(s_99_13), .d(s_99_12), .cin(t_1443), .o(t_1453), .co(t_1454), .cout(t_1455));
compressor_4_2 u2_505(.a(s_100_3), .b(s_100_2), .c(s_100_1), .d(s_100_0), .cin(t_1446), .o(t_1456), .co(t_1457), .cout(t_1458));
compressor_4_2 u2_506(.a(s_100_7), .b(s_100_6), .c(s_100_5), .d(s_100_4), .cin(t_1449), .o(t_1459), .co(t_1460), .cout(t_1461));
compressor_4_2 u2_507(.a(s_100_11), .b(s_100_10), .c(s_100_9), .d(s_100_8), .cin(t_1452), .o(t_1462), .co(t_1463), .cout(t_1464));
compressor_3_2 u1_508(.a(s_100_13), .b(s_100_12), .cin(t_1455), .o(t_1465), .cout(t_1466));
compressor_4_2 u2_509(.a(s_101_3), .b(s_101_2), .c(s_101_1), .d(s_101_0), .cin(t_1458), .o(t_1467), .co(t_1468), .cout(t_1469));
compressor_4_2 u2_510(.a(s_101_7), .b(s_101_6), .c(s_101_5), .d(s_101_4), .cin(t_1461), .o(t_1470), .co(t_1471), .cout(t_1472));
compressor_4_2 u2_511(.a(s_101_11), .b(s_101_10), .c(s_101_9), .d(s_101_8), .cin(t_1464), .o(t_1473), .co(t_1474), .cout(t_1475));
compressor_3_2 u1_512(.a(s_101_14), .b(s_101_13), .cin(s_101_12), .o(t_1476), .cout(t_1477));
compressor_4_2 u2_513(.a(s_102_3), .b(s_102_2), .c(s_102_1), .d(s_102_0), .cin(t_1469), .o(t_1478), .co(t_1479), .cout(t_1480));
compressor_4_2 u2_514(.a(s_102_7), .b(s_102_6), .c(s_102_5), .d(s_102_4), .cin(t_1472), .o(t_1481), .co(t_1482), .cout(t_1483));
compressor_4_2 u2_515(.a(s_102_11), .b(s_102_10), .c(s_102_9), .d(s_102_8), .cin(t_1475), .o(t_1484), .co(t_1485), .cout(t_1486));
half_adder u0_516(.a(s_102_13), .b(s_102_12), .o(t_1487), .cout(t_1488));
compressor_4_2 u2_517(.a(s_103_3), .b(s_103_2), .c(s_103_1), .d(s_103_0), .cin(t_1480), .o(t_1489), .co(t_1490), .cout(t_1491));
compressor_4_2 u2_518(.a(s_103_7), .b(s_103_6), .c(s_103_5), .d(s_103_4), .cin(t_1483), .o(t_1492), .co(t_1493), .cout(t_1494));
compressor_4_2 u2_519(.a(s_103_11), .b(s_103_10), .c(s_103_9), .d(s_103_8), .cin(t_1486), .o(t_1495), .co(t_1496), .cout(t_1497));
half_adder u0_520(.a(s_103_13), .b(s_103_12), .o(t_1498), .cout(t_1499));
compressor_4_2 u2_521(.a(s_104_3), .b(s_104_2), .c(s_104_1), .d(s_104_0), .cin(t_1491), .o(t_1500), .co(t_1501), .cout(t_1502));
compressor_4_2 u2_522(.a(s_104_7), .b(s_104_6), .c(s_104_5), .d(s_104_4), .cin(t_1494), .o(t_1503), .co(t_1504), .cout(t_1505));
compressor_4_2 u2_523(.a(s_104_11), .b(s_104_10), .c(s_104_9), .d(s_104_8), .cin(t_1497), .o(t_1506), .co(t_1507), .cout(t_1508));
compressor_4_2 u2_524(.a(s_105_3), .b(s_105_2), .c(s_105_1), .d(s_105_0), .cin(t_1502), .o(t_1509), .co(t_1510), .cout(t_1511));
compressor_4_2 u2_525(.a(s_105_7), .b(s_105_6), .c(s_105_5), .d(s_105_4), .cin(t_1505), .o(t_1512), .co(t_1513), .cout(t_1514));
compressor_4_2 u2_526(.a(s_105_11), .b(s_105_10), .c(s_105_9), .d(s_105_8), .cin(t_1508), .o(t_1515), .co(t_1516), .cout(t_1517));
compressor_4_2 u2_527(.a(s_106_3), .b(s_106_2), .c(s_106_1), .d(s_106_0), .cin(t_1511), .o(t_1518), .co(t_1519), .cout(t_1520));
compressor_4_2 u2_528(.a(s_106_7), .b(s_106_6), .c(s_106_5), .d(s_106_4), .cin(t_1514), .o(t_1521), .co(t_1522), .cout(t_1523));
compressor_4_2 u2_529(.a(s_106_11), .b(s_106_10), .c(s_106_9), .d(s_106_8), .cin(t_1517), .o(t_1524), .co(t_1525), .cout(t_1526));
compressor_4_2 u2_530(.a(s_107_3), .b(s_107_2), .c(s_107_1), .d(s_107_0), .cin(t_1520), .o(t_1527), .co(t_1528), .cout(t_1529));
compressor_4_2 u2_531(.a(s_107_7), .b(s_107_6), .c(s_107_5), .d(s_107_4), .cin(t_1523), .o(t_1530), .co(t_1531), .cout(t_1532));
compressor_4_2 u2_532(.a(s_107_11), .b(s_107_10), .c(s_107_9), .d(s_107_8), .cin(t_1526), .o(t_1533), .co(t_1534), .cout(t_1535));
compressor_4_2 u2_533(.a(s_108_3), .b(s_108_2), .c(s_108_1), .d(s_108_0), .cin(t_1529), .o(t_1536), .co(t_1537), .cout(t_1538));
compressor_4_2 u2_534(.a(s_108_7), .b(s_108_6), .c(s_108_5), .d(s_108_4), .cin(t_1532), .o(t_1539), .co(t_1540), .cout(t_1541));
compressor_3_2 u1_535(.a(s_108_9), .b(s_108_8), .cin(t_1535), .o(t_1542), .cout(t_1543));
compressor_4_2 u2_536(.a(s_109_3), .b(s_109_2), .c(s_109_1), .d(s_109_0), .cin(t_1538), .o(t_1544), .co(t_1545), .cout(t_1546));
compressor_4_2 u2_537(.a(s_109_7), .b(s_109_6), .c(s_109_5), .d(s_109_4), .cin(t_1541), .o(t_1547), .co(t_1548), .cout(t_1549));
compressor_3_2 u1_538(.a(s_109_10), .b(s_109_9), .cin(s_109_8), .o(t_1550), .cout(t_1551));
compressor_4_2 u2_539(.a(s_110_3), .b(s_110_2), .c(s_110_1), .d(s_110_0), .cin(t_1546), .o(t_1552), .co(t_1553), .cout(t_1554));
compressor_4_2 u2_540(.a(s_110_7), .b(s_110_6), .c(s_110_5), .d(s_110_4), .cin(t_1549), .o(t_1555), .co(t_1556), .cout(t_1557));
half_adder u0_541(.a(s_110_9), .b(s_110_8), .o(t_1558), .cout(t_1559));
compressor_4_2 u2_542(.a(s_111_3), .b(s_111_2), .c(s_111_1), .d(s_111_0), .cin(t_1554), .o(t_1560), .co(t_1561), .cout(t_1562));
compressor_4_2 u2_543(.a(s_111_7), .b(s_111_6), .c(s_111_5), .d(s_111_4), .cin(t_1557), .o(t_1563), .co(t_1564), .cout(t_1565));
half_adder u0_544(.a(s_111_9), .b(s_111_8), .o(t_1566), .cout(t_1567));
compressor_4_2 u2_545(.a(s_112_3), .b(s_112_2), .c(s_112_1), .d(s_112_0), .cin(t_1562), .o(t_1568), .co(t_1569), .cout(t_1570));
compressor_4_2 u2_546(.a(s_112_7), .b(s_112_6), .c(s_112_5), .d(s_112_4), .cin(t_1565), .o(t_1571), .co(t_1572), .cout(t_1573));
compressor_4_2 u2_547(.a(s_113_3), .b(s_113_2), .c(s_113_1), .d(s_113_0), .cin(t_1570), .o(t_1574), .co(t_1575), .cout(t_1576));
compressor_4_2 u2_548(.a(s_113_7), .b(s_113_6), .c(s_113_5), .d(s_113_4), .cin(t_1573), .o(t_1577), .co(t_1578), .cout(t_1579));
compressor_4_2 u2_549(.a(s_114_3), .b(s_114_2), .c(s_114_1), .d(s_114_0), .cin(t_1576), .o(t_1580), .co(t_1581), .cout(t_1582));
compressor_4_2 u2_550(.a(s_114_7), .b(s_114_6), .c(s_114_5), .d(s_114_4), .cin(t_1579), .o(t_1583), .co(t_1584), .cout(t_1585));
compressor_4_2 u2_551(.a(s_115_3), .b(s_115_2), .c(s_115_1), .d(s_115_0), .cin(t_1582), .o(t_1586), .co(t_1587), .cout(t_1588));
compressor_4_2 u2_552(.a(s_115_7), .b(s_115_6), .c(s_115_5), .d(s_115_4), .cin(t_1585), .o(t_1589), .co(t_1590), .cout(t_1591));
compressor_4_2 u2_553(.a(s_116_3), .b(s_116_2), .c(s_116_1), .d(s_116_0), .cin(t_1588), .o(t_1592), .co(t_1593), .cout(t_1594));
compressor_3_2 u1_554(.a(s_116_5), .b(s_116_4), .cin(t_1591), .o(t_1595), .cout(t_1596));
compressor_4_2 u2_555(.a(s_117_3), .b(s_117_2), .c(s_117_1), .d(s_117_0), .cin(t_1594), .o(t_1597), .co(t_1598), .cout(t_1599));
compressor_3_2 u1_556(.a(s_117_6), .b(s_117_5), .cin(s_117_4), .o(t_1600), .cout(t_1601));
compressor_4_2 u2_557(.a(s_118_3), .b(s_118_2), .c(s_118_1), .d(s_118_0), .cin(t_1599), .o(t_1602), .co(t_1603), .cout(t_1604));
half_adder u0_558(.a(s_118_5), .b(s_118_4), .o(t_1605), .cout(t_1606));
compressor_4_2 u2_559(.a(s_119_3), .b(s_119_2), .c(s_119_1), .d(s_119_0), .cin(t_1604), .o(t_1607), .co(t_1608), .cout(t_1609));
half_adder u0_560(.a(s_119_5), .b(s_119_4), .o(t_1610), .cout(t_1611));
compressor_4_2 u2_561(.a(s_120_3), .b(s_120_2), .c(s_120_1), .d(s_120_0), .cin(t_1609), .o(t_1612), .co(t_1613), .cout(t_1614));
compressor_4_2 u2_562(.a(s_121_3), .b(s_121_2), .c(s_121_1), .d(s_121_0), .cin(t_1614), .o(t_1615), .co(t_1616), .cout(t_1617));
compressor_4_2 u2_563(.a(s_122_3), .b(s_122_2), .c(s_122_1), .d(s_122_0), .cin(t_1617), .o(t_1618), .co(t_1619), .cout(t_1620));
compressor_4_2 u2_564(.a(s_123_3), .b(s_123_2), .c(s_123_1), .d(s_123_0), .cin(t_1620), .o(t_1621), .co(t_1622), .cout(t_1623));
compressor_3_2 u1_565(.a(s_124_1), .b(s_124_0), .cin(t_1623), .o(t_1624), .cout(t_1625));
compressor_3_2 u1_566(.a(s_125_2), .b(s_125_1), .cin(s_125_0), .o(t_1626), .cout(t_1627));
half_adder u0_567(.a(s_126_1), .b(s_126_0), .o(t_1628), .cout(t_1629));
half_adder u0_568(.a(s_127_1), .b(s_127_0), .o(t_1630), .cout());

/* u0_569 Output nets */
wire t_1631,   t_1632;
/* u0_570 Output nets */
wire t_1633,   t_1634;
/* u1_571 Output nets */
wire t_1635,   t_1636;
/* u0_572 Output nets */
wire t_1637,   t_1638;
/* u0_573 Output nets */
wire t_1639,   t_1640;
/* u0_574 Output nets */
wire t_1641,   t_1642;
/* u1_575 Output nets */
wire t_1643,   t_1644;
/* u1_576 Output nets */
wire t_1645,   t_1646;
/* u1_577 Output nets */
wire t_1647,   t_1648;
/* u1_578 Output nets */
wire t_1649,   t_1650;
/* u2_579 Output nets */
wire t_1651,   t_1652,   t_1653;
/* u2_580 Output nets */
wire t_1654,   t_1655,   t_1656;
/* u2_581 Output nets */
wire t_1657,   t_1658,   t_1659;
/* u2_582 Output nets */
wire t_1660,   t_1661,   t_1662;
/* u2_583 Output nets */
wire t_1663,   t_1664,   t_1665;
/* u2_584 Output nets */
wire t_1666,   t_1667,   t_1668;
/* u0_585 Output nets */
wire t_1669,   t_1670;
/* u2_586 Output nets */
wire t_1671,   t_1672,   t_1673;
/* u2_587 Output nets */
wire t_1674,   t_1675,   t_1676;
/* u0_588 Output nets */
wire t_1677,   t_1678;
/* u2_589 Output nets */
wire t_1679,   t_1680,   t_1681;
/* u1_590 Output nets */
wire t_1682,   t_1683;
/* u2_591 Output nets */
wire t_1684,   t_1685,   t_1686;
/* u0_592 Output nets */
wire t_1687,   t_1688;
/* u2_593 Output nets */
wire t_1689,   t_1690,   t_1691;
/* u0_594 Output nets */
wire t_1692,   t_1693;
/* u2_595 Output nets */
wire t_1694,   t_1695,   t_1696;
/* u0_596 Output nets */
wire t_1697,   t_1698;
/* u2_597 Output nets */
wire t_1699,   t_1700,   t_1701;
/* u1_598 Output nets */
wire t_1702,   t_1703;
/* u2_599 Output nets */
wire t_1704,   t_1705,   t_1706;
/* u1_600 Output nets */
wire t_1707,   t_1708;
/* u2_601 Output nets */
wire t_1709,   t_1710,   t_1711;
/* u1_602 Output nets */
wire t_1712,   t_1713;
/* u2_603 Output nets */
wire t_1714,   t_1715,   t_1716;
/* u1_604 Output nets */
wire t_1717,   t_1718;
/* u2_605 Output nets */
wire t_1719,   t_1720,   t_1721;
/* u2_606 Output nets */
wire t_1722,   t_1723,   t_1724;
/* u2_607 Output nets */
wire t_1725,   t_1726,   t_1727;
/* u2_608 Output nets */
wire t_1728,   t_1729,   t_1730;
/* u2_609 Output nets */
wire t_1731,   t_1732,   t_1733;
/* u2_610 Output nets */
wire t_1734,   t_1735,   t_1736;
/* u2_611 Output nets */
wire t_1737,   t_1738,   t_1739;
/* u2_612 Output nets */
wire t_1740,   t_1741,   t_1742;
/* u2_613 Output nets */
wire t_1743,   t_1744,   t_1745;
/* u2_614 Output nets */
wire t_1746,   t_1747,   t_1748;
/* u2_615 Output nets */
wire t_1749,   t_1750,   t_1751;
/* u2_616 Output nets */
wire t_1752,   t_1753,   t_1754;
/* u0_617 Output nets */
wire t_1755,   t_1756;
/* u2_618 Output nets */
wire t_1757,   t_1758,   t_1759;
/* u2_619 Output nets */
wire t_1760,   t_1761,   t_1762;
/* u2_620 Output nets */
wire t_1763,   t_1764,   t_1765;
/* u2_621 Output nets */
wire t_1766,   t_1767,   t_1768;
/* u0_622 Output nets */
wire t_1769,   t_1770;
/* u2_623 Output nets */
wire t_1771,   t_1772,   t_1773;
/* u2_624 Output nets */
wire t_1774,   t_1775,   t_1776;
/* u1_625 Output nets */
wire t_1777,   t_1778;
/* u2_626 Output nets */
wire t_1779,   t_1780,   t_1781;
/* u2_627 Output nets */
wire t_1782,   t_1783,   t_1784;
/* u0_628 Output nets */
wire t_1785,   t_1786;
/* u2_629 Output nets */
wire t_1787,   t_1788,   t_1789;
/* u2_630 Output nets */
wire t_1790,   t_1791,   t_1792;
/* u0_631 Output nets */
wire t_1793,   t_1794;
/* u2_632 Output nets */
wire t_1795,   t_1796,   t_1797;
/* u2_633 Output nets */
wire t_1798,   t_1799,   t_1800;
/* u0_634 Output nets */
wire t_1801,   t_1802;
/* u2_635 Output nets */
wire t_1803,   t_1804,   t_1805;
/* u2_636 Output nets */
wire t_1806,   t_1807,   t_1808;
/* u1_637 Output nets */
wire t_1809,   t_1810;
/* u2_638 Output nets */
wire t_1811,   t_1812,   t_1813;
/* u2_639 Output nets */
wire t_1814,   t_1815,   t_1816;
/* u1_640 Output nets */
wire t_1817,   t_1818;
/* u2_641 Output nets */
wire t_1819,   t_1820,   t_1821;
/* u2_642 Output nets */
wire t_1822,   t_1823,   t_1824;
/* u1_643 Output nets */
wire t_1825,   t_1826;
/* u2_644 Output nets */
wire t_1827,   t_1828,   t_1829;
/* u2_645 Output nets */
wire t_1830,   t_1831,   t_1832;
/* u1_646 Output nets */
wire t_1833,   t_1834;
/* u2_647 Output nets */
wire t_1835,   t_1836,   t_1837;
/* u2_648 Output nets */
wire t_1838,   t_1839,   t_1840;
/* u2_649 Output nets */
wire t_1841,   t_1842,   t_1843;
/* u2_650 Output nets */
wire t_1844,   t_1845,   t_1846;
/* u2_651 Output nets */
wire t_1847,   t_1848,   t_1849;
/* u2_652 Output nets */
wire t_1850,   t_1851,   t_1852;
/* u2_653 Output nets */
wire t_1853,   t_1854,   t_1855;
/* u2_654 Output nets */
wire t_1856,   t_1857,   t_1858;
/* u2_655 Output nets */
wire t_1859,   t_1860,   t_1861;
/* u2_656 Output nets */
wire t_1862,   t_1863,   t_1864;
/* u2_657 Output nets */
wire t_1865,   t_1866,   t_1867;
/* u2_658 Output nets */
wire t_1868,   t_1869,   t_1870;
/* u2_659 Output nets */
wire t_1871,   t_1872,   t_1873;
/* u2_660 Output nets */
wire t_1874,   t_1875,   t_1876;
/* u2_661 Output nets */
wire t_1877,   t_1878,   t_1879;
/* u2_662 Output nets */
wire t_1880,   t_1881,   t_1882;
/* u2_663 Output nets */
wire t_1883,   t_1884,   t_1885;
/* u2_664 Output nets */
wire t_1886,   t_1887,   t_1888;
/* u0_665 Output nets */
wire t_1889,   t_1890;
/* u2_666 Output nets */
wire t_1891,   t_1892,   t_1893;
/* u2_667 Output nets */
wire t_1894,   t_1895,   t_1896;
/* u2_668 Output nets */
wire t_1897,   t_1898,   t_1899;
/* u2_669 Output nets */
wire t_1900,   t_1901,   t_1902;
/* u2_670 Output nets */
wire t_1903,   t_1904,   t_1905;
/* u2_671 Output nets */
wire t_1906,   t_1907,   t_1908;
/* u0_672 Output nets */
wire t_1909,   t_1910;
/* u2_673 Output nets */
wire t_1911,   t_1912,   t_1913;
/* u2_674 Output nets */
wire t_1914,   t_1915,   t_1916;
/* u2_675 Output nets */
wire t_1917,   t_1918,   t_1919;
/* u1_676 Output nets */
wire t_1920,   t_1921;
/* u2_677 Output nets */
wire t_1922,   t_1923,   t_1924;
/* u2_678 Output nets */
wire t_1925,   t_1926,   t_1927;
/* u2_679 Output nets */
wire t_1928,   t_1929,   t_1930;
/* u0_680 Output nets */
wire t_1931,   t_1932;
/* u2_681 Output nets */
wire t_1933,   t_1934,   t_1935;
/* u2_682 Output nets */
wire t_1936,   t_1937,   t_1938;
/* u2_683 Output nets */
wire t_1939,   t_1940,   t_1941;
/* u0_684 Output nets */
wire t_1942,   t_1943;
/* u2_685 Output nets */
wire t_1944,   t_1945,   t_1946;
/* u2_686 Output nets */
wire t_1947,   t_1948,   t_1949;
/* u2_687 Output nets */
wire t_1950,   t_1951,   t_1952;
/* u0_688 Output nets */
wire t_1953,   t_1954;
/* u2_689 Output nets */
wire t_1955,   t_1956,   t_1957;
/* u2_690 Output nets */
wire t_1958,   t_1959,   t_1960;
/* u2_691 Output nets */
wire t_1961,   t_1962,   t_1963;
/* u1_692 Output nets */
wire t_1964,   t_1965;
/* u2_693 Output nets */
wire t_1966,   t_1967,   t_1968;
/* u2_694 Output nets */
wire t_1969,   t_1970,   t_1971;
/* u2_695 Output nets */
wire t_1972,   t_1973,   t_1974;
/* u1_696 Output nets */
wire t_1975,   t_1976;
/* u2_697 Output nets */
wire t_1977,   t_1978,   t_1979;
/* u2_698 Output nets */
wire t_1980,   t_1981,   t_1982;
/* u2_699 Output nets */
wire t_1983,   t_1984,   t_1985;
/* u1_700 Output nets */
wire t_1986,   t_1987;
/* u2_701 Output nets */
wire t_1988,   t_1989,   t_1990;
/* u2_702 Output nets */
wire t_1991,   t_1992,   t_1993;
/* u2_703 Output nets */
wire t_1994,   t_1995,   t_1996;
/* u1_704 Output nets */
wire t_1997,   t_1998;
/* u2_705 Output nets */
wire t_1999,   t_2000,   t_2001;
/* u2_706 Output nets */
wire t_2002,   t_2003,   t_2004;
/* u2_707 Output nets */
wire t_2005,   t_2006,   t_2007;
/* u2_708 Output nets */
wire t_2008,   t_2009,   t_2010;
/* u2_709 Output nets */
wire t_2011,   t_2012,   t_2013;
/* u2_710 Output nets */
wire t_2014,   t_2015,   t_2016;
/* u2_711 Output nets */
wire t_2017,   t_2018,   t_2019;
/* u2_712 Output nets */
wire t_2020,   t_2021,   t_2022;
/* u2_713 Output nets */
wire t_2023,   t_2024,   t_2025;
/* u2_714 Output nets */
wire t_2026,   t_2027,   t_2028;
/* u2_715 Output nets */
wire t_2029,   t_2030,   t_2031;
/* u2_716 Output nets */
wire t_2032,   t_2033,   t_2034;
/* u2_717 Output nets */
wire t_2035,   t_2036,   t_2037;
/* u2_718 Output nets */
wire t_2038,   t_2039,   t_2040;
/* u2_719 Output nets */
wire t_2041,   t_2042,   t_2043;
/* u2_720 Output nets */
wire t_2044,   t_2045,   t_2046;
/* u2_721 Output nets */
wire t_2047,   t_2048,   t_2049;
/* u2_722 Output nets */
wire t_2050,   t_2051,   t_2052;
/* u2_723 Output nets */
wire t_2053,   t_2054,   t_2055;
/* u2_724 Output nets */
wire t_2056,   t_2057,   t_2058;
/* u2_725 Output nets */
wire t_2059,   t_2060,   t_2061;
/* u2_726 Output nets */
wire t_2062,   t_2063,   t_2064;
/* u2_727 Output nets */
wire t_2065,   t_2066,   t_2067;
/* u2_728 Output nets */
wire t_2068,   t_2069,   t_2070;
/* u2_729 Output nets */
wire t_2071,   t_2072,   t_2073;
/* u2_730 Output nets */
wire t_2074,   t_2075,   t_2076;
/* u2_731 Output nets */
wire t_2077,   t_2078,   t_2079;
/* u2_732 Output nets */
wire t_2080,   t_2081,   t_2082;
/* u2_733 Output nets */
wire t_2083,   t_2084,   t_2085;
/* u2_734 Output nets */
wire t_2086,   t_2087,   t_2088;
/* u2_735 Output nets */
wire t_2089,   t_2090,   t_2091;
/* u2_736 Output nets */
wire t_2092,   t_2093,   t_2094;
/* u2_737 Output nets */
wire t_2095,   t_2096,   t_2097;
/* u2_738 Output nets */
wire t_2098,   t_2099,   t_2100;
/* u2_739 Output nets */
wire t_2101,   t_2102,   t_2103;
/* u2_740 Output nets */
wire t_2104,   t_2105,   t_2106;
/* u2_741 Output nets */
wire t_2107,   t_2108,   t_2109;
/* u2_742 Output nets */
wire t_2110,   t_2111,   t_2112;
/* u2_743 Output nets */
wire t_2113,   t_2114,   t_2115;
/* u2_744 Output nets */
wire t_2116,   t_2117,   t_2118;
/* u2_745 Output nets */
wire t_2119,   t_2120,   t_2121;
/* u2_746 Output nets */
wire t_2122,   t_2123,   t_2124;
/* u2_747 Output nets */
wire t_2125,   t_2126,   t_2127;
/* u2_748 Output nets */
wire t_2128,   t_2129,   t_2130;
/* u2_749 Output nets */
wire t_2131,   t_2132,   t_2133;
/* u2_750 Output nets */
wire t_2134,   t_2135,   t_2136;
/* u2_751 Output nets */
wire t_2137,   t_2138,   t_2139;
/* u2_752 Output nets */
wire t_2140,   t_2141,   t_2142;
/* u2_753 Output nets */
wire t_2143,   t_2144,   t_2145;
/* u2_754 Output nets */
wire t_2146,   t_2147,   t_2148;
/* u2_755 Output nets */
wire t_2149,   t_2150,   t_2151;
/* u2_756 Output nets */
wire t_2152,   t_2153,   t_2154;
/* u2_757 Output nets */
wire t_2155,   t_2156,   t_2157;
/* u2_758 Output nets */
wire t_2158,   t_2159,   t_2160;
/* u2_759 Output nets */
wire t_2161,   t_2162,   t_2163;
/* u1_760 Output nets */
wire t_2164,   t_2165;
/* u2_761 Output nets */
wire t_2166,   t_2167,   t_2168;
/* u2_762 Output nets */
wire t_2169,   t_2170,   t_2171;
/* u2_763 Output nets */
wire t_2172,   t_2173,   t_2174;
/* u0_764 Output nets */
wire t_2175,   t_2176;
/* u2_765 Output nets */
wire t_2177,   t_2178,   t_2179;
/* u2_766 Output nets */
wire t_2180,   t_2181,   t_2182;
/* u2_767 Output nets */
wire t_2183,   t_2184,   t_2185;
/* u0_768 Output nets */
wire t_2186,   t_2187;
/* u2_769 Output nets */
wire t_2188,   t_2189,   t_2190;
/* u2_770 Output nets */
wire t_2191,   t_2192,   t_2193;
/* u2_771 Output nets */
wire t_2194,   t_2195,   t_2196;
/* u1_772 Output nets */
wire t_2197,   t_2198;
/* u2_773 Output nets */
wire t_2199,   t_2200,   t_2201;
/* u2_774 Output nets */
wire t_2202,   t_2203,   t_2204;
/* u2_775 Output nets */
wire t_2205,   t_2206,   t_2207;
/* u0_776 Output nets */
wire t_2208,   t_2209;
/* u2_777 Output nets */
wire t_2210,   t_2211,   t_2212;
/* u2_778 Output nets */
wire t_2213,   t_2214,   t_2215;
/* u2_779 Output nets */
wire t_2216,   t_2217,   t_2218;
/* u0_780 Output nets */
wire t_2219,   t_2220;
/* u2_781 Output nets */
wire t_2221,   t_2222,   t_2223;
/* u2_782 Output nets */
wire t_2224,   t_2225,   t_2226;
/* u2_783 Output nets */
wire t_2227,   t_2228,   t_2229;
/* u0_784 Output nets */
wire t_2230,   t_2231;
/* u2_785 Output nets */
wire t_2232,   t_2233,   t_2234;
/* u2_786 Output nets */
wire t_2235,   t_2236,   t_2237;
/* u2_787 Output nets */
wire t_2238,   t_2239,   t_2240;
/* u0_788 Output nets */
wire t_2241,   t_2242;
/* u2_789 Output nets */
wire t_2243,   t_2244,   t_2245;
/* u2_790 Output nets */
wire t_2246,   t_2247,   t_2248;
/* u2_791 Output nets */
wire t_2249,   t_2250,   t_2251;
/* u2_792 Output nets */
wire t_2252,   t_2253,   t_2254;
/* u2_793 Output nets */
wire t_2255,   t_2256,   t_2257;
/* u2_794 Output nets */
wire t_2258,   t_2259,   t_2260;
/* u2_795 Output nets */
wire t_2261,   t_2262,   t_2263;
/* u2_796 Output nets */
wire t_2264,   t_2265,   t_2266;
/* u2_797 Output nets */
wire t_2267,   t_2268,   t_2269;
/* u2_798 Output nets */
wire t_2270,   t_2271,   t_2272;
/* u2_799 Output nets */
wire t_2273,   t_2274,   t_2275;
/* u2_800 Output nets */
wire t_2276,   t_2277,   t_2278;
/* u2_801 Output nets */
wire t_2279,   t_2280,   t_2281;
/* u2_802 Output nets */
wire t_2282,   t_2283,   t_2284;
/* u2_803 Output nets */
wire t_2285,   t_2286,   t_2287;
/* u2_804 Output nets */
wire t_2288,   t_2289,   t_2290;
/* u2_805 Output nets */
wire t_2291,   t_2292,   t_2293;
/* u2_806 Output nets */
wire t_2294,   t_2295,   t_2296;
/* u2_807 Output nets */
wire t_2297,   t_2298,   t_2299;
/* u2_808 Output nets */
wire t_2300,   t_2301,   t_2302;
/* u2_809 Output nets */
wire t_2303,   t_2304,   t_2305;
/* u2_810 Output nets */
wire t_2306,   t_2307,   t_2308;
/* u2_811 Output nets */
wire t_2309,   t_2310,   t_2311;
/* u2_812 Output nets */
wire t_2312,   t_2313,   t_2314;
/* u2_813 Output nets */
wire t_2315,   t_2316,   t_2317;
/* u2_814 Output nets */
wire t_2318,   t_2319,   t_2320;
/* u1_815 Output nets */
wire t_2321,   t_2322;
/* u2_816 Output nets */
wire t_2323,   t_2324,   t_2325;
/* u2_817 Output nets */
wire t_2326,   t_2327,   t_2328;
/* u0_818 Output nets */
wire t_2329,   t_2330;
/* u2_819 Output nets */
wire t_2331,   t_2332,   t_2333;
/* u2_820 Output nets */
wire t_2334,   t_2335,   t_2336;
/* u0_821 Output nets */
wire t_2337,   t_2338;
/* u2_822 Output nets */
wire t_2339,   t_2340,   t_2341;
/* u2_823 Output nets */
wire t_2342,   t_2343,   t_2344;
/* u1_824 Output nets */
wire t_2345,   t_2346;
/* u2_825 Output nets */
wire t_2347,   t_2348,   t_2349;
/* u2_826 Output nets */
wire t_2350,   t_2351,   t_2352;
/* u0_827 Output nets */
wire t_2353,   t_2354;
/* u2_828 Output nets */
wire t_2355,   t_2356,   t_2357;
/* u2_829 Output nets */
wire t_2358,   t_2359,   t_2360;
/* u0_830 Output nets */
wire t_2361,   t_2362;
/* u2_831 Output nets */
wire t_2363,   t_2364,   t_2365;
/* u2_832 Output nets */
wire t_2366,   t_2367,   t_2368;
/* u0_833 Output nets */
wire t_2369,   t_2370;
/* u2_834 Output nets */
wire t_2371,   t_2372,   t_2373;
/* u2_835 Output nets */
wire t_2374,   t_2375,   t_2376;
/* u0_836 Output nets */
wire t_2377,   t_2378;
/* u2_837 Output nets */
wire t_2379,   t_2380,   t_2381;
/* u2_838 Output nets */
wire t_2382,   t_2383,   t_2384;
/* u2_839 Output nets */
wire t_2385,   t_2386,   t_2387;
/* u2_840 Output nets */
wire t_2388,   t_2389,   t_2390;
/* u2_841 Output nets */
wire t_2391,   t_2392,   t_2393;
/* u2_842 Output nets */
wire t_2394,   t_2395,   t_2396;
/* u2_843 Output nets */
wire t_2397,   t_2398,   t_2399;
/* u2_844 Output nets */
wire t_2400,   t_2401,   t_2402;
/* u2_845 Output nets */
wire t_2403,   t_2404,   t_2405;
/* u2_846 Output nets */
wire t_2406,   t_2407,   t_2408;
/* u2_847 Output nets */
wire t_2409,   t_2410,   t_2411;
/* u2_848 Output nets */
wire t_2412,   t_2413,   t_2414;
/* u2_849 Output nets */
wire t_2415,   t_2416,   t_2417;
/* u2_850 Output nets */
wire t_2418,   t_2419,   t_2420;
/* u2_851 Output nets */
wire t_2421,   t_2422,   t_2423;
/* u2_852 Output nets */
wire t_2424,   t_2425,   t_2426;
/* u2_853 Output nets */
wire t_2427,   t_2428,   t_2429;
/* u1_854 Output nets */
wire t_2430,   t_2431;
/* u2_855 Output nets */
wire t_2432,   t_2433,   t_2434;
/* u0_856 Output nets */
wire t_2435,   t_2436;
/* u2_857 Output nets */
wire t_2437,   t_2438,   t_2439;
/* u0_858 Output nets */
wire t_2440,   t_2441;
/* u2_859 Output nets */
wire t_2442,   t_2443,   t_2444;
/* u1_860 Output nets */
wire t_2445,   t_2446;
/* u2_861 Output nets */
wire t_2447,   t_2448,   t_2449;
/* u0_862 Output nets */
wire t_2450,   t_2451;
/* u2_863 Output nets */
wire t_2452,   t_2453,   t_2454;
/* u0_864 Output nets */
wire t_2455,   t_2456;
/* u2_865 Output nets */
wire t_2457,   t_2458,   t_2459;
/* u0_866 Output nets */
wire t_2460,   t_2461;
/* u2_867 Output nets */
wire t_2462,   t_2463,   t_2464;
/* u0_868 Output nets */
wire t_2465,   t_2466;
/* u2_869 Output nets */
wire t_2467,   t_2468,   t_2469;
/* u2_870 Output nets */
wire t_2470,   t_2471,   t_2472;
/* u2_871 Output nets */
wire t_2473,   t_2474,   t_2475;
/* u2_872 Output nets */
wire t_2476,   t_2477,   t_2478;
/* u2_873 Output nets */
wire t_2479,   t_2480,   t_2481;
/* u2_874 Output nets */
wire t_2482,   t_2483,   t_2484;
/* u2_875 Output nets */
wire t_2485,   t_2486,   t_2487;
/* u2_876 Output nets */
wire t_2488,   t_2489,   t_2490;
/* u1_877 Output nets */
wire t_2491,   t_2492;
/* u0_878 Output nets */
wire t_2493,   t_2494;
/* u0_879 Output nets */
wire t_2495,   t_2496;
/* u1_880 Output nets */
wire t_2497,   t_2498;
/* u0_881 Output nets */
wire t_2499,   t_2500;
/* u0_882 Output nets */
wire t_2501,   t_2502;
/* u0_883 Output nets */
wire t_2503;

/* compress stage 2 */
half_adder u0_569(.a(t_1), .b(s_1_0), .o(t_1631), .cout(t_1632));
half_adder u0_570(.a(t_4), .b(t_3), .o(t_1633), .cout(t_1634));
compressor_3_2 u1_571(.a(t_6), .b(t_5), .cin(s_4_3), .o(t_1635), .cout(t_1636));
half_adder u0_572(.a(t_8), .b(t_7), .o(t_1637), .cout(t_1638));
half_adder u0_573(.a(t_10), .b(t_9), .o(t_1639), .cout(t_1640));
half_adder u0_574(.a(t_13), .b(t_11), .o(t_1641), .cout(t_1642));
compressor_3_2 u1_575(.a(t_19), .b(t_16), .cin(t_14), .o(t_1643), .cout(t_1644));
compressor_3_2 u1_576(.a(t_20), .b(t_17), .cin(s_9_4), .o(t_1645), .cout(t_1646));
compressor_3_2 u1_577(.a(t_27), .b(t_24), .cin(t_22), .o(t_1647), .cout(t_1648));
compressor_3_2 u1_578(.a(t_29), .b(t_28), .cin(t_25), .o(t_1649), .cout(t_1650));
compressor_4_2 u2_579(.a(t_37), .b(t_34), .c(t_33), .d(t_30), .cin(s_12_7), .o(t_1651), .co(t_1652), .cout(t_1653));
compressor_4_2 u2_580(.a(t_42), .b(t_39), .c(t_38), .d(t_35), .cin(t_1653), .o(t_1654), .co(t_1655), .cout(t_1656));
compressor_4_2 u2_581(.a(t_47), .b(t_44), .c(t_43), .d(t_40), .cin(t_1656), .o(t_1657), .co(t_1658), .cout(t_1659));
compressor_4_2 u2_582(.a(t_53), .b(t_50), .c(t_48), .d(t_45), .cin(t_1659), .o(t_1660), .co(t_1661), .cout(t_1662));
compressor_4_2 u2_583(.a(t_59), .b(t_56), .c(t_54), .d(t_51), .cin(t_1662), .o(t_1663), .co(t_1664), .cout(t_1665));
compressor_4_2 u2_584(.a(t_63), .b(t_60), .c(t_57), .d(s_17_8), .cin(t_1665), .o(t_1666), .co(t_1667), .cout(t_1668));
half_adder u0_585(.a(t_67), .b(t_64), .o(t_1669), .cout(t_1670));
compressor_4_2 u2_586(.a(t_73), .b(t_70), .c(t_68), .d(t_65), .cin(t_1668), .o(t_1671), .co(t_1672), .cout(t_1673));
compressor_4_2 u2_587(.a(t_78), .b(t_77), .c(t_74), .d(t_71), .cin(t_1673), .o(t_1674), .co(t_1675), .cout(t_1676));
half_adder u0_588(.a(t_84), .b(t_81), .o(t_1677), .cout(t_1678));
compressor_4_2 u2_589(.a(t_85), .b(t_82), .c(t_79), .d(s_20_11), .cin(t_1676), .o(t_1679), .co(t_1680), .cout(t_1681));
compressor_3_2 u1_590(.a(t_92), .b(t_89), .cin(t_86), .o(t_1682), .cout(t_1683));
compressor_4_2 u2_591(.a(t_94), .b(t_93), .c(t_90), .d(t_87), .cin(t_1681), .o(t_1684), .co(t_1685), .cout(t_1686));
half_adder u0_592(.a(t_100), .b(t_97), .o(t_1687), .cout(t_1688));
compressor_4_2 u2_593(.a(t_102), .b(t_101), .c(t_98), .d(t_95), .cin(t_1686), .o(t_1689), .co(t_1690), .cout(t_1691));
half_adder u0_594(.a(t_108), .b(t_105), .o(t_1692), .cout(t_1693));
compressor_4_2 u2_595(.a(t_111), .b(t_109), .c(t_106), .d(t_103), .cin(t_1691), .o(t_1694), .co(t_1695), .cout(t_1696));
half_adder u0_596(.a(t_117), .b(t_114), .o(t_1697), .cout(t_1698));
compressor_4_2 u2_597(.a(t_120), .b(t_118), .c(t_115), .d(t_112), .cin(t_1696), .o(t_1699), .co(t_1700), .cout(t_1701));
compressor_3_2 u1_598(.a(t_129), .b(t_126), .cin(t_123), .o(t_1702), .cout(t_1703));
compressor_4_2 u2_599(.a(t_127), .b(t_124), .c(t_121), .d(s_25_12), .cin(t_1701), .o(t_1704), .co(t_1705), .cout(t_1706));
compressor_3_2 u1_600(.a(t_134), .b(t_131), .cin(t_130), .o(t_1707), .cout(t_1708));
compressor_4_2 u2_601(.a(t_140), .b(t_138), .c(t_135), .d(t_132), .cin(t_1706), .o(t_1709), .co(t_1710), .cout(t_1711));
compressor_3_2 u1_602(.a(t_149), .b(t_146), .cin(t_143), .o(t_1712), .cout(t_1713));
compressor_4_2 u2_603(.a(t_150), .b(t_147), .c(t_144), .d(t_141), .cin(t_1711), .o(t_1714), .co(t_1715), .cout(t_1716));
compressor_3_2 u1_604(.a(t_157), .b(t_154), .cin(t_151), .o(t_1717), .cout(t_1718));
compressor_4_2 u2_605(.a(t_158), .b(t_155), .c(t_152), .d(s_28_15), .cin(t_1716), .o(t_1719), .co(t_1720), .cout(t_1721));
compressor_4_2 u2_606(.a(t_171), .b(t_168), .c(t_165), .d(t_162), .cin(t_161), .o(t_1722), .co(t_1723), .cout(t_1724));
compressor_4_2 u2_607(.a(t_172), .b(t_169), .c(t_166), .d(t_163), .cin(t_1721), .o(t_1725), .co(t_1726), .cout(t_1727));
compressor_4_2 u2_608(.a(t_182), .b(t_179), .c(t_176), .d(t_173), .cin(t_1724), .o(t_1728), .co(t_1729), .cout(t_1730));
compressor_4_2 u2_609(.a(t_183), .b(t_180), .c(t_177), .d(t_174), .cin(t_1727), .o(t_1731), .co(t_1732), .cout(t_1733));
compressor_4_2 u2_610(.a(t_193), .b(t_190), .c(t_187), .d(t_184), .cin(t_1730), .o(t_1734), .co(t_1735), .cout(t_1736));
compressor_4_2 u2_611(.a(t_194), .b(t_191), .c(t_188), .d(t_185), .cin(t_1733), .o(t_1737), .co(t_1738), .cout(t_1739));
compressor_4_2 u2_612(.a(t_205), .b(t_202), .c(t_199), .d(t_196), .cin(t_1736), .o(t_1740), .co(t_1741), .cout(t_1742));
compressor_4_2 u2_613(.a(t_206), .b(t_203), .c(t_200), .d(t_197), .cin(t_1739), .o(t_1743), .co(t_1744), .cout(t_1745));
compressor_4_2 u2_614(.a(t_217), .b(t_214), .c(t_211), .d(t_208), .cin(t_1742), .o(t_1746), .co(t_1747), .cout(t_1748));
compressor_4_2 u2_615(.a(t_215), .b(t_212), .c(t_209), .d(s_33_16), .cin(t_1745), .o(t_1749), .co(t_1750), .cout(t_1751));
compressor_4_2 u2_616(.a(t_225), .b(t_222), .c(t_221), .d(t_218), .cin(t_1748), .o(t_1752), .co(t_1753), .cout(t_1754));
half_adder u0_617(.a(t_231), .b(t_228), .o(t_1755), .cout(t_1756));
compressor_4_2 u2_618(.a(t_232), .b(t_229), .c(t_226), .d(t_223), .cin(t_1751), .o(t_1757), .co(t_1758), .cout(t_1759));
compressor_4_2 u2_619(.a(t_243), .b(t_240), .c(t_237), .d(t_234), .cin(t_1754), .o(t_1760), .co(t_1761), .cout(t_1762));
compressor_4_2 u2_620(.a(t_244), .b(t_241), .c(t_238), .d(t_235), .cin(t_1759), .o(t_1763), .co(t_1764), .cout(t_1765));
compressor_4_2 u2_621(.a(t_254), .b(t_251), .c(t_248), .d(t_247), .cin(t_1762), .o(t_1766), .co(t_1767), .cout(t_1768));
half_adder u0_622(.a(t_260), .b(t_257), .o(t_1769), .cout(t_1770));
compressor_4_2 u2_623(.a(t_255), .b(t_252), .c(t_249), .d(s_36_19), .cin(t_1765), .o(t_1771), .co(t_1772), .cout(t_1773));
compressor_4_2 u2_624(.a(t_265), .b(t_262), .c(t_261), .d(t_258), .cin(t_1768), .o(t_1774), .co(t_1775), .cout(t_1776));
compressor_3_2 u1_625(.a(t_274), .b(t_271), .cin(t_268), .o(t_1777), .cout(t_1778));
compressor_4_2 u2_626(.a(t_272), .b(t_269), .c(t_266), .d(t_263), .cin(t_1773), .o(t_1779), .co(t_1780), .cout(t_1781));
compressor_4_2 u2_627(.a(t_282), .b(t_279), .c(t_276), .d(t_275), .cin(t_1776), .o(t_1782), .co(t_1783), .cout(t_1784));
half_adder u0_628(.a(t_288), .b(t_285), .o(t_1785), .cout(t_1786));
compressor_4_2 u2_629(.a(t_286), .b(t_283), .c(t_280), .d(t_277), .cin(t_1781), .o(t_1787), .co(t_1788), .cout(t_1789));
compressor_4_2 u2_630(.a(t_296), .b(t_293), .c(t_290), .d(t_289), .cin(t_1784), .o(t_1790), .co(t_1791), .cout(t_1792));
half_adder u0_631(.a(t_302), .b(t_299), .o(t_1793), .cout(t_1794));
compressor_4_2 u2_632(.a(t_300), .b(t_297), .c(t_294), .d(t_291), .cin(t_1789), .o(t_1795), .co(t_1796), .cout(t_1797));
compressor_4_2 u2_633(.a(t_311), .b(t_308), .c(t_305), .d(t_303), .cin(t_1792), .o(t_1798), .co(t_1799), .cout(t_1800));
half_adder u0_634(.a(t_317), .b(t_314), .o(t_1801), .cout(t_1802));
compressor_4_2 u2_635(.a(t_315), .b(t_312), .c(t_309), .d(t_306), .cin(t_1797), .o(t_1803), .co(t_1804), .cout(t_1805));
compressor_4_2 u2_636(.a(t_326), .b(t_323), .c(t_320), .d(t_318), .cin(t_1800), .o(t_1806), .co(t_1807), .cout(t_1808));
compressor_3_2 u1_637(.a(t_335), .b(t_332), .cin(t_329), .o(t_1809), .cout(t_1810));
compressor_4_2 u2_638(.a(t_327), .b(t_324), .c(t_321), .d(s_41_20), .cin(t_1805), .o(t_1811), .co(t_1812), .cout(t_1813));
compressor_4_2 u2_639(.a(t_337), .b(t_336), .c(t_333), .d(t_330), .cin(t_1808), .o(t_1814), .co(t_1815), .cout(t_1816));
compressor_3_2 u1_640(.a(t_346), .b(t_343), .cin(t_340), .o(t_1817), .cout(t_1818));
compressor_4_2 u2_641(.a(t_347), .b(t_344), .c(t_341), .d(t_338), .cin(t_1813), .o(t_1819), .co(t_1820), .cout(t_1821));
compressor_4_2 u2_642(.a(t_358), .b(t_355), .c(t_352), .d(t_350), .cin(t_1816), .o(t_1822), .co(t_1823), .cout(t_1824));
compressor_3_2 u1_643(.a(t_367), .b(t_364), .cin(t_361), .o(t_1825), .cout(t_1826));
compressor_4_2 u2_644(.a(t_362), .b(t_359), .c(t_356), .d(t_353), .cin(t_1821), .o(t_1827), .co(t_1828), .cout(t_1829));
compressor_4_2 u2_645(.a(t_372), .b(t_369), .c(t_368), .d(t_365), .cin(t_1824), .o(t_1830), .co(t_1831), .cout(t_1832));
compressor_3_2 u1_646(.a(t_381), .b(t_378), .cin(t_375), .o(t_1833), .cout(t_1834));
compressor_4_2 u2_647(.a(t_376), .b(t_373), .c(t_370), .d(s_44_23), .cin(t_1829), .o(t_1835), .co(t_1836), .cout(t_1837));
compressor_4_2 u2_648(.a(t_386), .b(t_385), .c(t_382), .d(t_379), .cin(t_1832), .o(t_1838), .co(t_1839), .cout(t_1840));
compressor_4_2 u2_649(.a(t_401), .b(t_398), .c(t_395), .d(t_392), .cin(t_389), .o(t_1841), .co(t_1842), .cout(t_1843));
compressor_4_2 u2_650(.a(t_396), .b(t_393), .c(t_390), .d(t_387), .cin(t_1837), .o(t_1844), .co(t_1845), .cout(t_1846));
compressor_4_2 u2_651(.a(t_406), .b(t_403), .c(t_402), .d(t_399), .cin(t_1840), .o(t_1847), .co(t_1848), .cout(t_1849));
compressor_4_2 u2_652(.a(t_418), .b(t_415), .c(t_412), .d(t_409), .cin(t_1843), .o(t_1850), .co(t_1851), .cout(t_1852));
compressor_4_2 u2_653(.a(t_413), .b(t_410), .c(t_407), .d(t_404), .cin(t_1846), .o(t_1853), .co(t_1854), .cout(t_1855));
compressor_4_2 u2_654(.a(t_423), .b(t_420), .c(t_419), .d(t_416), .cin(t_1849), .o(t_1856), .co(t_1857), .cout(t_1858));
compressor_4_2 u2_655(.a(t_435), .b(t_432), .c(t_429), .d(t_426), .cin(t_1852), .o(t_1859), .co(t_1860), .cout(t_1861));
compressor_4_2 u2_656(.a(t_430), .b(t_427), .c(t_424), .d(t_421), .cin(t_1855), .o(t_1862), .co(t_1863), .cout(t_1864));
compressor_4_2 u2_657(.a(t_441), .b(t_438), .c(t_436), .d(t_433), .cin(t_1858), .o(t_1865), .co(t_1866), .cout(t_1867));
compressor_4_2 u2_658(.a(t_453), .b(t_450), .c(t_447), .d(t_444), .cin(t_1861), .o(t_1868), .co(t_1869), .cout(t_1870));
compressor_4_2 u2_659(.a(t_448), .b(t_445), .c(t_442), .d(t_439), .cin(t_1864), .o(t_1871), .co(t_1872), .cout(t_1873));
compressor_4_2 u2_660(.a(t_459), .b(t_456), .c(t_454), .d(t_451), .cin(t_1867), .o(t_1874), .co(t_1875), .cout(t_1876));
compressor_4_2 u2_661(.a(t_471), .b(t_468), .c(t_465), .d(t_462), .cin(t_1870), .o(t_1877), .co(t_1878), .cout(t_1879));
compressor_4_2 u2_662(.a(t_463), .b(t_460), .c(t_457), .d(s_49_24), .cin(t_1873), .o(t_1880), .co(t_1881), .cout(t_1882));
compressor_4_2 u2_663(.a(t_475), .b(t_472), .c(t_469), .d(t_466), .cin(t_1876), .o(t_1883), .co(t_1884), .cout(t_1885));
compressor_4_2 u2_664(.a(t_485), .b(t_482), .c(t_479), .d(t_476), .cin(t_1879), .o(t_1886), .co(t_1887), .cout(t_1888));
half_adder u0_665(.a(t_491), .b(t_488), .o(t_1889), .cout(t_1890));
compressor_4_2 u2_666(.a(t_486), .b(t_483), .c(t_480), .d(t_477), .cin(t_1882), .o(t_1891), .co(t_1892), .cout(t_1893));
compressor_4_2 u2_667(.a(t_497), .b(t_494), .c(t_492), .d(t_489), .cin(t_1885), .o(t_1894), .co(t_1895), .cout(t_1896));
compressor_4_2 u2_668(.a(t_509), .b(t_506), .c(t_503), .d(t_500), .cin(t_1888), .o(t_1897), .co(t_1898), .cout(t_1899));
compressor_4_2 u2_669(.a(t_504), .b(t_501), .c(t_498), .d(t_495), .cin(t_1893), .o(t_1900), .co(t_1901), .cout(t_1902));
compressor_4_2 u2_670(.a(t_514), .b(t_513), .c(t_510), .d(t_507), .cin(t_1896), .o(t_1903), .co(t_1904), .cout(t_1905));
compressor_4_2 u2_671(.a(t_526), .b(t_523), .c(t_520), .d(t_517), .cin(t_1899), .o(t_1906), .co(t_1907), .cout(t_1908));
half_adder u0_672(.a(t_532), .b(t_529), .o(t_1909), .cout(t_1910));
compressor_4_2 u2_673(.a(t_521), .b(t_518), .c(t_515), .d(s_52_27), .cin(t_1902), .o(t_1911), .co(t_1912), .cout(t_1913));
compressor_4_2 u2_674(.a(t_533), .b(t_530), .c(t_527), .d(t_524), .cin(t_1905), .o(t_1914), .co(t_1915), .cout(t_1916));
compressor_4_2 u2_675(.a(t_543), .b(t_540), .c(t_537), .d(t_534), .cin(t_1908), .o(t_1917), .co(t_1918), .cout(t_1919));
compressor_3_2 u1_676(.a(t_552), .b(t_549), .cin(t_546), .o(t_1920), .cout(t_1921));
compressor_4_2 u2_677(.a(t_544), .b(t_541), .c(t_538), .d(t_535), .cin(t_1913), .o(t_1922), .co(t_1923), .cout(t_1924));
compressor_4_2 u2_678(.a(t_554), .b(t_553), .c(t_550), .d(t_547), .cin(t_1916), .o(t_1925), .co(t_1926), .cout(t_1927));
compressor_4_2 u2_679(.a(t_566), .b(t_563), .c(t_560), .d(t_557), .cin(t_1919), .o(t_1928), .co(t_1929), .cout(t_1930));
half_adder u0_680(.a(t_572), .b(t_569), .o(t_1931), .cout(t_1932));
compressor_4_2 u2_681(.a(t_564), .b(t_561), .c(t_558), .d(t_555), .cin(t_1924), .o(t_1933), .co(t_1934), .cout(t_1935));
compressor_4_2 u2_682(.a(t_574), .b(t_573), .c(t_570), .d(t_567), .cin(t_1927), .o(t_1936), .co(t_1937), .cout(t_1938));
compressor_4_2 u2_683(.a(t_586), .b(t_583), .c(t_580), .d(t_577), .cin(t_1930), .o(t_1939), .co(t_1940), .cout(t_1941));
half_adder u0_684(.a(t_592), .b(t_589), .o(t_1942), .cout(t_1943));
compressor_4_2 u2_685(.a(t_584), .b(t_581), .c(t_578), .d(t_575), .cin(t_1935), .o(t_1944), .co(t_1945), .cout(t_1946));
compressor_4_2 u2_686(.a(t_595), .b(t_593), .c(t_590), .d(t_587), .cin(t_1938), .o(t_1947), .co(t_1948), .cout(t_1949));
compressor_4_2 u2_687(.a(t_607), .b(t_604), .c(t_601), .d(t_598), .cin(t_1941), .o(t_1950), .co(t_1951), .cout(t_1952));
half_adder u0_688(.a(t_613), .b(t_610), .o(t_1953), .cout(t_1954));
compressor_4_2 u2_689(.a(t_605), .b(t_602), .c(t_599), .d(t_596), .cin(t_1946), .o(t_1955), .co(t_1956), .cout(t_1957));
compressor_4_2 u2_690(.a(t_616), .b(t_614), .c(t_611), .d(t_608), .cin(t_1949), .o(t_1958), .co(t_1959), .cout(t_1960));
compressor_4_2 u2_691(.a(t_628), .b(t_625), .c(t_622), .d(t_619), .cin(t_1952), .o(t_1961), .co(t_1962), .cout(t_1963));
compressor_3_2 u1_692(.a(t_637), .b(t_634), .cin(t_631), .o(t_1964), .cout(t_1965));
compressor_4_2 u2_693(.a(t_623), .b(t_620), .c(t_617), .d(s_57_28), .cin(t_1957), .o(t_1966), .co(t_1967), .cout(t_1968));
compressor_4_2 u2_694(.a(t_635), .b(t_632), .c(t_629), .d(t_626), .cin(t_1960), .o(t_1969), .co(t_1970), .cout(t_1971));
compressor_4_2 u2_695(.a(t_645), .b(t_642), .c(t_639), .d(t_638), .cin(t_1963), .o(t_1972), .co(t_1973), .cout(t_1974));
compressor_3_2 u1_696(.a(t_654), .b(t_651), .cin(t_648), .o(t_1975), .cout(t_1976));
compressor_4_2 u2_697(.a(t_649), .b(t_646), .c(t_643), .d(t_640), .cin(t_1968), .o(t_1977), .co(t_1978), .cout(t_1979));
compressor_4_2 u2_698(.a(t_660), .b(t_658), .c(t_655), .d(t_652), .cin(t_1971), .o(t_1980), .co(t_1981), .cout(t_1982));
compressor_4_2 u2_699(.a(t_672), .b(t_669), .c(t_666), .d(t_663), .cin(t_1974), .o(t_1983), .co(t_1984), .cout(t_1985));
compressor_3_2 u1_700(.a(t_681), .b(t_678), .cin(t_675), .o(t_1986), .cout(t_1987));
compressor_4_2 u2_701(.a(t_670), .b(t_667), .c(t_664), .d(t_661), .cin(t_1979), .o(t_1988), .co(t_1989), .cout(t_1990));
compressor_4_2 u2_702(.a(t_682), .b(t_679), .c(t_676), .d(t_673), .cin(t_1982), .o(t_1991), .co(t_1992), .cout(t_1993));
compressor_4_2 u2_703(.a(t_692), .b(t_689), .c(t_686), .d(t_683), .cin(t_1985), .o(t_1994), .co(t_1995), .cout(t_1996));
compressor_3_2 u1_704(.a(t_701), .b(t_698), .cin(t_695), .o(t_1997), .cout(t_1998));
compressor_4_2 u2_705(.a(t_690), .b(t_687), .c(t_684), .d(s_60_31), .cin(t_1990), .o(t_1999), .co(t_2000), .cout(t_2001));
compressor_4_2 u2_706(.a(t_702), .b(t_699), .c(t_696), .d(t_693), .cin(t_1993), .o(t_2002), .co(t_2003), .cout(t_2004));
compressor_4_2 u2_707(.a(t_712), .b(t_709), .c(t_706), .d(t_705), .cin(t_1996), .o(t_2005), .co(t_2006), .cout(t_2007));
compressor_4_2 u2_708(.a(t_727), .b(t_724), .c(t_721), .d(t_718), .cin(t_715), .o(t_2008), .co(t_2009), .cout(t_2010));
compressor_4_2 u2_709(.a(t_716), .b(t_713), .c(t_710), .d(t_707), .cin(t_2001), .o(t_2011), .co(t_2012), .cout(t_2013));
compressor_4_2 u2_710(.a(t_728), .b(t_725), .c(t_722), .d(t_719), .cin(t_2004), .o(t_2014), .co(t_2015), .cout(t_2016));
compressor_4_2 u2_711(.a(t_738), .b(t_735), .c(t_732), .d(t_729), .cin(t_2007), .o(t_2017), .co(t_2018), .cout(t_2019));
compressor_4_2 u2_712(.a(t_750), .b(t_747), .c(t_744), .d(t_741), .cin(t_2010), .o(t_2020), .co(t_2021), .cout(t_2022));
compressor_4_2 u2_713(.a(t_739), .b(t_736), .c(t_733), .d(t_730), .cin(t_2013), .o(t_2023), .co(t_2024), .cout(t_2025));
compressor_4_2 u2_714(.a(t_751), .b(t_748), .c(t_745), .d(t_742), .cin(t_2016), .o(t_2026), .co(t_2027), .cout(t_2028));
compressor_4_2 u2_715(.a(t_761), .b(t_758), .c(t_755), .d(t_752), .cin(t_2019), .o(t_2029), .co(t_2030), .cout(t_2031));
compressor_4_2 u2_716(.a(t_773), .b(t_770), .c(t_767), .d(t_764), .cin(t_2022), .o(t_2032), .co(t_2033), .cout(t_2034));
compressor_4_2 u2_717(.a(t_762), .b(t_759), .c(t_756), .d(t_753), .cin(t_2025), .o(t_2035), .co(t_2036), .cout(t_2037));
compressor_4_2 u2_718(.a(t_774), .b(t_771), .c(t_768), .d(t_765), .cin(t_2028), .o(t_2038), .co(t_2039), .cout(t_2040));
compressor_4_2 u2_719(.a(t_785), .b(t_782), .c(t_779), .d(t_776), .cin(t_2031), .o(t_2041), .co(t_2042), .cout(t_2043));
compressor_4_2 u2_720(.a(t_797), .b(t_794), .c(t_791), .d(t_788), .cin(t_2034), .o(t_2044), .co(t_2045), .cout(t_2046));
compressor_4_2 u2_721(.a(t_783), .b(t_780), .c(t_777), .d(s_64_32), .cin(t_2037), .o(t_2047), .co(t_2048), .cout(t_2049));
compressor_4_2 u2_722(.a(t_795), .b(t_792), .c(t_789), .d(t_786), .cin(t_2040), .o(t_2050), .co(t_2051), .cout(t_2052));
compressor_4_2 u2_723(.a(t_806), .b(t_803), .c(t_800), .d(t_798), .cin(t_2043), .o(t_2053), .co(t_2054), .cout(t_2055));
compressor_4_2 u2_724(.a(t_818), .b(t_815), .c(t_812), .d(t_809), .cin(t_2046), .o(t_2056), .co(t_2057), .cout(t_2058));
compressor_4_2 u2_725(.a(t_807), .b(t_804), .c(t_801), .d(s_65_32), .cin(t_2049), .o(t_2059), .co(t_2060), .cout(t_2061));
compressor_4_2 u2_726(.a(t_819), .b(t_816), .c(t_813), .d(t_810), .cin(t_2052), .o(t_2062), .co(t_2063), .cout(t_2064));
compressor_4_2 u2_727(.a(t_830), .b(t_827), .c(t_824), .d(t_822), .cin(t_2055), .o(t_2065), .co(t_2066), .cout(t_2067));
compressor_4_2 u2_728(.a(t_842), .b(t_839), .c(t_836), .d(t_833), .cin(t_2058), .o(t_2068), .co(t_2069), .cout(t_2070));
compressor_4_2 u2_729(.a(t_834), .b(t_831), .c(t_828), .d(t_825), .cin(t_2061), .o(t_2071), .co(t_2072), .cout(t_2073));
compressor_4_2 u2_730(.a(t_846), .b(t_843), .c(t_840), .d(t_837), .cin(t_2064), .o(t_2074), .co(t_2075), .cout(t_2076));
compressor_4_2 u2_731(.a(t_857), .b(t_854), .c(t_851), .d(t_848), .cin(t_2067), .o(t_2077), .co(t_2078), .cout(t_2079));
compressor_4_2 u2_732(.a(t_869), .b(t_866), .c(t_863), .d(t_860), .cin(t_2070), .o(t_2080), .co(t_2081), .cout(t_2082));
compressor_4_2 u2_733(.a(t_858), .b(t_855), .c(t_852), .d(t_849), .cin(t_2073), .o(t_2083), .co(t_2084), .cout(t_2085));
compressor_4_2 u2_734(.a(t_870), .b(t_867), .c(t_864), .d(t_861), .cin(t_2076), .o(t_2086), .co(t_2087), .cout(t_2088));
compressor_4_2 u2_735(.a(t_881), .b(t_878), .c(t_875), .d(t_872), .cin(t_2079), .o(t_2089), .co(t_2090), .cout(t_2091));
compressor_4_2 u2_736(.a(t_893), .b(t_890), .c(t_887), .d(t_884), .cin(t_2082), .o(t_2092), .co(t_2093), .cout(t_2094));
compressor_4_2 u2_737(.a(t_879), .b(t_876), .c(t_873), .d(s_68_30), .cin(t_2085), .o(t_2095), .co(t_2096), .cout(t_2097));
compressor_4_2 u2_738(.a(t_891), .b(t_888), .c(t_885), .d(t_882), .cin(t_2088), .o(t_2098), .co(t_2099), .cout(t_2100));
compressor_4_2 u2_739(.a(t_902), .b(t_899), .c(t_896), .d(t_894), .cin(t_2091), .o(t_2101), .co(t_2102), .cout(t_2103));
compressor_4_2 u2_740(.a(t_914), .b(t_911), .c(t_908), .d(t_905), .cin(t_2094), .o(t_2104), .co(t_2105), .cout(t_2106));
compressor_4_2 u2_741(.a(t_906), .b(t_903), .c(t_900), .d(t_897), .cin(t_2097), .o(t_2107), .co(t_2108), .cout(t_2109));
compressor_4_2 u2_742(.a(t_918), .b(t_915), .c(t_912), .d(t_909), .cin(t_2100), .o(t_2110), .co(t_2111), .cout(t_2112));
compressor_4_2 u2_743(.a(t_928), .b(t_925), .c(t_922), .d(t_919), .cin(t_2103), .o(t_2113), .co(t_2114), .cout(t_2115));
compressor_4_2 u2_744(.a(t_940), .b(t_937), .c(t_934), .d(t_931), .cin(t_2106), .o(t_2116), .co(t_2117), .cout(t_2118));
compressor_4_2 u2_745(.a(t_929), .b(t_926), .c(t_923), .d(t_920), .cin(t_2109), .o(t_2119), .co(t_2120), .cout(t_2121));
compressor_4_2 u2_746(.a(t_941), .b(t_938), .c(t_935), .d(t_932), .cin(t_2112), .o(t_2122), .co(t_2123), .cout(t_2124));
compressor_4_2 u2_747(.a(t_951), .b(t_948), .c(t_945), .d(t_942), .cin(t_2115), .o(t_2125), .co(t_2126), .cout(t_2127));
compressor_4_2 u2_748(.a(t_963), .b(t_960), .c(t_957), .d(t_954), .cin(t_2118), .o(t_2128), .co(t_2129), .cout(t_2130));
compressor_4_2 u2_749(.a(t_952), .b(t_949), .c(t_946), .d(t_943), .cin(t_2121), .o(t_2131), .co(t_2132), .cout(t_2133));
compressor_4_2 u2_750(.a(t_964), .b(t_961), .c(t_958), .d(t_955), .cin(t_2124), .o(t_2134), .co(t_2135), .cout(t_2136));
compressor_4_2 u2_751(.a(t_974), .b(t_971), .c(t_968), .d(t_965), .cin(t_2127), .o(t_2137), .co(t_2138), .cout(t_2139));
compressor_4_2 u2_752(.a(t_986), .b(t_983), .c(t_980), .d(t_977), .cin(t_2130), .o(t_2140), .co(t_2141), .cout(t_2142));
compressor_4_2 u2_753(.a(t_972), .b(t_969), .c(t_966), .d(s_72_28), .cin(t_2133), .o(t_2143), .co(t_2144), .cout(t_2145));
compressor_4_2 u2_754(.a(t_984), .b(t_981), .c(t_978), .d(t_975), .cin(t_2136), .o(t_2146), .co(t_2147), .cout(t_2148));
compressor_4_2 u2_755(.a(t_994), .b(t_991), .c(t_988), .d(t_987), .cin(t_2139), .o(t_2149), .co(t_2150), .cout(t_2151));
compressor_4_2 u2_756(.a(t_1006), .b(t_1003), .c(t_1000), .d(t_997), .cin(t_2142), .o(t_2152), .co(t_2153), .cout(t_2154));
compressor_4_2 u2_757(.a(t_995), .b(t_992), .c(t_989), .d(s_73_28), .cin(t_2145), .o(t_2155), .co(t_2156), .cout(t_2157));
compressor_4_2 u2_758(.a(t_1007), .b(t_1004), .c(t_1001), .d(t_998), .cin(t_2148), .o(t_2158), .co(t_2159), .cout(t_2160));
compressor_4_2 u2_759(.a(t_1018), .b(t_1015), .c(t_1012), .d(t_1009), .cin(t_2151), .o(t_2161), .co(t_2162), .cout(t_2163));
compressor_3_2 u1_760(.a(t_1024), .b(t_1021), .cin(t_2154), .o(t_2164), .cout(t_2165));
compressor_4_2 u2_761(.a(t_1019), .b(t_1016), .c(t_1013), .d(t_1010), .cin(t_2157), .o(t_2166), .co(t_2167), .cout(t_2168));
compressor_4_2 u2_762(.a(t_1030), .b(t_1028), .c(t_1025), .d(t_1022), .cin(t_2160), .o(t_2169), .co(t_2170), .cout(t_2171));
compressor_4_2 u2_763(.a(t_1042), .b(t_1039), .c(t_1036), .d(t_1033), .cin(t_2163), .o(t_2172), .co(t_2173), .cout(t_2174));
half_adder u0_764(.a(t_1048), .b(t_1045), .o(t_2175), .cout(t_2176));
compressor_4_2 u2_765(.a(t_1040), .b(t_1037), .c(t_1034), .d(t_1031), .cin(t_2168), .o(t_2177), .co(t_2178), .cout(t_2179));
compressor_4_2 u2_766(.a(t_1051), .b(t_1049), .c(t_1046), .d(t_1043), .cin(t_2171), .o(t_2180), .co(t_2181), .cout(t_2182));
compressor_4_2 u2_767(.a(t_1063), .b(t_1060), .c(t_1057), .d(t_1054), .cin(t_2174), .o(t_2183), .co(t_2184), .cout(t_2185));
half_adder u0_768(.a(t_1069), .b(t_1066), .o(t_2186), .cout(t_2187));
compressor_4_2 u2_769(.a(t_1058), .b(t_1055), .c(t_1052), .d(s_76_26), .cin(t_2179), .o(t_2188), .co(t_2189), .cout(t_2190));
compressor_4_2 u2_770(.a(t_1070), .b(t_1067), .c(t_1064), .d(t_1061), .cin(t_2182), .o(t_2191), .co(t_2192), .cout(t_2193));
compressor_4_2 u2_771(.a(t_1081), .b(t_1078), .c(t_1075), .d(t_1072), .cin(t_2185), .o(t_2194), .co(t_2195), .cout(t_2196));
compressor_3_2 u1_772(.a(t_1090), .b(t_1087), .cin(t_1084), .o(t_2197), .cout(t_2198));
compressor_4_2 u2_773(.a(t_1082), .b(t_1079), .c(t_1076), .d(t_1073), .cin(t_2190), .o(t_2199), .co(t_2200), .cout(t_2201));
compressor_4_2 u2_774(.a(t_1092), .b(t_1091), .c(t_1088), .d(t_1085), .cin(t_2193), .o(t_2202), .co(t_2203), .cout(t_2204));
compressor_4_2 u2_775(.a(t_1104), .b(t_1101), .c(t_1098), .d(t_1095), .cin(t_2196), .o(t_2205), .co(t_2206), .cout(t_2207));
half_adder u0_776(.a(t_1110), .b(t_1107), .o(t_2208), .cout(t_2209));
compressor_4_2 u2_777(.a(t_1102), .b(t_1099), .c(t_1096), .d(t_1093), .cin(t_2201), .o(t_2210), .co(t_2211), .cout(t_2212));
compressor_4_2 u2_778(.a(t_1112), .b(t_1111), .c(t_1108), .d(t_1105), .cin(t_2204), .o(t_2213), .co(t_2214), .cout(t_2215));
compressor_4_2 u2_779(.a(t_1124), .b(t_1121), .c(t_1118), .d(t_1115), .cin(t_2207), .o(t_2216), .co(t_2217), .cout(t_2218));
half_adder u0_780(.a(t_1130), .b(t_1127), .o(t_2219), .cout(t_2220));
compressor_4_2 u2_781(.a(t_1122), .b(t_1119), .c(t_1116), .d(t_1113), .cin(t_2212), .o(t_2221), .co(t_2222), .cout(t_2223));
compressor_4_2 u2_782(.a(t_1132), .b(t_1131), .c(t_1128), .d(t_1125), .cin(t_2215), .o(t_2224), .co(t_2225), .cout(t_2226));
compressor_4_2 u2_783(.a(t_1144), .b(t_1141), .c(t_1138), .d(t_1135), .cin(t_2218), .o(t_2227), .co(t_2228), .cout(t_2229));
half_adder u0_784(.a(t_1150), .b(t_1147), .o(t_2230), .cout(t_2231));
compressor_4_2 u2_785(.a(t_1139), .b(t_1136), .c(t_1133), .d(s_80_24), .cin(t_2223), .o(t_2232), .co(t_2233), .cout(t_2234));
compressor_4_2 u2_786(.a(t_1151), .b(t_1148), .c(t_1145), .d(t_1142), .cin(t_2226), .o(t_2235), .co(t_2236), .cout(t_2237));
compressor_4_2 u2_787(.a(t_1161), .b(t_1158), .c(t_1155), .d(t_1152), .cin(t_2229), .o(t_2238), .co(t_2239), .cout(t_2240));
half_adder u0_788(.a(t_1167), .b(t_1164), .o(t_2241), .cout(t_2242));
compressor_4_2 u2_789(.a(t_1159), .b(t_1156), .c(t_1153), .d(s_81_24), .cin(t_2234), .o(t_2243), .co(t_2244), .cout(t_2245));
compressor_4_2 u2_790(.a(t_1170), .b(t_1168), .c(t_1165), .d(t_1162), .cin(t_2237), .o(t_2246), .co(t_2247), .cout(t_2248));
compressor_4_2 u2_791(.a(t_1182), .b(t_1179), .c(t_1176), .d(t_1173), .cin(t_2240), .o(t_2249), .co(t_2250), .cout(t_2251));
compressor_4_2 u2_792(.a(t_1180), .b(t_1177), .c(t_1174), .d(t_1171), .cin(t_2245), .o(t_2252), .co(t_2253), .cout(t_2254));
compressor_4_2 u2_793(.a(t_1191), .b(t_1188), .c(t_1186), .d(t_1183), .cin(t_2248), .o(t_2255), .co(t_2256), .cout(t_2257));
compressor_4_2 u2_794(.a(t_1203), .b(t_1200), .c(t_1197), .d(t_1194), .cin(t_2251), .o(t_2258), .co(t_2259), .cout(t_2260));
compressor_4_2 u2_795(.a(t_1198), .b(t_1195), .c(t_1192), .d(t_1189), .cin(t_2254), .o(t_2261), .co(t_2262), .cout(t_2263));
compressor_4_2 u2_796(.a(t_1209), .b(t_1206), .c(t_1204), .d(t_1201), .cin(t_2257), .o(t_2264), .co(t_2265), .cout(t_2266));
compressor_4_2 u2_797(.a(t_1221), .b(t_1218), .c(t_1215), .d(t_1212), .cin(t_2260), .o(t_2267), .co(t_2268), .cout(t_2269));
compressor_4_2 u2_798(.a(t_1213), .b(t_1210), .c(t_1207), .d(s_84_22), .cin(t_2263), .o(t_2270), .co(t_2271), .cout(t_2272));
compressor_4_2 u2_799(.a(t_1224), .b(t_1222), .c(t_1219), .d(t_1216), .cin(t_2266), .o(t_2273), .co(t_2274), .cout(t_2275));
compressor_4_2 u2_800(.a(t_1236), .b(t_1233), .c(t_1230), .d(t_1227), .cin(t_2269), .o(t_2276), .co(t_2277), .cout(t_2278));
compressor_4_2 u2_801(.a(t_1234), .b(t_1231), .c(t_1228), .d(t_1225), .cin(t_2272), .o(t_2279), .co(t_2280), .cout(t_2281));
compressor_4_2 u2_802(.a(t_1244), .b(t_1241), .c(t_1240), .d(t_1237), .cin(t_2275), .o(t_2282), .co(t_2283), .cout(t_2284));
compressor_4_2 u2_803(.a(t_1256), .b(t_1253), .c(t_1250), .d(t_1247), .cin(t_2278), .o(t_2285), .co(t_2286), .cout(t_2287));
compressor_4_2 u2_804(.a(t_1251), .b(t_1248), .c(t_1245), .d(t_1242), .cin(t_2281), .o(t_2288), .co(t_2289), .cout(t_2290));
compressor_4_2 u2_805(.a(t_1261), .b(t_1258), .c(t_1257), .d(t_1254), .cin(t_2284), .o(t_2291), .co(t_2292), .cout(t_2293));
compressor_4_2 u2_806(.a(t_1273), .b(t_1270), .c(t_1267), .d(t_1264), .cin(t_2287), .o(t_2294), .co(t_2295), .cout(t_2296));
compressor_4_2 u2_807(.a(t_1268), .b(t_1265), .c(t_1262), .d(t_1259), .cin(t_2290), .o(t_2297), .co(t_2298), .cout(t_2299));
compressor_4_2 u2_808(.a(t_1278), .b(t_1275), .c(t_1274), .d(t_1271), .cin(t_2293), .o(t_2300), .co(t_2301), .cout(t_2302));
compressor_4_2 u2_809(.a(t_1290), .b(t_1287), .c(t_1284), .d(t_1281), .cin(t_2296), .o(t_2303), .co(t_2304), .cout(t_2305));
compressor_4_2 u2_810(.a(t_1282), .b(t_1279), .c(t_1276), .d(s_88_20), .cin(t_2299), .o(t_2306), .co(t_2307), .cout(t_2308));
compressor_4_2 u2_811(.a(t_1292), .b(t_1291), .c(t_1288), .d(t_1285), .cin(t_2302), .o(t_2309), .co(t_2310), .cout(t_2311));
compressor_4_2 u2_812(.a(t_1304), .b(t_1301), .c(t_1298), .d(t_1295), .cin(t_2305), .o(t_2312), .co(t_2313), .cout(t_2314));
compressor_4_2 u2_813(.a(t_1299), .b(t_1296), .c(t_1293), .d(s_89_20), .cin(t_2308), .o(t_2315), .co(t_2316), .cout(t_2317));
compressor_4_2 u2_814(.a(t_1310), .b(t_1307), .c(t_1305), .d(t_1302), .cin(t_2311), .o(t_2318), .co(t_2319), .cout(t_2320));
compressor_3_2 u1_815(.a(t_1316), .b(t_1313), .cin(t_2314), .o(t_2321), .cout(t_2322));
compressor_4_2 u2_816(.a(t_1317), .b(t_1314), .c(t_1311), .d(t_1308), .cin(t_2317), .o(t_2323), .co(t_2324), .cout(t_2325));
compressor_4_2 u2_817(.a(t_1328), .b(t_1325), .c(t_1322), .d(t_1320), .cin(t_2320), .o(t_2326), .co(t_2327), .cout(t_2328));
half_adder u0_818(.a(t_1334), .b(t_1331), .o(t_2329), .cout(t_2330));
compressor_4_2 u2_819(.a(t_1332), .b(t_1329), .c(t_1326), .d(t_1323), .cin(t_2325), .o(t_2331), .co(t_2332), .cout(t_2333));
compressor_4_2 u2_820(.a(t_1343), .b(t_1340), .c(t_1337), .d(t_1335), .cin(t_2328), .o(t_2334), .co(t_2335), .cout(t_2336));
half_adder u0_821(.a(t_1349), .b(t_1346), .o(t_2337), .cout(t_2338));
compressor_4_2 u2_822(.a(t_1344), .b(t_1341), .c(t_1338), .d(s_92_18), .cin(t_2333), .o(t_2339), .co(t_2340), .cout(t_2341));
compressor_4_2 u2_823(.a(t_1355), .b(t_1352), .c(t_1350), .d(t_1347), .cin(t_2336), .o(t_2342), .co(t_2343), .cout(t_2344));
compressor_3_2 u1_824(.a(t_1364), .b(t_1361), .cin(t_1358), .o(t_2345), .cout(t_2346));
compressor_4_2 u2_825(.a(t_1362), .b(t_1359), .c(t_1356), .d(t_1353), .cin(t_2341), .o(t_2347), .co(t_2348), .cout(t_2349));
compressor_4_2 u2_826(.a(t_1372), .b(t_1369), .c(t_1366), .d(t_1365), .cin(t_2344), .o(t_2350), .co(t_2351), .cout(t_2352));
half_adder u0_827(.a(t_1378), .b(t_1375), .o(t_2353), .cout(t_2354));
compressor_4_2 u2_828(.a(t_1376), .b(t_1373), .c(t_1370), .d(t_1367), .cin(t_2349), .o(t_2355), .co(t_2356), .cout(t_2357));
compressor_4_2 u2_829(.a(t_1386), .b(t_1383), .c(t_1380), .d(t_1379), .cin(t_2352), .o(t_2358), .co(t_2359), .cout(t_2360));
half_adder u0_830(.a(t_1392), .b(t_1389), .o(t_2361), .cout(t_2362));
compressor_4_2 u2_831(.a(t_1390), .b(t_1387), .c(t_1384), .d(t_1381), .cin(t_2357), .o(t_2363), .co(t_2364), .cout(t_2365));
compressor_4_2 u2_832(.a(t_1400), .b(t_1397), .c(t_1394), .d(t_1393), .cin(t_2360), .o(t_2366), .co(t_2367), .cout(t_2368));
half_adder u0_833(.a(t_1406), .b(t_1403), .o(t_2369), .cout(t_2370));
compressor_4_2 u2_834(.a(t_1401), .b(t_1398), .c(t_1395), .d(s_96_16), .cin(t_2365), .o(t_2371), .co(t_2372), .cout(t_2373));
compressor_4_2 u2_835(.a(t_1411), .b(t_1408), .c(t_1407), .d(t_1404), .cin(t_2368), .o(t_2374), .co(t_2375), .cout(t_2376));
half_adder u0_836(.a(t_1417), .b(t_1414), .o(t_2377), .cout(t_2378));
compressor_4_2 u2_837(.a(t_1415), .b(t_1412), .c(t_1409), .d(s_97_16), .cin(t_2373), .o(t_2379), .co(t_2380), .cout(t_2381));
compressor_4_2 u2_838(.a(t_1426), .b(t_1423), .c(t_1420), .d(t_1418), .cin(t_2376), .o(t_2382), .co(t_2383), .cout(t_2384));
compressor_4_2 u2_839(.a(t_1430), .b(t_1427), .c(t_1424), .d(t_1421), .cin(t_2381), .o(t_2385), .co(t_2386), .cout(t_2387));
compressor_4_2 u2_840(.a(t_1441), .b(t_1438), .c(t_1435), .d(t_1432), .cin(t_2384), .o(t_2388), .co(t_2389), .cout(t_2390));
compressor_4_2 u2_841(.a(t_1442), .b(t_1439), .c(t_1436), .d(t_1433), .cin(t_2387), .o(t_2391), .co(t_2392), .cout(t_2393));
compressor_4_2 u2_842(.a(t_1453), .b(t_1450), .c(t_1447), .d(t_1444), .cin(t_2390), .o(t_2394), .co(t_2395), .cout(t_2396));
compressor_4_2 u2_843(.a(t_1451), .b(t_1448), .c(t_1445), .d(s_100_14), .cin(t_2393), .o(t_2397), .co(t_2398), .cout(t_2399));
compressor_4_2 u2_844(.a(t_1462), .b(t_1459), .c(t_1456), .d(t_1454), .cin(t_2396), .o(t_2400), .co(t_2401), .cout(t_2402));
compressor_4_2 u2_845(.a(t_1466), .b(t_1463), .c(t_1460), .d(t_1457), .cin(t_2399), .o(t_2403), .co(t_2404), .cout(t_2405));
compressor_4_2 u2_846(.a(t_1476), .b(t_1473), .c(t_1470), .d(t_1467), .cin(t_2402), .o(t_2406), .co(t_2407), .cout(t_2408));
compressor_4_2 u2_847(.a(t_1477), .b(t_1474), .c(t_1471), .d(t_1468), .cin(t_2405), .o(t_2409), .co(t_2410), .cout(t_2411));
compressor_4_2 u2_848(.a(t_1487), .b(t_1484), .c(t_1481), .d(t_1478), .cin(t_2408), .o(t_2412), .co(t_2413), .cout(t_2414));
compressor_4_2 u2_849(.a(t_1488), .b(t_1485), .c(t_1482), .d(t_1479), .cin(t_2411), .o(t_2415), .co(t_2416), .cout(t_2417));
compressor_4_2 u2_850(.a(t_1498), .b(t_1495), .c(t_1492), .d(t_1489), .cin(t_2414), .o(t_2418), .co(t_2419), .cout(t_2420));
compressor_4_2 u2_851(.a(t_1496), .b(t_1493), .c(t_1490), .d(s_104_12), .cin(t_2417), .o(t_2421), .co(t_2422), .cout(t_2423));
compressor_4_2 u2_852(.a(t_1506), .b(t_1503), .c(t_1500), .d(t_1499), .cin(t_2420), .o(t_2424), .co(t_2425), .cout(t_2426));
compressor_4_2 u2_853(.a(t_1507), .b(t_1504), .c(t_1501), .d(s_105_12), .cin(t_2423), .o(t_2427), .co(t_2428), .cout(t_2429));
compressor_3_2 u1_854(.a(t_1512), .b(t_1509), .cin(t_2426), .o(t_2430), .cout(t_2431));
compressor_4_2 u2_855(.a(t_1518), .b(t_1516), .c(t_1513), .d(t_1510), .cin(t_2429), .o(t_2432), .co(t_2433), .cout(t_2434));
half_adder u0_856(.a(t_1524), .b(t_1521), .o(t_2435), .cout(t_2436));
compressor_4_2 u2_857(.a(t_1527), .b(t_1525), .c(t_1522), .d(t_1519), .cin(t_2434), .o(t_2437), .co(t_2438), .cout(t_2439));
half_adder u0_858(.a(t_1533), .b(t_1530), .o(t_2440), .cout(t_2441));
compressor_4_2 u2_859(.a(t_1534), .b(t_1531), .c(t_1528), .d(s_108_10), .cin(t_2439), .o(t_2442), .co(t_2443), .cout(t_2444));
compressor_3_2 u1_860(.a(t_1542), .b(t_1539), .cin(t_1536), .o(t_2445), .cout(t_2446));
compressor_4_2 u2_861(.a(t_1544), .b(t_1543), .c(t_1540), .d(t_1537), .cin(t_2444), .o(t_2447), .co(t_2448), .cout(t_2449));
half_adder u0_862(.a(t_1550), .b(t_1547), .o(t_2450), .cout(t_2451));
compressor_4_2 u2_863(.a(t_1552), .b(t_1551), .c(t_1548), .d(t_1545), .cin(t_2449), .o(t_2452), .co(t_2453), .cout(t_2454));
half_adder u0_864(.a(t_1558), .b(t_1555), .o(t_2455), .cout(t_2456));
compressor_4_2 u2_865(.a(t_1560), .b(t_1559), .c(t_1556), .d(t_1553), .cin(t_2454), .o(t_2457), .co(t_2458), .cout(t_2459));
half_adder u0_866(.a(t_1566), .b(t_1563), .o(t_2460), .cout(t_2461));
compressor_4_2 u2_867(.a(t_1567), .b(t_1564), .c(t_1561), .d(s_112_8), .cin(t_2459), .o(t_2462), .co(t_2463), .cout(t_2464));
half_adder u0_868(.a(t_1571), .b(t_1568), .o(t_2465), .cout(t_2466));
compressor_4_2 u2_869(.a(t_1574), .b(t_1572), .c(t_1569), .d(s_113_8), .cin(t_2464), .o(t_2467), .co(t_2468), .cout(t_2469));
compressor_4_2 u2_870(.a(t_1583), .b(t_1580), .c(t_1578), .d(t_1575), .cin(t_2469), .o(t_2470), .co(t_2471), .cout(t_2472));
compressor_4_2 u2_871(.a(t_1589), .b(t_1586), .c(t_1584), .d(t_1581), .cin(t_2472), .o(t_2473), .co(t_2474), .cout(t_2475));
compressor_4_2 u2_872(.a(t_1592), .b(t_1590), .c(t_1587), .d(s_116_6), .cin(t_2475), .o(t_2476), .co(t_2477), .cout(t_2478));
compressor_4_2 u2_873(.a(t_1600), .b(t_1597), .c(t_1596), .d(t_1593), .cin(t_2478), .o(t_2479), .co(t_2480), .cout(t_2481));
compressor_4_2 u2_874(.a(t_1605), .b(t_1602), .c(t_1601), .d(t_1598), .cin(t_2481), .o(t_2482), .co(t_2483), .cout(t_2484));
compressor_4_2 u2_875(.a(t_1610), .b(t_1607), .c(t_1606), .d(t_1603), .cin(t_2484), .o(t_2485), .co(t_2486), .cout(t_2487));
compressor_4_2 u2_876(.a(t_1612), .b(t_1611), .c(t_1608), .d(s_120_4), .cin(t_2487), .o(t_2488), .co(t_2489), .cout(t_2490));
compressor_3_2 u1_877(.a(t_1613), .b(s_121_4), .cin(t_2490), .o(t_2491), .cout(t_2492));
half_adder u0_878(.a(t_1618), .b(t_1616), .o(t_2493), .cout(t_2494));
half_adder u0_879(.a(t_1621), .b(t_1619), .o(t_2495), .cout(t_2496));
compressor_3_2 u1_880(.a(t_1624), .b(t_1622), .cin(s_124_2), .o(t_2497), .cout(t_2498));
half_adder u0_881(.a(t_1626), .b(t_1625), .o(t_2499), .cout(t_2500));
half_adder u0_882(.a(t_1628), .b(t_1627), .o(t_2501), .cout(t_2502));
half_adder u0_883(.a(t_1630), .b(t_1629), .o(t_2503), .cout());

/* u0_884 Output nets */
wire t_2504,   t_2505;
/* u0_885 Output nets */
wire t_2506,   t_2507;
/* u0_886 Output nets */
wire t_2508,   t_2509;
/* u0_887 Output nets */
wire t_2510,   t_2511;
/* u0_888 Output nets */
wire t_2512,   t_2513;
/* u0_889 Output nets */
wire t_2514,   t_2515;
/* u1_890 Output nets */
wire t_2516,   t_2517;
/* u0_891 Output nets */
wire t_2518,   t_2519;
/* u1_892 Output nets */
wire t_2520,   t_2521;
/* u0_893 Output nets */
wire t_2522,   t_2523;
/* u0_894 Output nets */
wire t_2524,   t_2525;
/* u0_895 Output nets */
wire t_2526,   t_2527;
/* u0_896 Output nets */
wire t_2528,   t_2529;
/* u1_897 Output nets */
wire t_2530,   t_2531;
/* u1_898 Output nets */
wire t_2532,   t_2533;
/* u1_899 Output nets */
wire t_2534,   t_2535;
/* u1_900 Output nets */
wire t_2536,   t_2537;
/* u1_901 Output nets */
wire t_2538,   t_2539;
/* u1_902 Output nets */
wire t_2540,   t_2541;
/* u1_903 Output nets */
wire t_2542,   t_2543;
/* u1_904 Output nets */
wire t_2544,   t_2545;
/* u1_905 Output nets */
wire t_2546,   t_2547;
/* u2_906 Output nets */
wire t_2548,   t_2549,   t_2550;
/* u2_907 Output nets */
wire t_2551,   t_2552,   t_2553;
/* u2_908 Output nets */
wire t_2554,   t_2555,   t_2556;
/* u2_909 Output nets */
wire t_2557,   t_2558,   t_2559;
/* u2_910 Output nets */
wire t_2560,   t_2561,   t_2562;
/* u2_911 Output nets */
wire t_2563,   t_2564,   t_2565;
/* u2_912 Output nets */
wire t_2566,   t_2567,   t_2568;
/* u2_913 Output nets */
wire t_2569,   t_2570,   t_2571;
/* u2_914 Output nets */
wire t_2572,   t_2573,   t_2574;
/* u2_915 Output nets */
wire t_2575,   t_2576,   t_2577;
/* u0_916 Output nets */
wire t_2578,   t_2579;
/* u2_917 Output nets */
wire t_2580,   t_2581,   t_2582;
/* u2_918 Output nets */
wire t_2583,   t_2584,   t_2585;
/* u0_919 Output nets */
wire t_2586,   t_2587;
/* u2_920 Output nets */
wire t_2588,   t_2589,   t_2590;
/* u0_921 Output nets */
wire t_2591,   t_2592;
/* u2_922 Output nets */
wire t_2593,   t_2594,   t_2595;
/* u0_923 Output nets */
wire t_2596,   t_2597;
/* u2_924 Output nets */
wire t_2598,   t_2599,   t_2600;
/* u0_925 Output nets */
wire t_2601,   t_2602;
/* u2_926 Output nets */
wire t_2603,   t_2604,   t_2605;
/* u0_927 Output nets */
wire t_2606,   t_2607;
/* u2_928 Output nets */
wire t_2608,   t_2609,   t_2610;
/* u1_929 Output nets */
wire t_2611,   t_2612;
/* u2_930 Output nets */
wire t_2613,   t_2614,   t_2615;
/* u0_931 Output nets */
wire t_2616,   t_2617;
/* u2_932 Output nets */
wire t_2618,   t_2619,   t_2620;
/* u1_933 Output nets */
wire t_2621,   t_2622;
/* u2_934 Output nets */
wire t_2623,   t_2624,   t_2625;
/* u0_935 Output nets */
wire t_2626,   t_2627;
/* u2_936 Output nets */
wire t_2628,   t_2629,   t_2630;
/* u0_937 Output nets */
wire t_2631,   t_2632;
/* u2_938 Output nets */
wire t_2633,   t_2634,   t_2635;
/* u0_939 Output nets */
wire t_2636,   t_2637;
/* u2_940 Output nets */
wire t_2638,   t_2639,   t_2640;
/* u0_941 Output nets */
wire t_2641,   t_2642;
/* u2_942 Output nets */
wire t_2643,   t_2644,   t_2645;
/* u1_943 Output nets */
wire t_2646,   t_2647;
/* u2_944 Output nets */
wire t_2648,   t_2649,   t_2650;
/* u1_945 Output nets */
wire t_2651,   t_2652;
/* u2_946 Output nets */
wire t_2653,   t_2654,   t_2655;
/* u1_947 Output nets */
wire t_2656,   t_2657;
/* u2_948 Output nets */
wire t_2658,   t_2659,   t_2660;
/* u1_949 Output nets */
wire t_2661,   t_2662;
/* u2_950 Output nets */
wire t_2663,   t_2664,   t_2665;
/* u1_951 Output nets */
wire t_2666,   t_2667;
/* u2_952 Output nets */
wire t_2668,   t_2669,   t_2670;
/* u1_953 Output nets */
wire t_2671,   t_2672;
/* u2_954 Output nets */
wire t_2673,   t_2674,   t_2675;
/* u1_955 Output nets */
wire t_2676,   t_2677;
/* u2_956 Output nets */
wire t_2678,   t_2679,   t_2680;
/* u1_957 Output nets */
wire t_2681,   t_2682;
/* u2_958 Output nets */
wire t_2683,   t_2684,   t_2685;
/* u1_959 Output nets */
wire t_2686,   t_2687;
/* u2_960 Output nets */
wire t_2688,   t_2689,   t_2690;
/* u2_961 Output nets */
wire t_2691,   t_2692,   t_2693;
/* u2_962 Output nets */
wire t_2694,   t_2695,   t_2696;
/* u2_963 Output nets */
wire t_2697,   t_2698,   t_2699;
/* u2_964 Output nets */
wire t_2700,   t_2701,   t_2702;
/* u2_965 Output nets */
wire t_2703,   t_2704,   t_2705;
/* u2_966 Output nets */
wire t_2706,   t_2707,   t_2708;
/* u2_967 Output nets */
wire t_2709,   t_2710,   t_2711;
/* u2_968 Output nets */
wire t_2712,   t_2713,   t_2714;
/* u2_969 Output nets */
wire t_2715,   t_2716,   t_2717;
/* u2_970 Output nets */
wire t_2718,   t_2719,   t_2720;
/* u2_971 Output nets */
wire t_2721,   t_2722,   t_2723;
/* u2_972 Output nets */
wire t_2724,   t_2725,   t_2726;
/* u2_973 Output nets */
wire t_2727,   t_2728,   t_2729;
/* u2_974 Output nets */
wire t_2730,   t_2731,   t_2732;
/* u2_975 Output nets */
wire t_2733,   t_2734,   t_2735;
/* u2_976 Output nets */
wire t_2736,   t_2737,   t_2738;
/* u2_977 Output nets */
wire t_2739,   t_2740,   t_2741;
/* u2_978 Output nets */
wire t_2742,   t_2743,   t_2744;
/* u2_979 Output nets */
wire t_2745,   t_2746,   t_2747;
/* u2_980 Output nets */
wire t_2748,   t_2749,   t_2750;
/* u2_981 Output nets */
wire t_2751,   t_2752,   t_2753;
/* u2_982 Output nets */
wire t_2754,   t_2755,   t_2756;
/* u2_983 Output nets */
wire t_2757,   t_2758,   t_2759;
/* u2_984 Output nets */
wire t_2760,   t_2761,   t_2762;
/* u2_985 Output nets */
wire t_2763,   t_2764,   t_2765;
/* u2_986 Output nets */
wire t_2766,   t_2767,   t_2768;
/* u2_987 Output nets */
wire t_2769,   t_2770,   t_2771;
/* u2_988 Output nets */
wire t_2772,   t_2773,   t_2774;
/* u2_989 Output nets */
wire t_2775,   t_2776,   t_2777;
/* u2_990 Output nets */
wire t_2778,   t_2779,   t_2780;
/* u2_991 Output nets */
wire t_2781,   t_2782,   t_2783;
/* u2_992 Output nets */
wire t_2784,   t_2785,   t_2786;
/* u2_993 Output nets */
wire t_2787,   t_2788,   t_2789;
/* u2_994 Output nets */
wire t_2790,   t_2791,   t_2792;
/* u2_995 Output nets */
wire t_2793,   t_2794,   t_2795;
/* u2_996 Output nets */
wire t_2796,   t_2797,   t_2798;
/* u2_997 Output nets */
wire t_2799,   t_2800,   t_2801;
/* u2_998 Output nets */
wire t_2802,   t_2803,   t_2804;
/* u2_999 Output nets */
wire t_2805,   t_2806,   t_2807;
/* u2_1000 Output nets */
wire t_2808,   t_2809,   t_2810;
/* u2_1001 Output nets */
wire t_2811,   t_2812,   t_2813;
/* u2_1002 Output nets */
wire t_2814,   t_2815,   t_2816;
/* u2_1003 Output nets */
wire t_2817,   t_2818,   t_2819;
/* u2_1004 Output nets */
wire t_2820,   t_2821,   t_2822;
/* u2_1005 Output nets */
wire t_2823,   t_2824,   t_2825;
/* u2_1006 Output nets */
wire t_2826,   t_2827,   t_2828;
/* u2_1007 Output nets */
wire t_2829,   t_2830,   t_2831;
/* u2_1008 Output nets */
wire t_2832,   t_2833,   t_2834;
/* u2_1009 Output nets */
wire t_2835,   t_2836,   t_2837;
/* u2_1010 Output nets */
wire t_2838,   t_2839,   t_2840;
/* u1_1011 Output nets */
wire t_2841,   t_2842;
/* u2_1012 Output nets */
wire t_2843,   t_2844,   t_2845;
/* u0_1013 Output nets */
wire t_2846,   t_2847;
/* u2_1014 Output nets */
wire t_2848,   t_2849,   t_2850;
/* u1_1015 Output nets */
wire t_2851,   t_2852;
/* u2_1016 Output nets */
wire t_2853,   t_2854,   t_2855;
/* u0_1017 Output nets */
wire t_2856,   t_2857;
/* u2_1018 Output nets */
wire t_2858,   t_2859,   t_2860;
/* u0_1019 Output nets */
wire t_2861,   t_2862;
/* u2_1020 Output nets */
wire t_2863,   t_2864,   t_2865;
/* u0_1021 Output nets */
wire t_2866,   t_2867;
/* u2_1022 Output nets */
wire t_2868,   t_2869,   t_2870;
/* u0_1023 Output nets */
wire t_2871,   t_2872;
/* u2_1024 Output nets */
wire t_2873,   t_2874,   t_2875;
/* u1_1025 Output nets */
wire t_2876,   t_2877;
/* u2_1026 Output nets */
wire t_2878,   t_2879,   t_2880;
/* u0_1027 Output nets */
wire t_2881,   t_2882;
/* u2_1028 Output nets */
wire t_2883,   t_2884,   t_2885;
/* u0_1029 Output nets */
wire t_2886,   t_2887;
/* u2_1030 Output nets */
wire t_2888,   t_2889,   t_2890;
/* u0_1031 Output nets */
wire t_2891,   t_2892;
/* u2_1032 Output nets */
wire t_2893,   t_2894,   t_2895;
/* u0_1033 Output nets */
wire t_2896,   t_2897;
/* u2_1034 Output nets */
wire t_2898,   t_2899,   t_2900;
/* u0_1035 Output nets */
wire t_2901,   t_2902;
/* u2_1036 Output nets */
wire t_2903,   t_2904,   t_2905;
/* u0_1037 Output nets */
wire t_2906,   t_2907;
/* u2_1038 Output nets */
wire t_2908,   t_2909,   t_2910;
/* u0_1039 Output nets */
wire t_2911,   t_2912;
/* u2_1040 Output nets */
wire t_2913,   t_2914,   t_2915;
/* u0_1041 Output nets */
wire t_2916,   t_2917;
/* u2_1042 Output nets */
wire t_2918,   t_2919,   t_2920;
/* u2_1043 Output nets */
wire t_2921,   t_2922,   t_2923;
/* u2_1044 Output nets */
wire t_2924,   t_2925,   t_2926;
/* u2_1045 Output nets */
wire t_2927,   t_2928,   t_2929;
/* u2_1046 Output nets */
wire t_2930,   t_2931,   t_2932;
/* u2_1047 Output nets */
wire t_2933,   t_2934,   t_2935;
/* u2_1048 Output nets */
wire t_2936,   t_2937,   t_2938;
/* u2_1049 Output nets */
wire t_2939,   t_2940,   t_2941;
/* u2_1050 Output nets */
wire t_2942,   t_2943,   t_2944;
/* u2_1051 Output nets */
wire t_2945,   t_2946,   t_2947;
/* u2_1052 Output nets */
wire t_2948,   t_2949,   t_2950;
/* u2_1053 Output nets */
wire t_2951,   t_2952,   t_2953;
/* u2_1054 Output nets */
wire t_2954,   t_2955,   t_2956;
/* u2_1055 Output nets */
wire t_2957,   t_2958,   t_2959;
/* u2_1056 Output nets */
wire t_2960,   t_2961,   t_2962;
/* u2_1057 Output nets */
wire t_2963,   t_2964,   t_2965;
/* u1_1058 Output nets */
wire t_2966,   t_2967;
/* u0_1059 Output nets */
wire t_2968,   t_2969;
/* u1_1060 Output nets */
wire t_2970,   t_2971;
/* u0_1061 Output nets */
wire t_2972,   t_2973;
/* u0_1062 Output nets */
wire t_2974,   t_2975;
/* u0_1063 Output nets */
wire t_2976,   t_2977;
/* u0_1064 Output nets */
wire t_2978,   t_2979;
/* u1_1065 Output nets */
wire t_2980,   t_2981;
/* u0_1066 Output nets */
wire t_2982,   t_2983;
/* u0_1067 Output nets */
wire t_2984,   t_2985;
/* u0_1068 Output nets */
wire t_2986,   t_2987;
/* u0_1069 Output nets */
wire t_2988,   t_2989;
/* u0_1070 Output nets */
wire t_2990,   t_2991;
/* u0_1071 Output nets */
wire t_2992;

/* compress stage 3 */
half_adder u0_884(.a(t_1632), .b(t_2), .o(t_2504), .cout(t_2505));
half_adder u0_885(.a(t_1635), .b(t_1634), .o(t_2506), .cout(t_2507));
half_adder u0_886(.a(t_1637), .b(t_1636), .o(t_2508), .cout(t_2509));
half_adder u0_887(.a(t_1639), .b(t_1638), .o(t_2510), .cout(t_2511));
half_adder u0_888(.a(t_1641), .b(t_1640), .o(t_2512), .cout(t_2513));
half_adder u0_889(.a(t_1643), .b(t_1642), .o(t_2514), .cout(t_2515));
compressor_3_2 u1_890(.a(t_1645), .b(t_1644), .cin(t_21), .o(t_2516), .cout(t_2517));
half_adder u0_891(.a(t_1647), .b(t_1646), .o(t_2518), .cout(t_2519));
compressor_3_2 u1_892(.a(t_1649), .b(t_1648), .cin(t_32), .o(t_2520), .cout(t_2521));
half_adder u0_893(.a(t_1651), .b(t_1650), .o(t_2522), .cout(t_2523));
half_adder u0_894(.a(t_1654), .b(t_1652), .o(t_2524), .cout(t_2525));
half_adder u0_895(.a(t_1657), .b(t_1655), .o(t_2526), .cout(t_2527));
half_adder u0_896(.a(t_1660), .b(t_1658), .o(t_2528), .cout(t_2529));
compressor_3_2 u1_897(.a(t_1663), .b(t_1661), .cin(t_62), .o(t_2530), .cout(t_2531));
compressor_3_2 u1_898(.a(t_1669), .b(t_1666), .cin(t_1664), .o(t_2532), .cout(t_2533));
compressor_3_2 u1_899(.a(t_1670), .b(t_1667), .cin(t_76), .o(t_2534), .cout(t_2535));
compressor_3_2 u1_900(.a(t_1677), .b(t_1674), .cin(t_1672), .o(t_2536), .cout(t_2537));
compressor_3_2 u1_901(.a(t_1679), .b(t_1678), .cin(t_1675), .o(t_2538), .cout(t_2539));
compressor_3_2 u1_902(.a(t_1684), .b(t_1683), .cin(t_1680), .o(t_2540), .cout(t_2541));
compressor_3_2 u1_903(.a(t_1689), .b(t_1688), .cin(t_1685), .o(t_2542), .cout(t_2543));
compressor_3_2 u1_904(.a(t_1694), .b(t_1693), .cin(t_1690), .o(t_2544), .cout(t_2545));
compressor_3_2 u1_905(.a(t_1699), .b(t_1698), .cin(t_1695), .o(t_2546), .cout(t_2547));
compressor_4_2 u2_906(.a(t_1707), .b(t_1704), .c(t_1703), .d(t_1700), .cin(t_137), .o(t_2548), .co(t_2549), .cout(t_2550));
compressor_4_2 u2_907(.a(t_1712), .b(t_1709), .c(t_1708), .d(t_1705), .cin(t_2550), .o(t_2551), .co(t_2552), .cout(t_2553));
compressor_4_2 u2_908(.a(t_1714), .b(t_1713), .c(t_1710), .d(t_160), .cin(t_2553), .o(t_2554), .co(t_2555), .cout(t_2556));
compressor_4_2 u2_909(.a(t_1722), .b(t_1719), .c(t_1718), .d(t_1715), .cin(t_2556), .o(t_2557), .co(t_2558), .cout(t_2559));
compressor_4_2 u2_910(.a(t_1728), .b(t_1725), .c(t_1723), .d(t_1720), .cin(t_2559), .o(t_2560), .co(t_2561), .cout(t_2562));
compressor_4_2 u2_911(.a(t_1734), .b(t_1731), .c(t_1729), .d(t_1726), .cin(t_2562), .o(t_2563), .co(t_2564), .cout(t_2565));
compressor_4_2 u2_912(.a(t_1740), .b(t_1737), .c(t_1735), .d(t_1732), .cin(t_2565), .o(t_2566), .co(t_2567), .cout(t_2568));
compressor_4_2 u2_913(.a(t_1743), .b(t_1741), .c(t_1738), .d(t_220), .cin(t_2568), .o(t_2569), .co(t_2570), .cout(t_2571));
compressor_4_2 u2_914(.a(t_1752), .b(t_1749), .c(t_1747), .d(t_1744), .cin(t_2571), .o(t_2572), .co(t_2573), .cout(t_2574));
compressor_4_2 u2_915(.a(t_1756), .b(t_1753), .c(t_1750), .d(t_246), .cin(t_2574), .o(t_2575), .co(t_2576), .cout(t_2577));
half_adder u0_916(.a(t_1760), .b(t_1757), .o(t_2578), .cout(t_2579));
compressor_4_2 u2_917(.a(t_1766), .b(t_1763), .c(t_1761), .d(t_1758), .cin(t_2577), .o(t_2580), .co(t_2581), .cout(t_2582));
compressor_4_2 u2_918(.a(t_1771), .b(t_1770), .c(t_1767), .d(t_1764), .cin(t_2582), .o(t_2583), .co(t_2584), .cout(t_2585));
half_adder u0_919(.a(t_1777), .b(t_1774), .o(t_2586), .cout(t_2587));
compressor_4_2 u2_920(.a(t_1779), .b(t_1778), .c(t_1775), .d(t_1772), .cin(t_2585), .o(t_2588), .co(t_2589), .cout(t_2590));
half_adder u0_921(.a(t_1785), .b(t_1782), .o(t_2591), .cout(t_2592));
compressor_4_2 u2_922(.a(t_1787), .b(t_1786), .c(t_1783), .d(t_1780), .cin(t_2590), .o(t_2593), .co(t_2594), .cout(t_2595));
half_adder u0_923(.a(t_1793), .b(t_1790), .o(t_2596), .cout(t_2597));
compressor_4_2 u2_924(.a(t_1795), .b(t_1794), .c(t_1791), .d(t_1788), .cin(t_2595), .o(t_2598), .co(t_2599), .cout(t_2600));
half_adder u0_925(.a(t_1801), .b(t_1798), .o(t_2601), .cout(t_2602));
compressor_4_2 u2_926(.a(t_1803), .b(t_1802), .c(t_1799), .d(t_1796), .cin(t_2600), .o(t_2603), .co(t_2604), .cout(t_2605));
half_adder u0_927(.a(t_1809), .b(t_1806), .o(t_2606), .cout(t_2607));
compressor_4_2 u2_928(.a(t_1810), .b(t_1807), .c(t_1804), .d(t_349), .cin(t_2605), .o(t_2608), .co(t_2609), .cout(t_2610));
compressor_3_2 u1_929(.a(t_1817), .b(t_1814), .cin(t_1811), .o(t_2611), .cout(t_2612));
compressor_4_2 u2_930(.a(t_1819), .b(t_1818), .c(t_1815), .d(t_1812), .cin(t_2610), .o(t_2613), .co(t_2614), .cout(t_2615));
half_adder u0_931(.a(t_1825), .b(t_1822), .o(t_2616), .cout(t_2617));
compressor_4_2 u2_932(.a(t_1826), .b(t_1823), .c(t_1820), .d(t_384), .cin(t_2615), .o(t_2618), .co(t_2619), .cout(t_2620));
compressor_3_2 u1_933(.a(t_1833), .b(t_1830), .cin(t_1827), .o(t_2621), .cout(t_2622));
compressor_4_2 u2_934(.a(t_1835), .b(t_1834), .c(t_1831), .d(t_1828), .cin(t_2620), .o(t_2623), .co(t_2624), .cout(t_2625));
half_adder u0_935(.a(t_1841), .b(t_1838), .o(t_2626), .cout(t_2627));
compressor_4_2 u2_936(.a(t_1844), .b(t_1842), .c(t_1839), .d(t_1836), .cin(t_2625), .o(t_2628), .co(t_2629), .cout(t_2630));
half_adder u0_937(.a(t_1850), .b(t_1847), .o(t_2631), .cout(t_2632));
compressor_4_2 u2_938(.a(t_1853), .b(t_1851), .c(t_1848), .d(t_1845), .cin(t_2630), .o(t_2633), .co(t_2634), .cout(t_2635));
half_adder u0_939(.a(t_1859), .b(t_1856), .o(t_2636), .cout(t_2637));
compressor_4_2 u2_940(.a(t_1862), .b(t_1860), .c(t_1857), .d(t_1854), .cin(t_2635), .o(t_2638), .co(t_2639), .cout(t_2640));
half_adder u0_941(.a(t_1868), .b(t_1865), .o(t_2641), .cout(t_2642));
compressor_4_2 u2_942(.a(t_1869), .b(t_1866), .c(t_1863), .d(t_474), .cin(t_2640), .o(t_2643), .co(t_2644), .cout(t_2645));
compressor_3_2 u1_943(.a(t_1877), .b(t_1874), .cin(t_1871), .o(t_2646), .cout(t_2647));
compressor_4_2 u2_944(.a(t_1880), .b(t_1878), .c(t_1875), .d(t_1872), .cin(t_2645), .o(t_2648), .co(t_2649), .cout(t_2650));
compressor_3_2 u1_945(.a(t_1889), .b(t_1886), .cin(t_1883), .o(t_2651), .cout(t_2652));
compressor_4_2 u2_946(.a(t_1887), .b(t_1884), .c(t_1881), .d(t_512), .cin(t_2650), .o(t_2653), .co(t_2654), .cout(t_2655));
compressor_3_2 u1_947(.a(t_1894), .b(t_1891), .cin(t_1890), .o(t_2656), .cout(t_2657));
compressor_4_2 u2_948(.a(t_1900), .b(t_1898), .c(t_1895), .d(t_1892), .cin(t_2655), .o(t_2658), .co(t_2659), .cout(t_2660));
compressor_3_2 u1_949(.a(t_1909), .b(t_1906), .cin(t_1903), .o(t_2661), .cout(t_2662));
compressor_4_2 u2_950(.a(t_1910), .b(t_1907), .c(t_1904), .d(t_1901), .cin(t_2660), .o(t_2663), .co(t_2664), .cout(t_2665));
compressor_3_2 u1_951(.a(t_1917), .b(t_1914), .cin(t_1911), .o(t_2666), .cout(t_2667));
compressor_4_2 u2_952(.a(t_1921), .b(t_1918), .c(t_1915), .d(t_1912), .cin(t_2665), .o(t_2668), .co(t_2669), .cout(t_2670));
compressor_3_2 u1_953(.a(t_1928), .b(t_1925), .cin(t_1922), .o(t_2671), .cout(t_2672));
compressor_4_2 u2_954(.a(t_1932), .b(t_1929), .c(t_1926), .d(t_1923), .cin(t_2670), .o(t_2673), .co(t_2674), .cout(t_2675));
compressor_3_2 u1_955(.a(t_1939), .b(t_1936), .cin(t_1933), .o(t_2676), .cout(t_2677));
compressor_4_2 u2_956(.a(t_1943), .b(t_1940), .c(t_1937), .d(t_1934), .cin(t_2675), .o(t_2678), .co(t_2679), .cout(t_2680));
compressor_3_2 u1_957(.a(t_1950), .b(t_1947), .cin(t_1944), .o(t_2681), .cout(t_2682));
compressor_4_2 u2_958(.a(t_1954), .b(t_1951), .c(t_1948), .d(t_1945), .cin(t_2680), .o(t_2683), .co(t_2684), .cout(t_2685));
compressor_3_2 u1_959(.a(t_1961), .b(t_1958), .cin(t_1955), .o(t_2686), .cout(t_2687));
compressor_4_2 u2_960(.a(t_1962), .b(t_1959), .c(t_1956), .d(t_657), .cin(t_2685), .o(t_2688), .co(t_2689), .cout(t_2690));
compressor_4_2 u2_961(.a(t_1975), .b(t_1972), .c(t_1969), .d(t_1966), .cin(t_1965), .o(t_2691), .co(t_2692), .cout(t_2693));
compressor_4_2 u2_962(.a(t_1976), .b(t_1973), .c(t_1970), .d(t_1967), .cin(t_2690), .o(t_2694), .co(t_2695), .cout(t_2696));
compressor_4_2 u2_963(.a(t_1986), .b(t_1983), .c(t_1980), .d(t_1977), .cin(t_2693), .o(t_2697), .co(t_2698), .cout(t_2699));
compressor_4_2 u2_964(.a(t_1984), .b(t_1981), .c(t_1978), .d(t_704), .cin(t_2696), .o(t_2700), .co(t_2701), .cout(t_2702));
compressor_4_2 u2_965(.a(t_1994), .b(t_1991), .c(t_1988), .d(t_1987), .cin(t_2699), .o(t_2703), .co(t_2704), .cout(t_2705));
compressor_4_2 u2_966(.a(t_1998), .b(t_1995), .c(t_1992), .d(t_1989), .cin(t_2702), .o(t_2706), .co(t_2707), .cout(t_2708));
compressor_4_2 u2_967(.a(t_2008), .b(t_2005), .c(t_2002), .d(t_1999), .cin(t_2705), .o(t_2709), .co(t_2710), .cout(t_2711));
compressor_4_2 u2_968(.a(t_2009), .b(t_2006), .c(t_2003), .d(t_2000), .cin(t_2708), .o(t_2712), .co(t_2713), .cout(t_2714));
compressor_4_2 u2_969(.a(t_2020), .b(t_2017), .c(t_2014), .d(t_2011), .cin(t_2711), .o(t_2715), .co(t_2716), .cout(t_2717));
compressor_4_2 u2_970(.a(t_2021), .b(t_2018), .c(t_2015), .d(t_2012), .cin(t_2714), .o(t_2718), .co(t_2719), .cout(t_2720));
compressor_4_2 u2_971(.a(t_2032), .b(t_2029), .c(t_2026), .d(t_2023), .cin(t_2717), .o(t_2721), .co(t_2722), .cout(t_2723));
compressor_4_2 u2_972(.a(t_2033), .b(t_2030), .c(t_2027), .d(t_2024), .cin(t_2720), .o(t_2724), .co(t_2725), .cout(t_2726));
compressor_4_2 u2_973(.a(t_2044), .b(t_2041), .c(t_2038), .d(t_2035), .cin(t_2723), .o(t_2727), .co(t_2728), .cout(t_2729));
compressor_4_2 u2_974(.a(t_2042), .b(t_2039), .c(t_2036), .d(t_821), .cin(t_2726), .o(t_2730), .co(t_2731), .cout(t_2732));
compressor_4_2 u2_975(.a(t_2053), .b(t_2050), .c(t_2047), .d(t_2045), .cin(t_2729), .o(t_2733), .co(t_2734), .cout(t_2735));
compressor_4_2 u2_976(.a(t_2054), .b(t_2051), .c(t_2048), .d(t_845), .cin(t_2732), .o(t_2736), .co(t_2737), .cout(t_2738));
compressor_4_2 u2_977(.a(t_2065), .b(t_2062), .c(t_2059), .d(t_2057), .cin(t_2735), .o(t_2739), .co(t_2740), .cout(t_2741));
compressor_4_2 u2_978(.a(t_2069), .b(t_2066), .c(t_2063), .d(t_2060), .cin(t_2738), .o(t_2742), .co(t_2743), .cout(t_2744));
compressor_4_2 u2_979(.a(t_2080), .b(t_2077), .c(t_2074), .d(t_2071), .cin(t_2741), .o(t_2745), .co(t_2746), .cout(t_2747));
compressor_4_2 u2_980(.a(t_2081), .b(t_2078), .c(t_2075), .d(t_2072), .cin(t_2744), .o(t_2748), .co(t_2749), .cout(t_2750));
compressor_4_2 u2_981(.a(t_2092), .b(t_2089), .c(t_2086), .d(t_2083), .cin(t_2747), .o(t_2751), .co(t_2752), .cout(t_2753));
compressor_4_2 u2_982(.a(t_2090), .b(t_2087), .c(t_2084), .d(t_917), .cin(t_2750), .o(t_2754), .co(t_2755), .cout(t_2756));
compressor_4_2 u2_983(.a(t_2101), .b(t_2098), .c(t_2095), .d(t_2093), .cin(t_2753), .o(t_2757), .co(t_2758), .cout(t_2759));
compressor_4_2 u2_984(.a(t_2105), .b(t_2102), .c(t_2099), .d(t_2096), .cin(t_2756), .o(t_2760), .co(t_2761), .cout(t_2762));
compressor_4_2 u2_985(.a(t_2116), .b(t_2113), .c(t_2110), .d(t_2107), .cin(t_2759), .o(t_2763), .co(t_2764), .cout(t_2765));
compressor_4_2 u2_986(.a(t_2117), .b(t_2114), .c(t_2111), .d(t_2108), .cin(t_2762), .o(t_2766), .co(t_2767), .cout(t_2768));
compressor_4_2 u2_987(.a(t_2128), .b(t_2125), .c(t_2122), .d(t_2119), .cin(t_2765), .o(t_2769), .co(t_2770), .cout(t_2771));
compressor_4_2 u2_988(.a(t_2129), .b(t_2126), .c(t_2123), .d(t_2120), .cin(t_2768), .o(t_2772), .co(t_2773), .cout(t_2774));
compressor_4_2 u2_989(.a(t_2140), .b(t_2137), .c(t_2134), .d(t_2131), .cin(t_2771), .o(t_2775), .co(t_2776), .cout(t_2777));
compressor_4_2 u2_990(.a(t_2141), .b(t_2138), .c(t_2135), .d(t_2132), .cin(t_2774), .o(t_2778), .co(t_2779), .cout(t_2780));
compressor_4_2 u2_991(.a(t_2152), .b(t_2149), .c(t_2146), .d(t_2143), .cin(t_2777), .o(t_2781), .co(t_2782), .cout(t_2783));
compressor_4_2 u2_992(.a(t_2150), .b(t_2147), .c(t_2144), .d(t_1027), .cin(t_2780), .o(t_2784), .co(t_2785), .cout(t_2786));
compressor_4_2 u2_993(.a(t_2161), .b(t_2158), .c(t_2155), .d(t_2153), .cin(t_2783), .o(t_2787), .co(t_2788), .cout(t_2789));
compressor_4_2 u2_994(.a(t_2165), .b(t_2162), .c(t_2159), .d(t_2156), .cin(t_2786), .o(t_2790), .co(t_2791), .cout(t_2792));
compressor_4_2 u2_995(.a(t_2175), .b(t_2172), .c(t_2169), .d(t_2166), .cin(t_2789), .o(t_2793), .co(t_2794), .cout(t_2795));
compressor_4_2 u2_996(.a(t_2176), .b(t_2173), .c(t_2170), .d(t_2167), .cin(t_2792), .o(t_2796), .co(t_2797), .cout(t_2798));
compressor_4_2 u2_997(.a(t_2186), .b(t_2183), .c(t_2180), .d(t_2177), .cin(t_2795), .o(t_2799), .co(t_2800), .cout(t_2801));
compressor_4_2 u2_998(.a(t_2187), .b(t_2184), .c(t_2181), .d(t_2178), .cin(t_2798), .o(t_2802), .co(t_2803), .cout(t_2804));
compressor_4_2 u2_999(.a(t_2197), .b(t_2194), .c(t_2191), .d(t_2188), .cin(t_2801), .o(t_2805), .co(t_2806), .cout(t_2807));
compressor_4_2 u2_1000(.a(t_2198), .b(t_2195), .c(t_2192), .d(t_2189), .cin(t_2804), .o(t_2808), .co(t_2809), .cout(t_2810));
compressor_4_2 u2_1001(.a(t_2208), .b(t_2205), .c(t_2202), .d(t_2199), .cin(t_2807), .o(t_2811), .co(t_2812), .cout(t_2813));
compressor_4_2 u2_1002(.a(t_2209), .b(t_2206), .c(t_2203), .d(t_2200), .cin(t_2810), .o(t_2814), .co(t_2815), .cout(t_2816));
compressor_4_2 u2_1003(.a(t_2219), .b(t_2216), .c(t_2213), .d(t_2210), .cin(t_2813), .o(t_2817), .co(t_2818), .cout(t_2819));
compressor_4_2 u2_1004(.a(t_2220), .b(t_2217), .c(t_2214), .d(t_2211), .cin(t_2816), .o(t_2820), .co(t_2821), .cout(t_2822));
compressor_4_2 u2_1005(.a(t_2230), .b(t_2227), .c(t_2224), .d(t_2221), .cin(t_2819), .o(t_2823), .co(t_2824), .cout(t_2825));
compressor_4_2 u2_1006(.a(t_2231), .b(t_2228), .c(t_2225), .d(t_2222), .cin(t_2822), .o(t_2826), .co(t_2827), .cout(t_2828));
compressor_4_2 u2_1007(.a(t_2241), .b(t_2238), .c(t_2235), .d(t_2232), .cin(t_2825), .o(t_2829), .co(t_2830), .cout(t_2831));
compressor_4_2 u2_1008(.a(t_2239), .b(t_2236), .c(t_2233), .d(t_1185), .cin(t_2828), .o(t_2832), .co(t_2833), .cout(t_2834));
compressor_4_2 u2_1009(.a(t_2249), .b(t_2246), .c(t_2243), .d(t_2242), .cin(t_2831), .o(t_2835), .co(t_2836), .cout(t_2837));
compressor_4_2 u2_1010(.a(t_2252), .b(t_2250), .c(t_2247), .d(t_2244), .cin(t_2834), .o(t_2838), .co(t_2839), .cout(t_2840));
compressor_3_2 u1_1011(.a(t_2258), .b(t_2255), .cin(t_2837), .o(t_2841), .cout(t_2842));
compressor_4_2 u2_1012(.a(t_2261), .b(t_2259), .c(t_2256), .d(t_2253), .cin(t_2840), .o(t_2843), .co(t_2844), .cout(t_2845));
half_adder u0_1013(.a(t_2267), .b(t_2264), .o(t_2846), .cout(t_2847));
compressor_4_2 u2_1014(.a(t_2268), .b(t_2265), .c(t_2262), .d(t_1239), .cin(t_2845), .o(t_2848), .co(t_2849), .cout(t_2850));
compressor_3_2 u1_1015(.a(t_2276), .b(t_2273), .cin(t_2270), .o(t_2851), .cout(t_2852));
compressor_4_2 u2_1016(.a(t_2279), .b(t_2277), .c(t_2274), .d(t_2271), .cin(t_2850), .o(t_2853), .co(t_2854), .cout(t_2855));
half_adder u0_1017(.a(t_2285), .b(t_2282), .o(t_2856), .cout(t_2857));
compressor_4_2 u2_1018(.a(t_2288), .b(t_2286), .c(t_2283), .d(t_2280), .cin(t_2855), .o(t_2858), .co(t_2859), .cout(t_2860));
half_adder u0_1019(.a(t_2294), .b(t_2291), .o(t_2861), .cout(t_2862));
compressor_4_2 u2_1020(.a(t_2297), .b(t_2295), .c(t_2292), .d(t_2289), .cin(t_2860), .o(t_2863), .co(t_2864), .cout(t_2865));
half_adder u0_1021(.a(t_2303), .b(t_2300), .o(t_2866), .cout(t_2867));
compressor_4_2 u2_1022(.a(t_2306), .b(t_2304), .c(t_2301), .d(t_2298), .cin(t_2865), .o(t_2868), .co(t_2869), .cout(t_2870));
half_adder u0_1023(.a(t_2312), .b(t_2309), .o(t_2871), .cout(t_2872));
compressor_4_2 u2_1024(.a(t_2313), .b(t_2310), .c(t_2307), .d(t_1319), .cin(t_2870), .o(t_2873), .co(t_2874), .cout(t_2875));
compressor_3_2 u1_1025(.a(t_2321), .b(t_2318), .cin(t_2315), .o(t_2876), .cout(t_2877));
compressor_4_2 u2_1026(.a(t_2323), .b(t_2322), .c(t_2319), .d(t_2316), .cin(t_2875), .o(t_2878), .co(t_2879), .cout(t_2880));
half_adder u0_1027(.a(t_2329), .b(t_2326), .o(t_2881), .cout(t_2882));
compressor_4_2 u2_1028(.a(t_2331), .b(t_2330), .c(t_2327), .d(t_2324), .cin(t_2880), .o(t_2883), .co(t_2884), .cout(t_2885));
half_adder u0_1029(.a(t_2337), .b(t_2334), .o(t_2886), .cout(t_2887));
compressor_4_2 u2_1030(.a(t_2339), .b(t_2338), .c(t_2335), .d(t_2332), .cin(t_2885), .o(t_2888), .co(t_2889), .cout(t_2890));
half_adder u0_1031(.a(t_2345), .b(t_2342), .o(t_2891), .cout(t_2892));
compressor_4_2 u2_1032(.a(t_2347), .b(t_2346), .c(t_2343), .d(t_2340), .cin(t_2890), .o(t_2893), .co(t_2894), .cout(t_2895));
half_adder u0_1033(.a(t_2353), .b(t_2350), .o(t_2896), .cout(t_2897));
compressor_4_2 u2_1034(.a(t_2355), .b(t_2354), .c(t_2351), .d(t_2348), .cin(t_2895), .o(t_2898), .co(t_2899), .cout(t_2900));
half_adder u0_1035(.a(t_2361), .b(t_2358), .o(t_2901), .cout(t_2902));
compressor_4_2 u2_1036(.a(t_2363), .b(t_2362), .c(t_2359), .d(t_2356), .cin(t_2900), .o(t_2903), .co(t_2904), .cout(t_2905));
half_adder u0_1037(.a(t_2369), .b(t_2366), .o(t_2906), .cout(t_2907));
compressor_4_2 u2_1038(.a(t_2371), .b(t_2370), .c(t_2367), .d(t_2364), .cin(t_2905), .o(t_2908), .co(t_2909), .cout(t_2910));
half_adder u0_1039(.a(t_2377), .b(t_2374), .o(t_2911), .cout(t_2912));
compressor_4_2 u2_1040(.a(t_2378), .b(t_2375), .c(t_2372), .d(t_1429), .cin(t_2910), .o(t_2913), .co(t_2914), .cout(t_2915));
half_adder u0_1041(.a(t_2382), .b(t_2379), .o(t_2916), .cout(t_2917));
compressor_4_2 u2_1042(.a(t_2388), .b(t_2385), .c(t_2383), .d(t_2380), .cin(t_2915), .o(t_2918), .co(t_2919), .cout(t_2920));
compressor_4_2 u2_1043(.a(t_2394), .b(t_2391), .c(t_2389), .d(t_2386), .cin(t_2920), .o(t_2921), .co(t_2922), .cout(t_2923));
compressor_4_2 u2_1044(.a(t_2397), .b(t_2395), .c(t_2392), .d(t_1465), .cin(t_2923), .o(t_2924), .co(t_2925), .cout(t_2926));
compressor_4_2 u2_1045(.a(t_2406), .b(t_2403), .c(t_2401), .d(t_2398), .cin(t_2926), .o(t_2927), .co(t_2928), .cout(t_2929));
compressor_4_2 u2_1046(.a(t_2412), .b(t_2409), .c(t_2407), .d(t_2404), .cin(t_2929), .o(t_2930), .co(t_2931), .cout(t_2932));
compressor_4_2 u2_1047(.a(t_2418), .b(t_2415), .c(t_2413), .d(t_2410), .cin(t_2932), .o(t_2933), .co(t_2934), .cout(t_2935));
compressor_4_2 u2_1048(.a(t_2424), .b(t_2421), .c(t_2419), .d(t_2416), .cin(t_2935), .o(t_2936), .co(t_2937), .cout(t_2938));
compressor_4_2 u2_1049(.a(t_2427), .b(t_2425), .c(t_2422), .d(t_1515), .cin(t_2938), .o(t_2939), .co(t_2940), .cout(t_2941));
compressor_4_2 u2_1050(.a(t_2435), .b(t_2432), .c(t_2431), .d(t_2428), .cin(t_2941), .o(t_2942), .co(t_2943), .cout(t_2944));
compressor_4_2 u2_1051(.a(t_2440), .b(t_2437), .c(t_2436), .d(t_2433), .cin(t_2944), .o(t_2945), .co(t_2946), .cout(t_2947));
compressor_4_2 u2_1052(.a(t_2445), .b(t_2442), .c(t_2441), .d(t_2438), .cin(t_2947), .o(t_2948), .co(t_2949), .cout(t_2950));
compressor_4_2 u2_1053(.a(t_2450), .b(t_2447), .c(t_2446), .d(t_2443), .cin(t_2950), .o(t_2951), .co(t_2952), .cout(t_2953));
compressor_4_2 u2_1054(.a(t_2455), .b(t_2452), .c(t_2451), .d(t_2448), .cin(t_2953), .o(t_2954), .co(t_2955), .cout(t_2956));
compressor_4_2 u2_1055(.a(t_2460), .b(t_2457), .c(t_2456), .d(t_2453), .cin(t_2956), .o(t_2957), .co(t_2958), .cout(t_2959));
compressor_4_2 u2_1056(.a(t_2465), .b(t_2462), .c(t_2461), .d(t_2458), .cin(t_2959), .o(t_2960), .co(t_2961), .cout(t_2962));
compressor_4_2 u2_1057(.a(t_2467), .b(t_2466), .c(t_2463), .d(t_1577), .cin(t_2962), .o(t_2963), .co(t_2964), .cout(t_2965));
compressor_3_2 u1_1058(.a(t_2470), .b(t_2468), .cin(t_2965), .o(t_2966), .cout(t_2967));
half_adder u0_1059(.a(t_2473), .b(t_2471), .o(t_2968), .cout(t_2969));
compressor_3_2 u1_1060(.a(t_2476), .b(t_2474), .cin(t_1595), .o(t_2970), .cout(t_2971));
half_adder u0_1061(.a(t_2479), .b(t_2477), .o(t_2972), .cout(t_2973));
half_adder u0_1062(.a(t_2482), .b(t_2480), .o(t_2974), .cout(t_2975));
half_adder u0_1063(.a(t_2485), .b(t_2483), .o(t_2976), .cout(t_2977));
half_adder u0_1064(.a(t_2488), .b(t_2486), .o(t_2978), .cout(t_2979));
compressor_3_2 u1_1065(.a(t_2491), .b(t_2489), .cin(t_1615), .o(t_2980), .cout(t_2981));
half_adder u0_1066(.a(t_2493), .b(t_2492), .o(t_2982), .cout(t_2983));
half_adder u0_1067(.a(t_2495), .b(t_2494), .o(t_2984), .cout(t_2985));
half_adder u0_1068(.a(t_2497), .b(t_2496), .o(t_2986), .cout(t_2987));
half_adder u0_1069(.a(t_2499), .b(t_2498), .o(t_2988), .cout(t_2989));
half_adder u0_1070(.a(t_2501), .b(t_2500), .o(t_2990), .cout(t_2991));
half_adder u0_1071(.a(t_2503), .b(t_2502), .o(t_2992), .cout());

/* u0_1072 Output nets */
wire t_2993,   t_2994;
/* u0_1073 Output nets */
wire t_2995,   t_2996;
/* u0_1074 Output nets */
wire t_2997,   t_2998;
/* u0_1075 Output nets */
wire t_2999,   t_3000;
/* u0_1076 Output nets */
wire t_3001,   t_3002;
/* u0_1077 Output nets */
wire t_3003,   t_3004;
/* u0_1078 Output nets */
wire t_3005,   t_3006;
/* u0_1079 Output nets */
wire t_3007,   t_3008;
/* u0_1080 Output nets */
wire t_3009,   t_3010;
/* u0_1081 Output nets */
wire t_3011,   t_3012;
/* u0_1082 Output nets */
wire t_3013,   t_3014;
/* u0_1083 Output nets */
wire t_3015,   t_3016;
/* u0_1084 Output nets */
wire t_3017,   t_3018;
/* u0_1085 Output nets */
wire t_3019,   t_3020;
/* u1_1086 Output nets */
wire t_3021,   t_3022;
/* u0_1087 Output nets */
wire t_3023,   t_3024;
/* u1_1088 Output nets */
wire t_3025,   t_3026;
/* u1_1089 Output nets */
wire t_3027,   t_3028;
/* u1_1090 Output nets */
wire t_3029,   t_3030;
/* u1_1091 Output nets */
wire t_3031,   t_3032;
/* u1_1092 Output nets */
wire t_3033,   t_3034;
/* u0_1093 Output nets */
wire t_3035,   t_3036;
/* u0_1094 Output nets */
wire t_3037,   t_3038;
/* u1_1095 Output nets */
wire t_3039,   t_3040;
/* u0_1096 Output nets */
wire t_3041,   t_3042;
/* u0_1097 Output nets */
wire t_3043,   t_3044;
/* u0_1098 Output nets */
wire t_3045,   t_3046;
/* u0_1099 Output nets */
wire t_3047,   t_3048;
/* u1_1100 Output nets */
wire t_3049,   t_3050;
/* u1_1101 Output nets */
wire t_3051,   t_3052;
/* u1_1102 Output nets */
wire t_3053,   t_3054;
/* u1_1103 Output nets */
wire t_3055,   t_3056;
/* u1_1104 Output nets */
wire t_3057,   t_3058;
/* u1_1105 Output nets */
wire t_3059,   t_3060;
/* u1_1106 Output nets */
wire t_3061,   t_3062;
/* u1_1107 Output nets */
wire t_3063,   t_3064;
/* u1_1108 Output nets */
wire t_3065,   t_3066;
/* u1_1109 Output nets */
wire t_3067,   t_3068;
/* u1_1110 Output nets */
wire t_3069,   t_3070;
/* u1_1111 Output nets */
wire t_3071,   t_3072;
/* u1_1112 Output nets */
wire t_3073,   t_3074;
/* u1_1113 Output nets */
wire t_3075,   t_3076;
/* u1_1114 Output nets */
wire t_3077,   t_3078;
/* u1_1115 Output nets */
wire t_3079,   t_3080;
/* u1_1116 Output nets */
wire t_3081,   t_3082;
/* u1_1117 Output nets */
wire t_3083,   t_3084;
/* u2_1118 Output nets */
wire t_3085,   t_3086,   t_3087;
/* u2_1119 Output nets */
wire t_3088,   t_3089,   t_3090;
/* u2_1120 Output nets */
wire t_3091,   t_3092,   t_3093;
/* u2_1121 Output nets */
wire t_3094,   t_3095,   t_3096;
/* u2_1122 Output nets */
wire t_3097,   t_3098,   t_3099;
/* u2_1123 Output nets */
wire t_3100,   t_3101,   t_3102;
/* u2_1124 Output nets */
wire t_3103,   t_3104,   t_3105;
/* u2_1125 Output nets */
wire t_3106,   t_3107,   t_3108;
/* u2_1126 Output nets */
wire t_3109,   t_3110,   t_3111;
/* u2_1127 Output nets */
wire t_3112,   t_3113,   t_3114;
/* u2_1128 Output nets */
wire t_3115,   t_3116,   t_3117;
/* u2_1129 Output nets */
wire t_3118,   t_3119,   t_3120;
/* u2_1130 Output nets */
wire t_3121,   t_3122,   t_3123;
/* u2_1131 Output nets */
wire t_3124,   t_3125,   t_3126;
/* u2_1132 Output nets */
wire t_3127,   t_3128,   t_3129;
/* u2_1133 Output nets */
wire t_3130,   t_3131,   t_3132;
/* u2_1134 Output nets */
wire t_3133,   t_3134,   t_3135;
/* u2_1135 Output nets */
wire t_3136,   t_3137,   t_3138;
/* u2_1136 Output nets */
wire t_3139,   t_3140,   t_3141;
/* u2_1137 Output nets */
wire t_3142,   t_3143,   t_3144;
/* u2_1138 Output nets */
wire t_3145,   t_3146,   t_3147;
/* u2_1139 Output nets */
wire t_3148,   t_3149,   t_3150;
/* u2_1140 Output nets */
wire t_3151,   t_3152,   t_3153;
/* u2_1141 Output nets */
wire t_3154,   t_3155,   t_3156;
/* u2_1142 Output nets */
wire t_3157,   t_3158,   t_3159;
/* u2_1143 Output nets */
wire t_3160,   t_3161,   t_3162;
/* u2_1144 Output nets */
wire t_3163,   t_3164,   t_3165;
/* u2_1145 Output nets */
wire t_3166,   t_3167,   t_3168;
/* u2_1146 Output nets */
wire t_3169,   t_3170,   t_3171;
/* u2_1147 Output nets */
wire t_3172,   t_3173,   t_3174;
/* u2_1148 Output nets */
wire t_3175,   t_3176,   t_3177;
/* u2_1149 Output nets */
wire t_3178,   t_3179,   t_3180;
/* u2_1150 Output nets */
wire t_3181,   t_3182,   t_3183;
/* u2_1151 Output nets */
wire t_3184,   t_3185,   t_3186;
/* u2_1152 Output nets */
wire t_3187,   t_3188,   t_3189;
/* u2_1153 Output nets */
wire t_3190,   t_3191,   t_3192;
/* u2_1154 Output nets */
wire t_3193,   t_3194,   t_3195;
/* u2_1155 Output nets */
wire t_3196,   t_3197,   t_3198;
/* u2_1156 Output nets */
wire t_3199,   t_3200,   t_3201;
/* u2_1157 Output nets */
wire t_3202,   t_3203,   t_3204;
/* u2_1158 Output nets */
wire t_3205,   t_3206,   t_3207;
/* u2_1159 Output nets */
wire t_3208,   t_3209,   t_3210;
/* u2_1160 Output nets */
wire t_3211,   t_3212,   t_3213;
/* u2_1161 Output nets */
wire t_3214,   t_3215,   t_3216;
/* u2_1162 Output nets */
wire t_3217,   t_3218,   t_3219;
/* u2_1163 Output nets */
wire t_3220,   t_3221,   t_3222;
/* u2_1164 Output nets */
wire t_3223,   t_3224,   t_3225;
/* u2_1165 Output nets */
wire t_3226,   t_3227,   t_3228;
/* u1_1166 Output nets */
wire t_3229,   t_3230;
/* u0_1167 Output nets */
wire t_3231,   t_3232;
/* u1_1168 Output nets */
wire t_3233,   t_3234;
/* u0_1169 Output nets */
wire t_3235,   t_3236;
/* u0_1170 Output nets */
wire t_3237,   t_3238;
/* u0_1171 Output nets */
wire t_3239,   t_3240;
/* u0_1172 Output nets */
wire t_3241,   t_3242;
/* u1_1173 Output nets */
wire t_3243,   t_3244;
/* u0_1174 Output nets */
wire t_3245,   t_3246;
/* u0_1175 Output nets */
wire t_3247,   t_3248;
/* u0_1176 Output nets */
wire t_3249,   t_3250;
/* u0_1177 Output nets */
wire t_3251,   t_3252;
/* u0_1178 Output nets */
wire t_3253,   t_3254;
/* u0_1179 Output nets */
wire t_3255,   t_3256;
/* u0_1180 Output nets */
wire t_3257,   t_3258;
/* u0_1181 Output nets */
wire t_3259,   t_3260;
/* u0_1182 Output nets */
wire t_3261,   t_3262;
/* u0_1183 Output nets */
wire t_3263,   t_3264;
/* u0_1184 Output nets */
wire t_3265,   t_3266;
/* u0_1185 Output nets */
wire t_3267,   t_3268;
/* u0_1186 Output nets */
wire t_3269,   t_3270;
/* u0_1187 Output nets */
wire t_3271,   t_3272;
/* u0_1188 Output nets */
wire t_3273,   t_3274;
/* u0_1189 Output nets */
wire t_3275,   t_3276;
/* u0_1190 Output nets */
wire t_3277,   t_3278;
/* u0_1191 Output nets */
wire t_3279,   t_3280;
/* u0_1192 Output nets */
wire t_3281,   t_3282;
/* u0_1193 Output nets */
wire t_3283,   t_3284;
/* u0_1194 Output nets */
wire t_3285,   t_3286;
/* u0_1195 Output nets */
wire t_3287;

/* compress stage 4 */
half_adder u0_1072(.a(t_2505), .b(t_1633), .o(t_2993), .cout(t_2994));
half_adder u0_1073(.a(t_2508), .b(t_2507), .o(t_2995), .cout(t_2996));
half_adder u0_1074(.a(t_2510), .b(t_2509), .o(t_2997), .cout(t_2998));
half_adder u0_1075(.a(t_2512), .b(t_2511), .o(t_2999), .cout(t_3000));
half_adder u0_1076(.a(t_2514), .b(t_2513), .o(t_3001), .cout(t_3002));
half_adder u0_1077(.a(t_2516), .b(t_2515), .o(t_3003), .cout(t_3004));
half_adder u0_1078(.a(t_2518), .b(t_2517), .o(t_3005), .cout(t_3006));
half_adder u0_1079(.a(t_2520), .b(t_2519), .o(t_3007), .cout(t_3008));
half_adder u0_1080(.a(t_2522), .b(t_2521), .o(t_3009), .cout(t_3010));
half_adder u0_1081(.a(t_2524), .b(t_2523), .o(t_3011), .cout(t_3012));
half_adder u0_1082(.a(t_2526), .b(t_2525), .o(t_3013), .cout(t_3014));
half_adder u0_1083(.a(t_2528), .b(t_2527), .o(t_3015), .cout(t_3016));
half_adder u0_1084(.a(t_2530), .b(t_2529), .o(t_3017), .cout(t_3018));
half_adder u0_1085(.a(t_2532), .b(t_2531), .o(t_3019), .cout(t_3020));
compressor_3_2 u1_1086(.a(t_2534), .b(t_2533), .cin(t_1671), .o(t_3021), .cout(t_3022));
half_adder u0_1087(.a(t_2536), .b(t_2535), .o(t_3023), .cout(t_3024));
compressor_3_2 u1_1088(.a(t_2538), .b(t_2537), .cin(t_1682), .o(t_3025), .cout(t_3026));
compressor_3_2 u1_1089(.a(t_2540), .b(t_2539), .cin(t_1687), .o(t_3027), .cout(t_3028));
compressor_3_2 u1_1090(.a(t_2542), .b(t_2541), .cin(t_1692), .o(t_3029), .cout(t_3030));
compressor_3_2 u1_1091(.a(t_2544), .b(t_2543), .cin(t_1697), .o(t_3031), .cout(t_3032));
compressor_3_2 u1_1092(.a(t_2546), .b(t_2545), .cin(t_1702), .o(t_3033), .cout(t_3034));
half_adder u0_1093(.a(t_2548), .b(t_2547), .o(t_3035), .cout(t_3036));
half_adder u0_1094(.a(t_2551), .b(t_2549), .o(t_3037), .cout(t_3038));
compressor_3_2 u1_1095(.a(t_2554), .b(t_2552), .cin(t_1717), .o(t_3039), .cout(t_3040));
half_adder u0_1096(.a(t_2557), .b(t_2555), .o(t_3041), .cout(t_3042));
half_adder u0_1097(.a(t_2560), .b(t_2558), .o(t_3043), .cout(t_3044));
half_adder u0_1098(.a(t_2563), .b(t_2561), .o(t_3045), .cout(t_3046));
half_adder u0_1099(.a(t_2566), .b(t_2564), .o(t_3047), .cout(t_3048));
compressor_3_2 u1_1100(.a(t_2569), .b(t_2567), .cin(t_1746), .o(t_3049), .cout(t_3050));
compressor_3_2 u1_1101(.a(t_2572), .b(t_2570), .cin(t_1755), .o(t_3051), .cout(t_3052));
compressor_3_2 u1_1102(.a(t_2578), .b(t_2575), .cin(t_2573), .o(t_3053), .cout(t_3054));
compressor_3_2 u1_1103(.a(t_2579), .b(t_2576), .cin(t_1769), .o(t_3055), .cout(t_3056));
compressor_3_2 u1_1104(.a(t_2586), .b(t_2583), .cin(t_2581), .o(t_3057), .cout(t_3058));
compressor_3_2 u1_1105(.a(t_2588), .b(t_2587), .cin(t_2584), .o(t_3059), .cout(t_3060));
compressor_3_2 u1_1106(.a(t_2593), .b(t_2592), .cin(t_2589), .o(t_3061), .cout(t_3062));
compressor_3_2 u1_1107(.a(t_2598), .b(t_2597), .cin(t_2594), .o(t_3063), .cout(t_3064));
compressor_3_2 u1_1108(.a(t_2603), .b(t_2602), .cin(t_2599), .o(t_3065), .cout(t_3066));
compressor_3_2 u1_1109(.a(t_2608), .b(t_2607), .cin(t_2604), .o(t_3067), .cout(t_3068));
compressor_3_2 u1_1110(.a(t_2613), .b(t_2612), .cin(t_2609), .o(t_3069), .cout(t_3070));
compressor_3_2 u1_1111(.a(t_2618), .b(t_2617), .cin(t_2614), .o(t_3071), .cout(t_3072));
compressor_3_2 u1_1112(.a(t_2623), .b(t_2622), .cin(t_2619), .o(t_3073), .cout(t_3074));
compressor_3_2 u1_1113(.a(t_2628), .b(t_2627), .cin(t_2624), .o(t_3075), .cout(t_3076));
compressor_3_2 u1_1114(.a(t_2633), .b(t_2632), .cin(t_2629), .o(t_3077), .cout(t_3078));
compressor_3_2 u1_1115(.a(t_2638), .b(t_2637), .cin(t_2634), .o(t_3079), .cout(t_3080));
compressor_3_2 u1_1116(.a(t_2643), .b(t_2642), .cin(t_2639), .o(t_3081), .cout(t_3082));
compressor_3_2 u1_1117(.a(t_2648), .b(t_2647), .cin(t_2644), .o(t_3083), .cout(t_3084));
compressor_4_2 u2_1118(.a(t_2656), .b(t_2653), .c(t_2652), .d(t_2649), .cin(t_1897), .o(t_3085), .co(t_3086), .cout(t_3087));
compressor_4_2 u2_1119(.a(t_2661), .b(t_2658), .c(t_2657), .d(t_2654), .cin(t_3087), .o(t_3088), .co(t_3089), .cout(t_3090));
compressor_4_2 u2_1120(.a(t_2663), .b(t_2662), .c(t_2659), .d(t_1920), .cin(t_3090), .o(t_3091), .co(t_3092), .cout(t_3093));
compressor_4_2 u2_1121(.a(t_2668), .b(t_2667), .c(t_2664), .d(t_1931), .cin(t_3093), .o(t_3094), .co(t_3095), .cout(t_3096));
compressor_4_2 u2_1122(.a(t_2673), .b(t_2672), .c(t_2669), .d(t_1942), .cin(t_3096), .o(t_3097), .co(t_3098), .cout(t_3099));
compressor_4_2 u2_1123(.a(t_2678), .b(t_2677), .c(t_2674), .d(t_1953), .cin(t_3099), .o(t_3100), .co(t_3101), .cout(t_3102));
compressor_4_2 u2_1124(.a(t_2683), .b(t_2682), .c(t_2679), .d(t_1964), .cin(t_3102), .o(t_3103), .co(t_3104), .cout(t_3105));
compressor_4_2 u2_1125(.a(t_2691), .b(t_2688), .c(t_2687), .d(t_2684), .cin(t_3105), .o(t_3106), .co(t_3107), .cout(t_3108));
compressor_4_2 u2_1126(.a(t_2697), .b(t_2694), .c(t_2692), .d(t_2689), .cin(t_3108), .o(t_3109), .co(t_3110), .cout(t_3111));
compressor_4_2 u2_1127(.a(t_2700), .b(t_2698), .c(t_2695), .d(t_1997), .cin(t_3111), .o(t_3112), .co(t_3113), .cout(t_3114));
compressor_4_2 u2_1128(.a(t_2709), .b(t_2706), .c(t_2704), .d(t_2701), .cin(t_3114), .o(t_3115), .co(t_3116), .cout(t_3117));
compressor_4_2 u2_1129(.a(t_2715), .b(t_2712), .c(t_2710), .d(t_2707), .cin(t_3117), .o(t_3118), .co(t_3119), .cout(t_3120));
compressor_4_2 u2_1130(.a(t_2721), .b(t_2718), .c(t_2716), .d(t_2713), .cin(t_3120), .o(t_3121), .co(t_3122), .cout(t_3123));
compressor_4_2 u2_1131(.a(t_2727), .b(t_2724), .c(t_2722), .d(t_2719), .cin(t_3123), .o(t_3124), .co(t_3125), .cout(t_3126));
compressor_4_2 u2_1132(.a(t_2730), .b(t_2728), .c(t_2725), .d(t_2056), .cin(t_3126), .o(t_3127), .co(t_3128), .cout(t_3129));
compressor_4_2 u2_1133(.a(t_2736), .b(t_2734), .c(t_2731), .d(t_2068), .cin(t_3129), .o(t_3130), .co(t_3131), .cout(t_3132));
compressor_4_2 u2_1134(.a(t_2745), .b(t_2742), .c(t_2740), .d(t_2737), .cin(t_3132), .o(t_3133), .co(t_3134), .cout(t_3135));
compressor_4_2 u2_1135(.a(t_2751), .b(t_2748), .c(t_2746), .d(t_2743), .cin(t_3135), .o(t_3136), .co(t_3137), .cout(t_3138));
compressor_4_2 u2_1136(.a(t_2754), .b(t_2752), .c(t_2749), .d(t_2104), .cin(t_3138), .o(t_3139), .co(t_3140), .cout(t_3141));
compressor_4_2 u2_1137(.a(t_2763), .b(t_2760), .c(t_2758), .d(t_2755), .cin(t_3141), .o(t_3142), .co(t_3143), .cout(t_3144));
compressor_4_2 u2_1138(.a(t_2769), .b(t_2766), .c(t_2764), .d(t_2761), .cin(t_3144), .o(t_3145), .co(t_3146), .cout(t_3147));
compressor_4_2 u2_1139(.a(t_2775), .b(t_2772), .c(t_2770), .d(t_2767), .cin(t_3147), .o(t_3148), .co(t_3149), .cout(t_3150));
compressor_4_2 u2_1140(.a(t_2781), .b(t_2778), .c(t_2776), .d(t_2773), .cin(t_3150), .o(t_3151), .co(t_3152), .cout(t_3153));
compressor_4_2 u2_1141(.a(t_2784), .b(t_2782), .c(t_2779), .d(t_2164), .cin(t_3153), .o(t_3154), .co(t_3155), .cout(t_3156));
compressor_4_2 u2_1142(.a(t_2793), .b(t_2790), .c(t_2788), .d(t_2785), .cin(t_3156), .o(t_3157), .co(t_3158), .cout(t_3159));
compressor_4_2 u2_1143(.a(t_2799), .b(t_2796), .c(t_2794), .d(t_2791), .cin(t_3159), .o(t_3160), .co(t_3161), .cout(t_3162));
compressor_4_2 u2_1144(.a(t_2805), .b(t_2802), .c(t_2800), .d(t_2797), .cin(t_3162), .o(t_3163), .co(t_3164), .cout(t_3165));
compressor_4_2 u2_1145(.a(t_2811), .b(t_2808), .c(t_2806), .d(t_2803), .cin(t_3165), .o(t_3166), .co(t_3167), .cout(t_3168));
compressor_4_2 u2_1146(.a(t_2817), .b(t_2814), .c(t_2812), .d(t_2809), .cin(t_3168), .o(t_3169), .co(t_3170), .cout(t_3171));
compressor_4_2 u2_1147(.a(t_2823), .b(t_2820), .c(t_2818), .d(t_2815), .cin(t_3171), .o(t_3172), .co(t_3173), .cout(t_3174));
compressor_4_2 u2_1148(.a(t_2829), .b(t_2826), .c(t_2824), .d(t_2821), .cin(t_3174), .o(t_3175), .co(t_3176), .cout(t_3177));
compressor_4_2 u2_1149(.a(t_2835), .b(t_2832), .c(t_2830), .d(t_2827), .cin(t_3177), .o(t_3178), .co(t_3179), .cout(t_3180));
compressor_4_2 u2_1150(.a(t_2841), .b(t_2838), .c(t_2836), .d(t_2833), .cin(t_3180), .o(t_3181), .co(t_3182), .cout(t_3183));
compressor_4_2 u2_1151(.a(t_2846), .b(t_2843), .c(t_2842), .d(t_2839), .cin(t_3183), .o(t_3184), .co(t_3185), .cout(t_3186));
compressor_4_2 u2_1152(.a(t_2851), .b(t_2848), .c(t_2847), .d(t_2844), .cin(t_3186), .o(t_3187), .co(t_3188), .cout(t_3189));
compressor_4_2 u2_1153(.a(t_2856), .b(t_2853), .c(t_2852), .d(t_2849), .cin(t_3189), .o(t_3190), .co(t_3191), .cout(t_3192));
compressor_4_2 u2_1154(.a(t_2861), .b(t_2858), .c(t_2857), .d(t_2854), .cin(t_3192), .o(t_3193), .co(t_3194), .cout(t_3195));
compressor_4_2 u2_1155(.a(t_2866), .b(t_2863), .c(t_2862), .d(t_2859), .cin(t_3195), .o(t_3196), .co(t_3197), .cout(t_3198));
compressor_4_2 u2_1156(.a(t_2871), .b(t_2868), .c(t_2867), .d(t_2864), .cin(t_3198), .o(t_3199), .co(t_3200), .cout(t_3201));
compressor_4_2 u2_1157(.a(t_2876), .b(t_2873), .c(t_2872), .d(t_2869), .cin(t_3201), .o(t_3202), .co(t_3203), .cout(t_3204));
compressor_4_2 u2_1158(.a(t_2881), .b(t_2878), .c(t_2877), .d(t_2874), .cin(t_3204), .o(t_3205), .co(t_3206), .cout(t_3207));
compressor_4_2 u2_1159(.a(t_2886), .b(t_2883), .c(t_2882), .d(t_2879), .cin(t_3207), .o(t_3208), .co(t_3209), .cout(t_3210));
compressor_4_2 u2_1160(.a(t_2891), .b(t_2888), .c(t_2887), .d(t_2884), .cin(t_3210), .o(t_3211), .co(t_3212), .cout(t_3213));
compressor_4_2 u2_1161(.a(t_2896), .b(t_2893), .c(t_2892), .d(t_2889), .cin(t_3213), .o(t_3214), .co(t_3215), .cout(t_3216));
compressor_4_2 u2_1162(.a(t_2901), .b(t_2898), .c(t_2897), .d(t_2894), .cin(t_3216), .o(t_3217), .co(t_3218), .cout(t_3219));
compressor_4_2 u2_1163(.a(t_2906), .b(t_2903), .c(t_2902), .d(t_2899), .cin(t_3219), .o(t_3220), .co(t_3221), .cout(t_3222));
compressor_4_2 u2_1164(.a(t_2911), .b(t_2908), .c(t_2907), .d(t_2904), .cin(t_3222), .o(t_3223), .co(t_3224), .cout(t_3225));
compressor_4_2 u2_1165(.a(t_2916), .b(t_2913), .c(t_2912), .d(t_2909), .cin(t_3225), .o(t_3226), .co(t_3227), .cout(t_3228));
compressor_3_2 u1_1166(.a(t_2917), .b(t_2914), .cin(t_3228), .o(t_3229), .cout(t_3230));
half_adder u0_1167(.a(t_2921), .b(t_2919), .o(t_3231), .cout(t_3232));
compressor_3_2 u1_1168(.a(t_2924), .b(t_2922), .cin(t_2400), .o(t_3233), .cout(t_3234));
half_adder u0_1169(.a(t_2927), .b(t_2925), .o(t_3235), .cout(t_3236));
half_adder u0_1170(.a(t_2930), .b(t_2928), .o(t_3237), .cout(t_3238));
half_adder u0_1171(.a(t_2933), .b(t_2931), .o(t_3239), .cout(t_3240));
half_adder u0_1172(.a(t_2936), .b(t_2934), .o(t_3241), .cout(t_3242));
compressor_3_2 u1_1173(.a(t_2939), .b(t_2937), .cin(t_2430), .o(t_3243), .cout(t_3244));
half_adder u0_1174(.a(t_2942), .b(t_2940), .o(t_3245), .cout(t_3246));
half_adder u0_1175(.a(t_2945), .b(t_2943), .o(t_3247), .cout(t_3248));
half_adder u0_1176(.a(t_2948), .b(t_2946), .o(t_3249), .cout(t_3250));
half_adder u0_1177(.a(t_2951), .b(t_2949), .o(t_3251), .cout(t_3252));
half_adder u0_1178(.a(t_2954), .b(t_2952), .o(t_3253), .cout(t_3254));
half_adder u0_1179(.a(t_2957), .b(t_2955), .o(t_3255), .cout(t_3256));
half_adder u0_1180(.a(t_2960), .b(t_2958), .o(t_3257), .cout(t_3258));
half_adder u0_1181(.a(t_2963), .b(t_2961), .o(t_3259), .cout(t_3260));
half_adder u0_1182(.a(t_2966), .b(t_2964), .o(t_3261), .cout(t_3262));
half_adder u0_1183(.a(t_2968), .b(t_2967), .o(t_3263), .cout(t_3264));
half_adder u0_1184(.a(t_2970), .b(t_2969), .o(t_3265), .cout(t_3266));
half_adder u0_1185(.a(t_2972), .b(t_2971), .o(t_3267), .cout(t_3268));
half_adder u0_1186(.a(t_2974), .b(t_2973), .o(t_3269), .cout(t_3270));
half_adder u0_1187(.a(t_2976), .b(t_2975), .o(t_3271), .cout(t_3272));
half_adder u0_1188(.a(t_2978), .b(t_2977), .o(t_3273), .cout(t_3274));
half_adder u0_1189(.a(t_2980), .b(t_2979), .o(t_3275), .cout(t_3276));
half_adder u0_1190(.a(t_2982), .b(t_2981), .o(t_3277), .cout(t_3278));
half_adder u0_1191(.a(t_2984), .b(t_2983), .o(t_3279), .cout(t_3280));
half_adder u0_1192(.a(t_2986), .b(t_2985), .o(t_3281), .cout(t_3282));
half_adder u0_1193(.a(t_2988), .b(t_2987), .o(t_3283), .cout(t_3284));
half_adder u0_1194(.a(t_2990), .b(t_2989), .o(t_3285), .cout(t_3286));
half_adder u0_1195(.a(t_2992), .b(t_2991), .o(t_3287), .cout());

/* u0_1196 Output nets */
wire t_3288,   t_3289;
/* u0_1197 Output nets */
wire t_3290,   t_3291;
/* u0_1198 Output nets */
wire t_3292,   t_3293;
/* u0_1199 Output nets */
wire t_3294,   t_3295;
/* u0_1200 Output nets */
wire t_3296,   t_3297;
/* u0_1201 Output nets */
wire t_3298,   t_3299;
/* u0_1202 Output nets */
wire t_3300,   t_3301;
/* u0_1203 Output nets */
wire t_3302,   t_3303;
/* u0_1204 Output nets */
wire t_3304,   t_3305;
/* u0_1205 Output nets */
wire t_3306,   t_3307;
/* u0_1206 Output nets */
wire t_3308,   t_3309;
/* u0_1207 Output nets */
wire t_3310,   t_3311;
/* u0_1208 Output nets */
wire t_3312,   t_3313;
/* u0_1209 Output nets */
wire t_3314,   t_3315;
/* u0_1210 Output nets */
wire t_3316,   t_3317;
/* u0_1211 Output nets */
wire t_3318,   t_3319;
/* u0_1212 Output nets */
wire t_3320,   t_3321;
/* u0_1213 Output nets */
wire t_3322,   t_3323;
/* u0_1214 Output nets */
wire t_3324,   t_3325;
/* u0_1215 Output nets */
wire t_3326,   t_3327;
/* u0_1216 Output nets */
wire t_3328,   t_3329;
/* u0_1217 Output nets */
wire t_3330,   t_3331;
/* u0_1218 Output nets */
wire t_3332,   t_3333;
/* u0_1219 Output nets */
wire t_3334,   t_3335;
/* u0_1220 Output nets */
wire t_3336,   t_3337;
/* u0_1221 Output nets */
wire t_3338,   t_3339;
/* u0_1222 Output nets */
wire t_3340,   t_3341;
/* u0_1223 Output nets */
wire t_3342,   t_3343;
/* u0_1224 Output nets */
wire t_3344,   t_3345;
/* u0_1225 Output nets */
wire t_3346,   t_3347;
/* u1_1226 Output nets */
wire t_3348,   t_3349;
/* u0_1227 Output nets */
wire t_3350,   t_3351;
/* u1_1228 Output nets */
wire t_3352,   t_3353;
/* u1_1229 Output nets */
wire t_3354,   t_3355;
/* u1_1230 Output nets */
wire t_3356,   t_3357;
/* u1_1231 Output nets */
wire t_3358,   t_3359;
/* u1_1232 Output nets */
wire t_3360,   t_3361;
/* u1_1233 Output nets */
wire t_3362,   t_3363;
/* u1_1234 Output nets */
wire t_3364,   t_3365;
/* u1_1235 Output nets */
wire t_3366,   t_3367;
/* u1_1236 Output nets */
wire t_3368,   t_3369;
/* u1_1237 Output nets */
wire t_3370,   t_3371;
/* u1_1238 Output nets */
wire t_3372,   t_3373;
/* u1_1239 Output nets */
wire t_3374,   t_3375;
/* u1_1240 Output nets */
wire t_3376,   t_3377;
/* u0_1241 Output nets */
wire t_3378,   t_3379;
/* u0_1242 Output nets */
wire t_3380,   t_3381;
/* u1_1243 Output nets */
wire t_3382,   t_3383;
/* u1_1244 Output nets */
wire t_3384,   t_3385;
/* u1_1245 Output nets */
wire t_3386,   t_3387;
/* u1_1246 Output nets */
wire t_3388,   t_3389;
/* u1_1247 Output nets */
wire t_3390,   t_3391;
/* u0_1248 Output nets */
wire t_3392,   t_3393;
/* u0_1249 Output nets */
wire t_3394,   t_3395;
/* u1_1250 Output nets */
wire t_3396,   t_3397;
/* u0_1251 Output nets */
wire t_3398,   t_3399;
/* u0_1252 Output nets */
wire t_3400,   t_3401;
/* u0_1253 Output nets */
wire t_3402,   t_3403;
/* u0_1254 Output nets */
wire t_3404,   t_3405;
/* u1_1255 Output nets */
wire t_3406,   t_3407;
/* u1_1256 Output nets */
wire t_3408,   t_3409;
/* u0_1257 Output nets */
wire t_3410,   t_3411;
/* u0_1258 Output nets */
wire t_3412,   t_3413;
/* u1_1259 Output nets */
wire t_3414,   t_3415;
/* u0_1260 Output nets */
wire t_3416,   t_3417;
/* u0_1261 Output nets */
wire t_3418,   t_3419;
/* u0_1262 Output nets */
wire t_3420,   t_3421;
/* u0_1263 Output nets */
wire t_3422,   t_3423;
/* u1_1264 Output nets */
wire t_3424,   t_3425;
/* u0_1265 Output nets */
wire t_3426,   t_3427;
/* u0_1266 Output nets */
wire t_3428,   t_3429;
/* u0_1267 Output nets */
wire t_3430,   t_3431;
/* u0_1268 Output nets */
wire t_3432,   t_3433;
/* u0_1269 Output nets */
wire t_3434,   t_3435;
/* u0_1270 Output nets */
wire t_3436,   t_3437;
/* u0_1271 Output nets */
wire t_3438,   t_3439;
/* u0_1272 Output nets */
wire t_3440,   t_3441;
/* u0_1273 Output nets */
wire t_3442,   t_3443;
/* u0_1274 Output nets */
wire t_3444,   t_3445;
/* u0_1275 Output nets */
wire t_3446,   t_3447;
/* u0_1276 Output nets */
wire t_3448,   t_3449;
/* u0_1277 Output nets */
wire t_3450,   t_3451;
/* u0_1278 Output nets */
wire t_3452,   t_3453;
/* u0_1279 Output nets */
wire t_3454,   t_3455;
/* u0_1280 Output nets */
wire t_3456,   t_3457;
/* u0_1281 Output nets */
wire t_3458,   t_3459;
/* u0_1282 Output nets */
wire t_3460,   t_3461;
/* u0_1283 Output nets */
wire t_3462,   t_3463;
/* u0_1284 Output nets */
wire t_3464,   t_3465;
/* u0_1285 Output nets */
wire t_3466,   t_3467;
/* u0_1286 Output nets */
wire t_3468,   t_3469;
/* u0_1287 Output nets */
wire t_3470,   t_3471;
/* u0_1288 Output nets */
wire t_3472,   t_3473;
/* u1_1289 Output nets */
wire t_3474,   t_3475;
/* u0_1290 Output nets */
wire t_3476,   t_3477;
/* u0_1291 Output nets */
wire t_3478,   t_3479;
/* u0_1292 Output nets */
wire t_3480,   t_3481;
/* u0_1293 Output nets */
wire t_3482,   t_3483;
/* u0_1294 Output nets */
wire t_3484,   t_3485;
/* u0_1295 Output nets */
wire t_3486,   t_3487;
/* u0_1296 Output nets */
wire t_3488,   t_3489;
/* u0_1297 Output nets */
wire t_3490,   t_3491;
/* u0_1298 Output nets */
wire t_3492,   t_3493;
/* u0_1299 Output nets */
wire t_3494,   t_3495;
/* u0_1300 Output nets */
wire t_3496,   t_3497;
/* u0_1301 Output nets */
wire t_3498,   t_3499;
/* u0_1302 Output nets */
wire t_3500,   t_3501;
/* u0_1303 Output nets */
wire t_3502,   t_3503;
/* u0_1304 Output nets */
wire t_3504,   t_3505;
/* u0_1305 Output nets */
wire t_3506,   t_3507;
/* u0_1306 Output nets */
wire t_3508,   t_3509;
/* u0_1307 Output nets */
wire t_3510,   t_3511;
/* u0_1308 Output nets */
wire t_3512,   t_3513;
/* u0_1309 Output nets */
wire t_3514,   t_3515;
/* u0_1310 Output nets */
wire t_3516,   t_3517;
/* u0_1311 Output nets */
wire t_3518,   t_3519;
/* u0_1312 Output nets */
wire t_3520,   t_3521;
/* u0_1313 Output nets */
wire t_3522,   t_3523;
/* u0_1314 Output nets */
wire t_3524,   t_3525;
/* u0_1315 Output nets */
wire t_3526,   t_3527;
/* u0_1316 Output nets */
wire t_3528,   t_3529;
/* u0_1317 Output nets */
wire t_3530,   t_3531;
/* u0_1318 Output nets */
wire t_3532;

/* compress stage 5 */
half_adder u0_1196(.a(t_2994), .b(t_2506), .o(t_3288), .cout(t_3289));
half_adder u0_1197(.a(t_2997), .b(t_2996), .o(t_3290), .cout(t_3291));
half_adder u0_1198(.a(t_2999), .b(t_2998), .o(t_3292), .cout(t_3293));
half_adder u0_1199(.a(t_3001), .b(t_3000), .o(t_3294), .cout(t_3295));
half_adder u0_1200(.a(t_3003), .b(t_3002), .o(t_3296), .cout(t_3297));
half_adder u0_1201(.a(t_3005), .b(t_3004), .o(t_3298), .cout(t_3299));
half_adder u0_1202(.a(t_3007), .b(t_3006), .o(t_3300), .cout(t_3301));
half_adder u0_1203(.a(t_3009), .b(t_3008), .o(t_3302), .cout(t_3303));
half_adder u0_1204(.a(t_3011), .b(t_3010), .o(t_3304), .cout(t_3305));
half_adder u0_1205(.a(t_3013), .b(t_3012), .o(t_3306), .cout(t_3307));
half_adder u0_1206(.a(t_3015), .b(t_3014), .o(t_3308), .cout(t_3309));
half_adder u0_1207(.a(t_3017), .b(t_3016), .o(t_3310), .cout(t_3311));
half_adder u0_1208(.a(t_3019), .b(t_3018), .o(t_3312), .cout(t_3313));
half_adder u0_1209(.a(t_3021), .b(t_3020), .o(t_3314), .cout(t_3315));
half_adder u0_1210(.a(t_3023), .b(t_3022), .o(t_3316), .cout(t_3317));
half_adder u0_1211(.a(t_3025), .b(t_3024), .o(t_3318), .cout(t_3319));
half_adder u0_1212(.a(t_3027), .b(t_3026), .o(t_3320), .cout(t_3321));
half_adder u0_1213(.a(t_3029), .b(t_3028), .o(t_3322), .cout(t_3323));
half_adder u0_1214(.a(t_3031), .b(t_3030), .o(t_3324), .cout(t_3325));
half_adder u0_1215(.a(t_3033), .b(t_3032), .o(t_3326), .cout(t_3327));
half_adder u0_1216(.a(t_3035), .b(t_3034), .o(t_3328), .cout(t_3329));
half_adder u0_1217(.a(t_3037), .b(t_3036), .o(t_3330), .cout(t_3331));
half_adder u0_1218(.a(t_3039), .b(t_3038), .o(t_3332), .cout(t_3333));
half_adder u0_1219(.a(t_3041), .b(t_3040), .o(t_3334), .cout(t_3335));
half_adder u0_1220(.a(t_3043), .b(t_3042), .o(t_3336), .cout(t_3337));
half_adder u0_1221(.a(t_3045), .b(t_3044), .o(t_3338), .cout(t_3339));
half_adder u0_1222(.a(t_3047), .b(t_3046), .o(t_3340), .cout(t_3341));
half_adder u0_1223(.a(t_3049), .b(t_3048), .o(t_3342), .cout(t_3343));
half_adder u0_1224(.a(t_3051), .b(t_3050), .o(t_3344), .cout(t_3345));
half_adder u0_1225(.a(t_3053), .b(t_3052), .o(t_3346), .cout(t_3347));
compressor_3_2 u1_1226(.a(t_3055), .b(t_3054), .cin(t_2580), .o(t_3348), .cout(t_3349));
half_adder u0_1227(.a(t_3057), .b(t_3056), .o(t_3350), .cout(t_3351));
compressor_3_2 u1_1228(.a(t_3059), .b(t_3058), .cin(t_2591), .o(t_3352), .cout(t_3353));
compressor_3_2 u1_1229(.a(t_3061), .b(t_3060), .cin(t_2596), .o(t_3354), .cout(t_3355));
compressor_3_2 u1_1230(.a(t_3063), .b(t_3062), .cin(t_2601), .o(t_3356), .cout(t_3357));
compressor_3_2 u1_1231(.a(t_3065), .b(t_3064), .cin(t_2606), .o(t_3358), .cout(t_3359));
compressor_3_2 u1_1232(.a(t_3067), .b(t_3066), .cin(t_2611), .o(t_3360), .cout(t_3361));
compressor_3_2 u1_1233(.a(t_3069), .b(t_3068), .cin(t_2616), .o(t_3362), .cout(t_3363));
compressor_3_2 u1_1234(.a(t_3071), .b(t_3070), .cin(t_2621), .o(t_3364), .cout(t_3365));
compressor_3_2 u1_1235(.a(t_3073), .b(t_3072), .cin(t_2626), .o(t_3366), .cout(t_3367));
compressor_3_2 u1_1236(.a(t_3075), .b(t_3074), .cin(t_2631), .o(t_3368), .cout(t_3369));
compressor_3_2 u1_1237(.a(t_3077), .b(t_3076), .cin(t_2636), .o(t_3370), .cout(t_3371));
compressor_3_2 u1_1238(.a(t_3079), .b(t_3078), .cin(t_2641), .o(t_3372), .cout(t_3373));
compressor_3_2 u1_1239(.a(t_3081), .b(t_3080), .cin(t_2646), .o(t_3374), .cout(t_3375));
compressor_3_2 u1_1240(.a(t_3083), .b(t_3082), .cin(t_2651), .o(t_3376), .cout(t_3377));
half_adder u0_1241(.a(t_3085), .b(t_3084), .o(t_3378), .cout(t_3379));
half_adder u0_1242(.a(t_3088), .b(t_3086), .o(t_3380), .cout(t_3381));
compressor_3_2 u1_1243(.a(t_3091), .b(t_3089), .cin(t_2666), .o(t_3382), .cout(t_3383));
compressor_3_2 u1_1244(.a(t_3094), .b(t_3092), .cin(t_2671), .o(t_3384), .cout(t_3385));
compressor_3_2 u1_1245(.a(t_3097), .b(t_3095), .cin(t_2676), .o(t_3386), .cout(t_3387));
compressor_3_2 u1_1246(.a(t_3100), .b(t_3098), .cin(t_2681), .o(t_3388), .cout(t_3389));
compressor_3_2 u1_1247(.a(t_3103), .b(t_3101), .cin(t_2686), .o(t_3390), .cout(t_3391));
half_adder u0_1248(.a(t_3106), .b(t_3104), .o(t_3392), .cout(t_3393));
half_adder u0_1249(.a(t_3109), .b(t_3107), .o(t_3394), .cout(t_3395));
compressor_3_2 u1_1250(.a(t_3112), .b(t_3110), .cin(t_2703), .o(t_3396), .cout(t_3397));
half_adder u0_1251(.a(t_3115), .b(t_3113), .o(t_3398), .cout(t_3399));
half_adder u0_1252(.a(t_3118), .b(t_3116), .o(t_3400), .cout(t_3401));
half_adder u0_1253(.a(t_3121), .b(t_3119), .o(t_3402), .cout(t_3403));
half_adder u0_1254(.a(t_3124), .b(t_3122), .o(t_3404), .cout(t_3405));
compressor_3_2 u1_1255(.a(t_3127), .b(t_3125), .cin(t_2733), .o(t_3406), .cout(t_3407));
compressor_3_2 u1_1256(.a(t_3130), .b(t_3128), .cin(t_2739), .o(t_3408), .cout(t_3409));
half_adder u0_1257(.a(t_3133), .b(t_3131), .o(t_3410), .cout(t_3411));
half_adder u0_1258(.a(t_3136), .b(t_3134), .o(t_3412), .cout(t_3413));
compressor_3_2 u1_1259(.a(t_3139), .b(t_3137), .cin(t_2757), .o(t_3414), .cout(t_3415));
half_adder u0_1260(.a(t_3142), .b(t_3140), .o(t_3416), .cout(t_3417));
half_adder u0_1261(.a(t_3145), .b(t_3143), .o(t_3418), .cout(t_3419));
half_adder u0_1262(.a(t_3148), .b(t_3146), .o(t_3420), .cout(t_3421));
half_adder u0_1263(.a(t_3151), .b(t_3149), .o(t_3422), .cout(t_3423));
compressor_3_2 u1_1264(.a(t_3154), .b(t_3152), .cin(t_2787), .o(t_3424), .cout(t_3425));
half_adder u0_1265(.a(t_3157), .b(t_3155), .o(t_3426), .cout(t_3427));
half_adder u0_1266(.a(t_3160), .b(t_3158), .o(t_3428), .cout(t_3429));
half_adder u0_1267(.a(t_3163), .b(t_3161), .o(t_3430), .cout(t_3431));
half_adder u0_1268(.a(t_3166), .b(t_3164), .o(t_3432), .cout(t_3433));
half_adder u0_1269(.a(t_3169), .b(t_3167), .o(t_3434), .cout(t_3435));
half_adder u0_1270(.a(t_3172), .b(t_3170), .o(t_3436), .cout(t_3437));
half_adder u0_1271(.a(t_3175), .b(t_3173), .o(t_3438), .cout(t_3439));
half_adder u0_1272(.a(t_3178), .b(t_3176), .o(t_3440), .cout(t_3441));
half_adder u0_1273(.a(t_3181), .b(t_3179), .o(t_3442), .cout(t_3443));
half_adder u0_1274(.a(t_3184), .b(t_3182), .o(t_3444), .cout(t_3445));
half_adder u0_1275(.a(t_3187), .b(t_3185), .o(t_3446), .cout(t_3447));
half_adder u0_1276(.a(t_3190), .b(t_3188), .o(t_3448), .cout(t_3449));
half_adder u0_1277(.a(t_3193), .b(t_3191), .o(t_3450), .cout(t_3451));
half_adder u0_1278(.a(t_3196), .b(t_3194), .o(t_3452), .cout(t_3453));
half_adder u0_1279(.a(t_3199), .b(t_3197), .o(t_3454), .cout(t_3455));
half_adder u0_1280(.a(t_3202), .b(t_3200), .o(t_3456), .cout(t_3457));
half_adder u0_1281(.a(t_3205), .b(t_3203), .o(t_3458), .cout(t_3459));
half_adder u0_1282(.a(t_3208), .b(t_3206), .o(t_3460), .cout(t_3461));
half_adder u0_1283(.a(t_3211), .b(t_3209), .o(t_3462), .cout(t_3463));
half_adder u0_1284(.a(t_3214), .b(t_3212), .o(t_3464), .cout(t_3465));
half_adder u0_1285(.a(t_3217), .b(t_3215), .o(t_3466), .cout(t_3467));
half_adder u0_1286(.a(t_3220), .b(t_3218), .o(t_3468), .cout(t_3469));
half_adder u0_1287(.a(t_3223), .b(t_3221), .o(t_3470), .cout(t_3471));
half_adder u0_1288(.a(t_3226), .b(t_3224), .o(t_3472), .cout(t_3473));
compressor_3_2 u1_1289(.a(t_3229), .b(t_3227), .cin(t_2918), .o(t_3474), .cout(t_3475));
half_adder u0_1290(.a(t_3231), .b(t_3230), .o(t_3476), .cout(t_3477));
half_adder u0_1291(.a(t_3233), .b(t_3232), .o(t_3478), .cout(t_3479));
half_adder u0_1292(.a(t_3235), .b(t_3234), .o(t_3480), .cout(t_3481));
half_adder u0_1293(.a(t_3237), .b(t_3236), .o(t_3482), .cout(t_3483));
half_adder u0_1294(.a(t_3239), .b(t_3238), .o(t_3484), .cout(t_3485));
half_adder u0_1295(.a(t_3241), .b(t_3240), .o(t_3486), .cout(t_3487));
half_adder u0_1296(.a(t_3243), .b(t_3242), .o(t_3488), .cout(t_3489));
half_adder u0_1297(.a(t_3245), .b(t_3244), .o(t_3490), .cout(t_3491));
half_adder u0_1298(.a(t_3247), .b(t_3246), .o(t_3492), .cout(t_3493));
half_adder u0_1299(.a(t_3249), .b(t_3248), .o(t_3494), .cout(t_3495));
half_adder u0_1300(.a(t_3251), .b(t_3250), .o(t_3496), .cout(t_3497));
half_adder u0_1301(.a(t_3253), .b(t_3252), .o(t_3498), .cout(t_3499));
half_adder u0_1302(.a(t_3255), .b(t_3254), .o(t_3500), .cout(t_3501));
half_adder u0_1303(.a(t_3257), .b(t_3256), .o(t_3502), .cout(t_3503));
half_adder u0_1304(.a(t_3259), .b(t_3258), .o(t_3504), .cout(t_3505));
half_adder u0_1305(.a(t_3261), .b(t_3260), .o(t_3506), .cout(t_3507));
half_adder u0_1306(.a(t_3263), .b(t_3262), .o(t_3508), .cout(t_3509));
half_adder u0_1307(.a(t_3265), .b(t_3264), .o(t_3510), .cout(t_3511));
half_adder u0_1308(.a(t_3267), .b(t_3266), .o(t_3512), .cout(t_3513));
half_adder u0_1309(.a(t_3269), .b(t_3268), .o(t_3514), .cout(t_3515));
half_adder u0_1310(.a(t_3271), .b(t_3270), .o(t_3516), .cout(t_3517));
half_adder u0_1311(.a(t_3273), .b(t_3272), .o(t_3518), .cout(t_3519));
half_adder u0_1312(.a(t_3275), .b(t_3274), .o(t_3520), .cout(t_3521));
half_adder u0_1313(.a(t_3277), .b(t_3276), .o(t_3522), .cout(t_3523));
half_adder u0_1314(.a(t_3279), .b(t_3278), .o(t_3524), .cout(t_3525));
half_adder u0_1315(.a(t_3281), .b(t_3280), .o(t_3526), .cout(t_3527));
half_adder u0_1316(.a(t_3283), .b(t_3282), .o(t_3528), .cout(t_3529));
half_adder u0_1317(.a(t_3285), .b(t_3284), .o(t_3530), .cout(t_3531));
half_adder u0_1318(.a(t_3287), .b(t_3286), .o(t_3532), .cout());

/* Output nets Compression result */
assign compress_a = {
  t_3531,  t_3529,  t_3527,  t_3525,
  t_3523,  t_3521,  t_3519,  t_3517,
  t_3515,  t_3513,  t_3511,  t_3509,
  t_3507,  t_3505,  t_3503,  t_3501,
  t_3499,  t_3497,  t_3495,  t_3493,
  t_3491,  t_3489,  t_3487,  t_3485,
  t_3483,  t_3481,  t_3479,  t_3477,
  t_3475,  t_3473,  t_3471,  t_3469,
  t_3467,  t_3465,  t_3463,  t_3461,
  t_3459,  t_3457,  t_3455,  t_3453,
  t_3451,  t_3449,  t_3447,  t_3445,
  t_3443,  t_3441,  t_3439,  t_3437,
  t_3435,  t_3433,  t_3431,  t_3429,
  t_3427,  t_3425,  t_3423,  t_3421,
  t_3419,  t_3417,  t_3415,  t_3413,
  t_3411,  t_3409,  t_3407,  t_3405,
  t_3403,  t_3401,  t_3399,  t_3397,
  t_3395,  t_3393,  t_3391,  t_3389,
  t_3387,  t_3385,  t_3383,  t_3381,
  t_3379,  t_3377,  t_3375,  t_3373,
  t_3371,  t_3369,  t_3367,  t_3365,
  t_3363,  t_3361,  t_3359,  t_3357,
  t_3355,  t_3353,  t_3351,  t_3349,
  t_3347,  t_3345,  t_3343,  t_3341,
  t_3339,  t_3337,  t_3335,  t_3333,
  t_3331,  t_3329,  t_3327,  t_3325,
  t_3323,  t_3321,  t_3319,  t_3317,
  t_3315,  t_3313,  t_3311,  t_3309,
  t_3307,  t_3305,  t_3303,  t_3301,
  t_3299,  t_3297,  t_3295,  t_3293,
  t_3291,  t_3290,  t_2995,  t_3288,
  t_2993,  t_2504,  t_1631,     t_0
};
assign compress_b = {
  t_3532,  t_3530,  t_3528,  t_3526,
  t_3524,  t_3522,  t_3520,  t_3518,
  t_3516,  t_3514,  t_3512,  t_3510,
  t_3508,  t_3506,  t_3504,  t_3502,
  t_3500,  t_3498,  t_3496,  t_3494,
  t_3492,  t_3490,  t_3488,  t_3486,
  t_3484,  t_3482,  t_3480,  t_3478,
  t_3476,  t_3474,  t_3472,  t_3470,
  t_3468,  t_3466,  t_3464,  t_3462,
  t_3460,  t_3458,  t_3456,  t_3454,
  t_3452,  t_3450,  t_3448,  t_3446,
  t_3444,  t_3442,  t_3440,  t_3438,
  t_3436,  t_3434,  t_3432,  t_3430,
  t_3428,  t_3426,  t_3424,  t_3422,
  t_3420,  t_3418,  t_3416,  t_3414,
  t_3412,  t_3410,  t_3408,  t_3406,
  t_3404,  t_3402,  t_3400,  t_3398,
  t_3396,  t_3394,  t_3392,  t_3390,
  t_3388,  t_3386,  t_3384,  t_3382,
  t_3380,  t_3378,  t_3376,  t_3374,
  t_3372,  t_3370,  t_3368,  t_3366,
  t_3364,  t_3362,  t_3360,  t_3358,
  t_3356,  t_3354,  t_3352,  t_3350,
  t_3348,  t_3346,  t_3344,  t_3342,
  t_3340,  t_3338,  t_3336,  t_3334,
  t_3332,  t_3330,  t_3328,  t_3326,
  t_3324,  t_3322,  t_3320,  t_3318,
  t_3316,  t_3314,  t_3312,  t_3310,
  t_3308,  t_3306,  t_3304,  t_3302,
  t_3300,  t_3298,  t_3296,  t_3294,
  t_3292,    1'b0,  t_3289,    1'b0,
    1'b0,    1'b0,    1'b0,    1'b0
};

endmodule

/********************************************************************************/

module _128_wallace_tree(
//inputs
	partial_products,
	carry,
//outputs
	compress_a,
	compress_b
);

localparam width = 128;

input wire [(width+2)*(width/2+1)-1:0] partial_products;
input wire [width/2-1:0] carry;
output wire [2*width-1:0] compress_a;
output wire [2*width-1:0] compress_b;

/* Input nets */
wire    s_0_0,    s_0_1,    s_1_0,    s_2_0,    s_2_1,    s_2_2;
wire    s_3_0,    s_3_1,    s_4_0,    s_4_1,    s_4_2,    s_4_3;
wire    s_5_0,    s_5_1,    s_5_2,    s_6_0,    s_6_1,    s_6_2;
wire    s_6_3,    s_6_4,    s_7_0,    s_7_1,    s_7_2,    s_7_3;
wire    s_8_0,    s_8_1,    s_8_2,    s_8_3,    s_8_4,    s_8_5;
wire    s_9_0,    s_9_1,    s_9_2,    s_9_3,    s_9_4,   s_10_0;
wire   s_10_1,   s_10_2,   s_10_3,   s_10_4,   s_10_5,   s_10_6;
wire   s_11_0,   s_11_1,   s_11_2,   s_11_3,   s_11_4,   s_11_5;
wire   s_12_0,   s_12_1,   s_12_2,   s_12_3,   s_12_4,   s_12_5;
wire   s_12_6,   s_12_7,   s_13_0,   s_13_1,   s_13_2,   s_13_3;
wire   s_13_4,   s_13_5,   s_13_6,   s_14_0,   s_14_1,   s_14_2;
wire   s_14_3,   s_14_4,   s_14_5,   s_14_6,   s_14_7,   s_14_8;
wire   s_15_0,   s_15_1,   s_15_2,   s_15_3,   s_15_4,   s_15_5;
wire   s_15_6,   s_15_7,   s_16_0,   s_16_1,   s_16_2,   s_16_3;
wire   s_16_4,   s_16_5,   s_16_6,   s_16_7,   s_16_8,   s_16_9;
wire   s_17_0,   s_17_1,   s_17_2,   s_17_3,   s_17_4,   s_17_5;
wire   s_17_6,   s_17_7,   s_17_8,   s_18_0,   s_18_1,   s_18_2;
wire   s_18_3,   s_18_4,   s_18_5,   s_18_6,   s_18_7,   s_18_8;
wire   s_18_9,  s_18_10,   s_19_0,   s_19_1,   s_19_2,   s_19_3;
wire   s_19_4,   s_19_5,   s_19_6,   s_19_7,   s_19_8,   s_19_9;
wire   s_20_0,   s_20_1,   s_20_2,   s_20_3,   s_20_4,   s_20_5;
wire   s_20_6,   s_20_7,   s_20_8,   s_20_9,  s_20_10,  s_20_11;
wire   s_21_0,   s_21_1,   s_21_2,   s_21_3,   s_21_4,   s_21_5;
wire   s_21_6,   s_21_7,   s_21_8,   s_21_9,  s_21_10,   s_22_0;
wire   s_22_1,   s_22_2,   s_22_3,   s_22_4,   s_22_5,   s_22_6;
wire   s_22_7,   s_22_8,   s_22_9,  s_22_10,  s_22_11,  s_22_12;
wire   s_23_0,   s_23_1,   s_23_2,   s_23_3,   s_23_4,   s_23_5;
wire   s_23_6,   s_23_7,   s_23_8,   s_23_9,  s_23_10,  s_23_11;
wire   s_24_0,   s_24_1,   s_24_2,   s_24_3,   s_24_4,   s_24_5;
wire   s_24_6,   s_24_7,   s_24_8,   s_24_9,  s_24_10,  s_24_11;
wire  s_24_12,  s_24_13,   s_25_0,   s_25_1,   s_25_2,   s_25_3;
wire   s_25_4,   s_25_5,   s_25_6,   s_25_7,   s_25_8,   s_25_9;
wire  s_25_10,  s_25_11,  s_25_12,   s_26_0,   s_26_1,   s_26_2;
wire   s_26_3,   s_26_4,   s_26_5,   s_26_6,   s_26_7,   s_26_8;
wire   s_26_9,  s_26_10,  s_26_11,  s_26_12,  s_26_13,  s_26_14;
wire   s_27_0,   s_27_1,   s_27_2,   s_27_3,   s_27_4,   s_27_5;
wire   s_27_6,   s_27_7,   s_27_8,   s_27_9,  s_27_10,  s_27_11;
wire  s_27_12,  s_27_13,   s_28_0,   s_28_1,   s_28_2,   s_28_3;
wire   s_28_4,   s_28_5,   s_28_6,   s_28_7,   s_28_8,   s_28_9;
wire  s_28_10,  s_28_11,  s_28_12,  s_28_13,  s_28_14,  s_28_15;
wire   s_29_0,   s_29_1,   s_29_2,   s_29_3,   s_29_4,   s_29_5;
wire   s_29_6,   s_29_7,   s_29_8,   s_29_9,  s_29_10,  s_29_11;
wire  s_29_12,  s_29_13,  s_29_14,   s_30_0,   s_30_1,   s_30_2;
wire   s_30_3,   s_30_4,   s_30_5,   s_30_6,   s_30_7,   s_30_8;
wire   s_30_9,  s_30_10,  s_30_11,  s_30_12,  s_30_13,  s_30_14;
wire  s_30_15,  s_30_16,   s_31_0,   s_31_1,   s_31_2,   s_31_3;
wire   s_31_4,   s_31_5,   s_31_6,   s_31_7,   s_31_8,   s_31_9;
wire  s_31_10,  s_31_11,  s_31_12,  s_31_13,  s_31_14,  s_31_15;
wire   s_32_0,   s_32_1,   s_32_2,   s_32_3,   s_32_4,   s_32_5;
wire   s_32_6,   s_32_7,   s_32_8,   s_32_9,  s_32_10,  s_32_11;
wire  s_32_12,  s_32_13,  s_32_14,  s_32_15,  s_32_16,  s_32_17;
wire   s_33_0,   s_33_1,   s_33_2,   s_33_3,   s_33_4,   s_33_5;
wire   s_33_6,   s_33_7,   s_33_8,   s_33_9,  s_33_10,  s_33_11;
wire  s_33_12,  s_33_13,  s_33_14,  s_33_15,  s_33_16,   s_34_0;
wire   s_34_1,   s_34_2,   s_34_3,   s_34_4,   s_34_5,   s_34_6;
wire   s_34_7,   s_34_8,   s_34_9,  s_34_10,  s_34_11,  s_34_12;
wire  s_34_13,  s_34_14,  s_34_15,  s_34_16,  s_34_17,  s_34_18;
wire   s_35_0,   s_35_1,   s_35_2,   s_35_3,   s_35_4,   s_35_5;
wire   s_35_6,   s_35_7,   s_35_8,   s_35_9,  s_35_10,  s_35_11;
wire  s_35_12,  s_35_13,  s_35_14,  s_35_15,  s_35_16,  s_35_17;
wire   s_36_0,   s_36_1,   s_36_2,   s_36_3,   s_36_4,   s_36_5;
wire   s_36_6,   s_36_7,   s_36_8,   s_36_9,  s_36_10,  s_36_11;
wire  s_36_12,  s_36_13,  s_36_14,  s_36_15,  s_36_16,  s_36_17;
wire  s_36_18,  s_36_19,   s_37_0,   s_37_1,   s_37_2,   s_37_3;
wire   s_37_4,   s_37_5,   s_37_6,   s_37_7,   s_37_8,   s_37_9;
wire  s_37_10,  s_37_11,  s_37_12,  s_37_13,  s_37_14,  s_37_15;
wire  s_37_16,  s_37_17,  s_37_18,   s_38_0,   s_38_1,   s_38_2;
wire   s_38_3,   s_38_4,   s_38_5,   s_38_6,   s_38_7,   s_38_8;
wire   s_38_9,  s_38_10,  s_38_11,  s_38_12,  s_38_13,  s_38_14;
wire  s_38_15,  s_38_16,  s_38_17,  s_38_18,  s_38_19,  s_38_20;
wire   s_39_0,   s_39_1,   s_39_2,   s_39_3,   s_39_4,   s_39_5;
wire   s_39_6,   s_39_7,   s_39_8,   s_39_9,  s_39_10,  s_39_11;
wire  s_39_12,  s_39_13,  s_39_14,  s_39_15,  s_39_16,  s_39_17;
wire  s_39_18,  s_39_19,   s_40_0,   s_40_1,   s_40_2,   s_40_3;
wire   s_40_4,   s_40_5,   s_40_6,   s_40_7,   s_40_8,   s_40_9;
wire  s_40_10,  s_40_11,  s_40_12,  s_40_13,  s_40_14,  s_40_15;
wire  s_40_16,  s_40_17,  s_40_18,  s_40_19,  s_40_20,  s_40_21;
wire   s_41_0,   s_41_1,   s_41_2,   s_41_3,   s_41_4,   s_41_5;
wire   s_41_6,   s_41_7,   s_41_8,   s_41_9,  s_41_10,  s_41_11;
wire  s_41_12,  s_41_13,  s_41_14,  s_41_15,  s_41_16,  s_41_17;
wire  s_41_18,  s_41_19,  s_41_20,   s_42_0,   s_42_1,   s_42_2;
wire   s_42_3,   s_42_4,   s_42_5,   s_42_6,   s_42_7,   s_42_8;
wire   s_42_9,  s_42_10,  s_42_11,  s_42_12,  s_42_13,  s_42_14;
wire  s_42_15,  s_42_16,  s_42_17,  s_42_18,  s_42_19,  s_42_20;
wire  s_42_21,  s_42_22,   s_43_0,   s_43_1,   s_43_2,   s_43_3;
wire   s_43_4,   s_43_5,   s_43_6,   s_43_7,   s_43_8,   s_43_9;
wire  s_43_10,  s_43_11,  s_43_12,  s_43_13,  s_43_14,  s_43_15;
wire  s_43_16,  s_43_17,  s_43_18,  s_43_19,  s_43_20,  s_43_21;
wire   s_44_0,   s_44_1,   s_44_2,   s_44_3,   s_44_4,   s_44_5;
wire   s_44_6,   s_44_7,   s_44_8,   s_44_9,  s_44_10,  s_44_11;
wire  s_44_12,  s_44_13,  s_44_14,  s_44_15,  s_44_16,  s_44_17;
wire  s_44_18,  s_44_19,  s_44_20,  s_44_21,  s_44_22,  s_44_23;
wire   s_45_0,   s_45_1,   s_45_2,   s_45_3,   s_45_4,   s_45_5;
wire   s_45_6,   s_45_7,   s_45_8,   s_45_9,  s_45_10,  s_45_11;
wire  s_45_12,  s_45_13,  s_45_14,  s_45_15,  s_45_16,  s_45_17;
wire  s_45_18,  s_45_19,  s_45_20,  s_45_21,  s_45_22,   s_46_0;
wire   s_46_1,   s_46_2,   s_46_3,   s_46_4,   s_46_5,   s_46_6;
wire   s_46_7,   s_46_8,   s_46_9,  s_46_10,  s_46_11,  s_46_12;
wire  s_46_13,  s_46_14,  s_46_15,  s_46_16,  s_46_17,  s_46_18;
wire  s_46_19,  s_46_20,  s_46_21,  s_46_22,  s_46_23,  s_46_24;
wire   s_47_0,   s_47_1,   s_47_2,   s_47_3,   s_47_4,   s_47_5;
wire   s_47_6,   s_47_7,   s_47_8,   s_47_9,  s_47_10,  s_47_11;
wire  s_47_12,  s_47_13,  s_47_14,  s_47_15,  s_47_16,  s_47_17;
wire  s_47_18,  s_47_19,  s_47_20,  s_47_21,  s_47_22,  s_47_23;
wire   s_48_0,   s_48_1,   s_48_2,   s_48_3,   s_48_4,   s_48_5;
wire   s_48_6,   s_48_7,   s_48_8,   s_48_9,  s_48_10,  s_48_11;
wire  s_48_12,  s_48_13,  s_48_14,  s_48_15,  s_48_16,  s_48_17;
wire  s_48_18,  s_48_19,  s_48_20,  s_48_21,  s_48_22,  s_48_23;
wire  s_48_24,  s_48_25,   s_49_0,   s_49_1,   s_49_2,   s_49_3;
wire   s_49_4,   s_49_5,   s_49_6,   s_49_7,   s_49_8,   s_49_9;
wire  s_49_10,  s_49_11,  s_49_12,  s_49_13,  s_49_14,  s_49_15;
wire  s_49_16,  s_49_17,  s_49_18,  s_49_19,  s_49_20,  s_49_21;
wire  s_49_22,  s_49_23,  s_49_24,   s_50_0,   s_50_1,   s_50_2;
wire   s_50_3,   s_50_4,   s_50_5,   s_50_6,   s_50_7,   s_50_8;
wire   s_50_9,  s_50_10,  s_50_11,  s_50_12,  s_50_13,  s_50_14;
wire  s_50_15,  s_50_16,  s_50_17,  s_50_18,  s_50_19,  s_50_20;
wire  s_50_21,  s_50_22,  s_50_23,  s_50_24,  s_50_25,  s_50_26;
wire   s_51_0,   s_51_1,   s_51_2,   s_51_3,   s_51_4,   s_51_5;
wire   s_51_6,   s_51_7,   s_51_8,   s_51_9,  s_51_10,  s_51_11;
wire  s_51_12,  s_51_13,  s_51_14,  s_51_15,  s_51_16,  s_51_17;
wire  s_51_18,  s_51_19,  s_51_20,  s_51_21,  s_51_22,  s_51_23;
wire  s_51_24,  s_51_25,   s_52_0,   s_52_1,   s_52_2,   s_52_3;
wire   s_52_4,   s_52_5,   s_52_6,   s_52_7,   s_52_8,   s_52_9;
wire  s_52_10,  s_52_11,  s_52_12,  s_52_13,  s_52_14,  s_52_15;
wire  s_52_16,  s_52_17,  s_52_18,  s_52_19,  s_52_20,  s_52_21;
wire  s_52_22,  s_52_23,  s_52_24,  s_52_25,  s_52_26,  s_52_27;
wire   s_53_0,   s_53_1,   s_53_2,   s_53_3,   s_53_4,   s_53_5;
wire   s_53_6,   s_53_7,   s_53_8,   s_53_9,  s_53_10,  s_53_11;
wire  s_53_12,  s_53_13,  s_53_14,  s_53_15,  s_53_16,  s_53_17;
wire  s_53_18,  s_53_19,  s_53_20,  s_53_21,  s_53_22,  s_53_23;
wire  s_53_24,  s_53_25,  s_53_26,   s_54_0,   s_54_1,   s_54_2;
wire   s_54_3,   s_54_4,   s_54_5,   s_54_6,   s_54_7,   s_54_8;
wire   s_54_9,  s_54_10,  s_54_11,  s_54_12,  s_54_13,  s_54_14;
wire  s_54_15,  s_54_16,  s_54_17,  s_54_18,  s_54_19,  s_54_20;
wire  s_54_21,  s_54_22,  s_54_23,  s_54_24,  s_54_25,  s_54_26;
wire  s_54_27,  s_54_28,   s_55_0,   s_55_1,   s_55_2,   s_55_3;
wire   s_55_4,   s_55_5,   s_55_6,   s_55_7,   s_55_8,   s_55_9;
wire  s_55_10,  s_55_11,  s_55_12,  s_55_13,  s_55_14,  s_55_15;
wire  s_55_16,  s_55_17,  s_55_18,  s_55_19,  s_55_20,  s_55_21;
wire  s_55_22,  s_55_23,  s_55_24,  s_55_25,  s_55_26,  s_55_27;
wire   s_56_0,   s_56_1,   s_56_2,   s_56_3,   s_56_4,   s_56_5;
wire   s_56_6,   s_56_7,   s_56_8,   s_56_9,  s_56_10,  s_56_11;
wire  s_56_12,  s_56_13,  s_56_14,  s_56_15,  s_56_16,  s_56_17;
wire  s_56_18,  s_56_19,  s_56_20,  s_56_21,  s_56_22,  s_56_23;
wire  s_56_24,  s_56_25,  s_56_26,  s_56_27,  s_56_28,  s_56_29;
wire   s_57_0,   s_57_1,   s_57_2,   s_57_3,   s_57_4,   s_57_5;
wire   s_57_6,   s_57_7,   s_57_8,   s_57_9,  s_57_10,  s_57_11;
wire  s_57_12,  s_57_13,  s_57_14,  s_57_15,  s_57_16,  s_57_17;
wire  s_57_18,  s_57_19,  s_57_20,  s_57_21,  s_57_22,  s_57_23;
wire  s_57_24,  s_57_25,  s_57_26,  s_57_27,  s_57_28,   s_58_0;
wire   s_58_1,   s_58_2,   s_58_3,   s_58_4,   s_58_5,   s_58_6;
wire   s_58_7,   s_58_8,   s_58_9,  s_58_10,  s_58_11,  s_58_12;
wire  s_58_13,  s_58_14,  s_58_15,  s_58_16,  s_58_17,  s_58_18;
wire  s_58_19,  s_58_20,  s_58_21,  s_58_22,  s_58_23,  s_58_24;
wire  s_58_25,  s_58_26,  s_58_27,  s_58_28,  s_58_29,  s_58_30;
wire   s_59_0,   s_59_1,   s_59_2,   s_59_3,   s_59_4,   s_59_5;
wire   s_59_6,   s_59_7,   s_59_8,   s_59_9,  s_59_10,  s_59_11;
wire  s_59_12,  s_59_13,  s_59_14,  s_59_15,  s_59_16,  s_59_17;
wire  s_59_18,  s_59_19,  s_59_20,  s_59_21,  s_59_22,  s_59_23;
wire  s_59_24,  s_59_25,  s_59_26,  s_59_27,  s_59_28,  s_59_29;
wire   s_60_0,   s_60_1,   s_60_2,   s_60_3,   s_60_4,   s_60_5;
wire   s_60_6,   s_60_7,   s_60_8,   s_60_9,  s_60_10,  s_60_11;
wire  s_60_12,  s_60_13,  s_60_14,  s_60_15,  s_60_16,  s_60_17;
wire  s_60_18,  s_60_19,  s_60_20,  s_60_21,  s_60_22,  s_60_23;
wire  s_60_24,  s_60_25,  s_60_26,  s_60_27,  s_60_28,  s_60_29;
wire  s_60_30,  s_60_31,   s_61_0,   s_61_1,   s_61_2,   s_61_3;
wire   s_61_4,   s_61_5,   s_61_6,   s_61_7,   s_61_8,   s_61_9;
wire  s_61_10,  s_61_11,  s_61_12,  s_61_13,  s_61_14,  s_61_15;
wire  s_61_16,  s_61_17,  s_61_18,  s_61_19,  s_61_20,  s_61_21;
wire  s_61_22,  s_61_23,  s_61_24,  s_61_25,  s_61_26,  s_61_27;
wire  s_61_28,  s_61_29,  s_61_30,   s_62_0,   s_62_1,   s_62_2;
wire   s_62_3,   s_62_4,   s_62_5,   s_62_6,   s_62_7,   s_62_8;
wire   s_62_9,  s_62_10,  s_62_11,  s_62_12,  s_62_13,  s_62_14;
wire  s_62_15,  s_62_16,  s_62_17,  s_62_18,  s_62_19,  s_62_20;
wire  s_62_21,  s_62_22,  s_62_23,  s_62_24,  s_62_25,  s_62_26;
wire  s_62_27,  s_62_28,  s_62_29,  s_62_30,  s_62_31,  s_62_32;
wire   s_63_0,   s_63_1,   s_63_2,   s_63_3,   s_63_4,   s_63_5;
wire   s_63_6,   s_63_7,   s_63_8,   s_63_9,  s_63_10,  s_63_11;
wire  s_63_12,  s_63_13,  s_63_14,  s_63_15,  s_63_16,  s_63_17;
wire  s_63_18,  s_63_19,  s_63_20,  s_63_21,  s_63_22,  s_63_23;
wire  s_63_24,  s_63_25,  s_63_26,  s_63_27,  s_63_28,  s_63_29;
wire  s_63_30,  s_63_31,   s_64_0,   s_64_1,   s_64_2,   s_64_3;
wire   s_64_4,   s_64_5,   s_64_6,   s_64_7,   s_64_8,   s_64_9;
wire  s_64_10,  s_64_11,  s_64_12,  s_64_13,  s_64_14,  s_64_15;
wire  s_64_16,  s_64_17,  s_64_18,  s_64_19,  s_64_20,  s_64_21;
wire  s_64_22,  s_64_23,  s_64_24,  s_64_25,  s_64_26,  s_64_27;
wire  s_64_28,  s_64_29,  s_64_30,  s_64_31,  s_64_32,  s_64_33;
wire   s_65_0,   s_65_1,   s_65_2,   s_65_3,   s_65_4,   s_65_5;
wire   s_65_6,   s_65_7,   s_65_8,   s_65_9,  s_65_10,  s_65_11;
wire  s_65_12,  s_65_13,  s_65_14,  s_65_15,  s_65_16,  s_65_17;
wire  s_65_18,  s_65_19,  s_65_20,  s_65_21,  s_65_22,  s_65_23;
wire  s_65_24,  s_65_25,  s_65_26,  s_65_27,  s_65_28,  s_65_29;
wire  s_65_30,  s_65_31,  s_65_32,   s_66_0,   s_66_1,   s_66_2;
wire   s_66_3,   s_66_4,   s_66_5,   s_66_6,   s_66_7,   s_66_8;
wire   s_66_9,  s_66_10,  s_66_11,  s_66_12,  s_66_13,  s_66_14;
wire  s_66_15,  s_66_16,  s_66_17,  s_66_18,  s_66_19,  s_66_20;
wire  s_66_21,  s_66_22,  s_66_23,  s_66_24,  s_66_25,  s_66_26;
wire  s_66_27,  s_66_28,  s_66_29,  s_66_30,  s_66_31,  s_66_32;
wire  s_66_33,  s_66_34,   s_67_0,   s_67_1,   s_67_2,   s_67_3;
wire   s_67_4,   s_67_5,   s_67_6,   s_67_7,   s_67_8,   s_67_9;
wire  s_67_10,  s_67_11,  s_67_12,  s_67_13,  s_67_14,  s_67_15;
wire  s_67_16,  s_67_17,  s_67_18,  s_67_19,  s_67_20,  s_67_21;
wire  s_67_22,  s_67_23,  s_67_24,  s_67_25,  s_67_26,  s_67_27;
wire  s_67_28,  s_67_29,  s_67_30,  s_67_31,  s_67_32,  s_67_33;
wire   s_68_0,   s_68_1,   s_68_2,   s_68_3,   s_68_4,   s_68_5;
wire   s_68_6,   s_68_7,   s_68_8,   s_68_9,  s_68_10,  s_68_11;
wire  s_68_12,  s_68_13,  s_68_14,  s_68_15,  s_68_16,  s_68_17;
wire  s_68_18,  s_68_19,  s_68_20,  s_68_21,  s_68_22,  s_68_23;
wire  s_68_24,  s_68_25,  s_68_26,  s_68_27,  s_68_28,  s_68_29;
wire  s_68_30,  s_68_31,  s_68_32,  s_68_33,  s_68_34,  s_68_35;
wire   s_69_0,   s_69_1,   s_69_2,   s_69_3,   s_69_4,   s_69_5;
wire   s_69_6,   s_69_7,   s_69_8,   s_69_9,  s_69_10,  s_69_11;
wire  s_69_12,  s_69_13,  s_69_14,  s_69_15,  s_69_16,  s_69_17;
wire  s_69_18,  s_69_19,  s_69_20,  s_69_21,  s_69_22,  s_69_23;
wire  s_69_24,  s_69_25,  s_69_26,  s_69_27,  s_69_28,  s_69_29;
wire  s_69_30,  s_69_31,  s_69_32,  s_69_33,  s_69_34,   s_70_0;
wire   s_70_1,   s_70_2,   s_70_3,   s_70_4,   s_70_5,   s_70_6;
wire   s_70_7,   s_70_8,   s_70_9,  s_70_10,  s_70_11,  s_70_12;
wire  s_70_13,  s_70_14,  s_70_15,  s_70_16,  s_70_17,  s_70_18;
wire  s_70_19,  s_70_20,  s_70_21,  s_70_22,  s_70_23,  s_70_24;
wire  s_70_25,  s_70_26,  s_70_27,  s_70_28,  s_70_29,  s_70_30;
wire  s_70_31,  s_70_32,  s_70_33,  s_70_34,  s_70_35,  s_70_36;
wire   s_71_0,   s_71_1,   s_71_2,   s_71_3,   s_71_4,   s_71_5;
wire   s_71_6,   s_71_7,   s_71_8,   s_71_9,  s_71_10,  s_71_11;
wire  s_71_12,  s_71_13,  s_71_14,  s_71_15,  s_71_16,  s_71_17;
wire  s_71_18,  s_71_19,  s_71_20,  s_71_21,  s_71_22,  s_71_23;
wire  s_71_24,  s_71_25,  s_71_26,  s_71_27,  s_71_28,  s_71_29;
wire  s_71_30,  s_71_31,  s_71_32,  s_71_33,  s_71_34,  s_71_35;
wire   s_72_0,   s_72_1,   s_72_2,   s_72_3,   s_72_4,   s_72_5;
wire   s_72_6,   s_72_7,   s_72_8,   s_72_9,  s_72_10,  s_72_11;
wire  s_72_12,  s_72_13,  s_72_14,  s_72_15,  s_72_16,  s_72_17;
wire  s_72_18,  s_72_19,  s_72_20,  s_72_21,  s_72_22,  s_72_23;
wire  s_72_24,  s_72_25,  s_72_26,  s_72_27,  s_72_28,  s_72_29;
wire  s_72_30,  s_72_31,  s_72_32,  s_72_33,  s_72_34,  s_72_35;
wire  s_72_36,  s_72_37,   s_73_0,   s_73_1,   s_73_2,   s_73_3;
wire   s_73_4,   s_73_5,   s_73_6,   s_73_7,   s_73_8,   s_73_9;
wire  s_73_10,  s_73_11,  s_73_12,  s_73_13,  s_73_14,  s_73_15;
wire  s_73_16,  s_73_17,  s_73_18,  s_73_19,  s_73_20,  s_73_21;
wire  s_73_22,  s_73_23,  s_73_24,  s_73_25,  s_73_26,  s_73_27;
wire  s_73_28,  s_73_29,  s_73_30,  s_73_31,  s_73_32,  s_73_33;
wire  s_73_34,  s_73_35,  s_73_36,   s_74_0,   s_74_1,   s_74_2;
wire   s_74_3,   s_74_4,   s_74_5,   s_74_6,   s_74_7,   s_74_8;
wire   s_74_9,  s_74_10,  s_74_11,  s_74_12,  s_74_13,  s_74_14;
wire  s_74_15,  s_74_16,  s_74_17,  s_74_18,  s_74_19,  s_74_20;
wire  s_74_21,  s_74_22,  s_74_23,  s_74_24,  s_74_25,  s_74_26;
wire  s_74_27,  s_74_28,  s_74_29,  s_74_30,  s_74_31,  s_74_32;
wire  s_74_33,  s_74_34,  s_74_35,  s_74_36,  s_74_37,  s_74_38;
wire   s_75_0,   s_75_1,   s_75_2,   s_75_3,   s_75_4,   s_75_5;
wire   s_75_6,   s_75_7,   s_75_8,   s_75_9,  s_75_10,  s_75_11;
wire  s_75_12,  s_75_13,  s_75_14,  s_75_15,  s_75_16,  s_75_17;
wire  s_75_18,  s_75_19,  s_75_20,  s_75_21,  s_75_22,  s_75_23;
wire  s_75_24,  s_75_25,  s_75_26,  s_75_27,  s_75_28,  s_75_29;
wire  s_75_30,  s_75_31,  s_75_32,  s_75_33,  s_75_34,  s_75_35;
wire  s_75_36,  s_75_37,   s_76_0,   s_76_1,   s_76_2,   s_76_3;
wire   s_76_4,   s_76_5,   s_76_6,   s_76_7,   s_76_8,   s_76_9;
wire  s_76_10,  s_76_11,  s_76_12,  s_76_13,  s_76_14,  s_76_15;
wire  s_76_16,  s_76_17,  s_76_18,  s_76_19,  s_76_20,  s_76_21;
wire  s_76_22,  s_76_23,  s_76_24,  s_76_25,  s_76_26,  s_76_27;
wire  s_76_28,  s_76_29,  s_76_30,  s_76_31,  s_76_32,  s_76_33;
wire  s_76_34,  s_76_35,  s_76_36,  s_76_37,  s_76_38,  s_76_39;
wire   s_77_0,   s_77_1,   s_77_2,   s_77_3,   s_77_4,   s_77_5;
wire   s_77_6,   s_77_7,   s_77_8,   s_77_9,  s_77_10,  s_77_11;
wire  s_77_12,  s_77_13,  s_77_14,  s_77_15,  s_77_16,  s_77_17;
wire  s_77_18,  s_77_19,  s_77_20,  s_77_21,  s_77_22,  s_77_23;
wire  s_77_24,  s_77_25,  s_77_26,  s_77_27,  s_77_28,  s_77_29;
wire  s_77_30,  s_77_31,  s_77_32,  s_77_33,  s_77_34,  s_77_35;
wire  s_77_36,  s_77_37,  s_77_38,   s_78_0,   s_78_1,   s_78_2;
wire   s_78_3,   s_78_4,   s_78_5,   s_78_6,   s_78_7,   s_78_8;
wire   s_78_9,  s_78_10,  s_78_11,  s_78_12,  s_78_13,  s_78_14;
wire  s_78_15,  s_78_16,  s_78_17,  s_78_18,  s_78_19,  s_78_20;
wire  s_78_21,  s_78_22,  s_78_23,  s_78_24,  s_78_25,  s_78_26;
wire  s_78_27,  s_78_28,  s_78_29,  s_78_30,  s_78_31,  s_78_32;
wire  s_78_33,  s_78_34,  s_78_35,  s_78_36,  s_78_37,  s_78_38;
wire  s_78_39,  s_78_40,   s_79_0,   s_79_1,   s_79_2,   s_79_3;
wire   s_79_4,   s_79_5,   s_79_6,   s_79_7,   s_79_8,   s_79_9;
wire  s_79_10,  s_79_11,  s_79_12,  s_79_13,  s_79_14,  s_79_15;
wire  s_79_16,  s_79_17,  s_79_18,  s_79_19,  s_79_20,  s_79_21;
wire  s_79_22,  s_79_23,  s_79_24,  s_79_25,  s_79_26,  s_79_27;
wire  s_79_28,  s_79_29,  s_79_30,  s_79_31,  s_79_32,  s_79_33;
wire  s_79_34,  s_79_35,  s_79_36,  s_79_37,  s_79_38,  s_79_39;
wire   s_80_0,   s_80_1,   s_80_2,   s_80_3,   s_80_4,   s_80_5;
wire   s_80_6,   s_80_7,   s_80_8,   s_80_9,  s_80_10,  s_80_11;
wire  s_80_12,  s_80_13,  s_80_14,  s_80_15,  s_80_16,  s_80_17;
wire  s_80_18,  s_80_19,  s_80_20,  s_80_21,  s_80_22,  s_80_23;
wire  s_80_24,  s_80_25,  s_80_26,  s_80_27,  s_80_28,  s_80_29;
wire  s_80_30,  s_80_31,  s_80_32,  s_80_33,  s_80_34,  s_80_35;
wire  s_80_36,  s_80_37,  s_80_38,  s_80_39,  s_80_40,  s_80_41;
wire   s_81_0,   s_81_1,   s_81_2,   s_81_3,   s_81_4,   s_81_5;
wire   s_81_6,   s_81_7,   s_81_8,   s_81_9,  s_81_10,  s_81_11;
wire  s_81_12,  s_81_13,  s_81_14,  s_81_15,  s_81_16,  s_81_17;
wire  s_81_18,  s_81_19,  s_81_20,  s_81_21,  s_81_22,  s_81_23;
wire  s_81_24,  s_81_25,  s_81_26,  s_81_27,  s_81_28,  s_81_29;
wire  s_81_30,  s_81_31,  s_81_32,  s_81_33,  s_81_34,  s_81_35;
wire  s_81_36,  s_81_37,  s_81_38,  s_81_39,  s_81_40,   s_82_0;
wire   s_82_1,   s_82_2,   s_82_3,   s_82_4,   s_82_5,   s_82_6;
wire   s_82_7,   s_82_8,   s_82_9,  s_82_10,  s_82_11,  s_82_12;
wire  s_82_13,  s_82_14,  s_82_15,  s_82_16,  s_82_17,  s_82_18;
wire  s_82_19,  s_82_20,  s_82_21,  s_82_22,  s_82_23,  s_82_24;
wire  s_82_25,  s_82_26,  s_82_27,  s_82_28,  s_82_29,  s_82_30;
wire  s_82_31,  s_82_32,  s_82_33,  s_82_34,  s_82_35,  s_82_36;
wire  s_82_37,  s_82_38,  s_82_39,  s_82_40,  s_82_41,  s_82_42;
wire   s_83_0,   s_83_1,   s_83_2,   s_83_3,   s_83_4,   s_83_5;
wire   s_83_6,   s_83_7,   s_83_8,   s_83_9,  s_83_10,  s_83_11;
wire  s_83_12,  s_83_13,  s_83_14,  s_83_15,  s_83_16,  s_83_17;
wire  s_83_18,  s_83_19,  s_83_20,  s_83_21,  s_83_22,  s_83_23;
wire  s_83_24,  s_83_25,  s_83_26,  s_83_27,  s_83_28,  s_83_29;
wire  s_83_30,  s_83_31,  s_83_32,  s_83_33,  s_83_34,  s_83_35;
wire  s_83_36,  s_83_37,  s_83_38,  s_83_39,  s_83_40,  s_83_41;
wire   s_84_0,   s_84_1,   s_84_2,   s_84_3,   s_84_4,   s_84_5;
wire   s_84_6,   s_84_7,   s_84_8,   s_84_9,  s_84_10,  s_84_11;
wire  s_84_12,  s_84_13,  s_84_14,  s_84_15,  s_84_16,  s_84_17;
wire  s_84_18,  s_84_19,  s_84_20,  s_84_21,  s_84_22,  s_84_23;
wire  s_84_24,  s_84_25,  s_84_26,  s_84_27,  s_84_28,  s_84_29;
wire  s_84_30,  s_84_31,  s_84_32,  s_84_33,  s_84_34,  s_84_35;
wire  s_84_36,  s_84_37,  s_84_38,  s_84_39,  s_84_40,  s_84_41;
wire  s_84_42,  s_84_43,   s_85_0,   s_85_1,   s_85_2,   s_85_3;
wire   s_85_4,   s_85_5,   s_85_6,   s_85_7,   s_85_8,   s_85_9;
wire  s_85_10,  s_85_11,  s_85_12,  s_85_13,  s_85_14,  s_85_15;
wire  s_85_16,  s_85_17,  s_85_18,  s_85_19,  s_85_20,  s_85_21;
wire  s_85_22,  s_85_23,  s_85_24,  s_85_25,  s_85_26,  s_85_27;
wire  s_85_28,  s_85_29,  s_85_30,  s_85_31,  s_85_32,  s_85_33;
wire  s_85_34,  s_85_35,  s_85_36,  s_85_37,  s_85_38,  s_85_39;
wire  s_85_40,  s_85_41,  s_85_42,   s_86_0,   s_86_1,   s_86_2;
wire   s_86_3,   s_86_4,   s_86_5,   s_86_6,   s_86_7,   s_86_8;
wire   s_86_9,  s_86_10,  s_86_11,  s_86_12,  s_86_13,  s_86_14;
wire  s_86_15,  s_86_16,  s_86_17,  s_86_18,  s_86_19,  s_86_20;
wire  s_86_21,  s_86_22,  s_86_23,  s_86_24,  s_86_25,  s_86_26;
wire  s_86_27,  s_86_28,  s_86_29,  s_86_30,  s_86_31,  s_86_32;
wire  s_86_33,  s_86_34,  s_86_35,  s_86_36,  s_86_37,  s_86_38;
wire  s_86_39,  s_86_40,  s_86_41,  s_86_42,  s_86_43,  s_86_44;
wire   s_87_0,   s_87_1,   s_87_2,   s_87_3,   s_87_4,   s_87_5;
wire   s_87_6,   s_87_7,   s_87_8,   s_87_9,  s_87_10,  s_87_11;
wire  s_87_12,  s_87_13,  s_87_14,  s_87_15,  s_87_16,  s_87_17;
wire  s_87_18,  s_87_19,  s_87_20,  s_87_21,  s_87_22,  s_87_23;
wire  s_87_24,  s_87_25,  s_87_26,  s_87_27,  s_87_28,  s_87_29;
wire  s_87_30,  s_87_31,  s_87_32,  s_87_33,  s_87_34,  s_87_35;
wire  s_87_36,  s_87_37,  s_87_38,  s_87_39,  s_87_40,  s_87_41;
wire  s_87_42,  s_87_43,   s_88_0,   s_88_1,   s_88_2,   s_88_3;
wire   s_88_4,   s_88_5,   s_88_6,   s_88_7,   s_88_8,   s_88_9;
wire  s_88_10,  s_88_11,  s_88_12,  s_88_13,  s_88_14,  s_88_15;
wire  s_88_16,  s_88_17,  s_88_18,  s_88_19,  s_88_20,  s_88_21;
wire  s_88_22,  s_88_23,  s_88_24,  s_88_25,  s_88_26,  s_88_27;
wire  s_88_28,  s_88_29,  s_88_30,  s_88_31,  s_88_32,  s_88_33;
wire  s_88_34,  s_88_35,  s_88_36,  s_88_37,  s_88_38,  s_88_39;
wire  s_88_40,  s_88_41,  s_88_42,  s_88_43,  s_88_44,  s_88_45;
wire   s_89_0,   s_89_1,   s_89_2,   s_89_3,   s_89_4,   s_89_5;
wire   s_89_6,   s_89_7,   s_89_8,   s_89_9,  s_89_10,  s_89_11;
wire  s_89_12,  s_89_13,  s_89_14,  s_89_15,  s_89_16,  s_89_17;
wire  s_89_18,  s_89_19,  s_89_20,  s_89_21,  s_89_22,  s_89_23;
wire  s_89_24,  s_89_25,  s_89_26,  s_89_27,  s_89_28,  s_89_29;
wire  s_89_30,  s_89_31,  s_89_32,  s_89_33,  s_89_34,  s_89_35;
wire  s_89_36,  s_89_37,  s_89_38,  s_89_39,  s_89_40,  s_89_41;
wire  s_89_42,  s_89_43,  s_89_44,   s_90_0,   s_90_1,   s_90_2;
wire   s_90_3,   s_90_4,   s_90_5,   s_90_6,   s_90_7,   s_90_8;
wire   s_90_9,  s_90_10,  s_90_11,  s_90_12,  s_90_13,  s_90_14;
wire  s_90_15,  s_90_16,  s_90_17,  s_90_18,  s_90_19,  s_90_20;
wire  s_90_21,  s_90_22,  s_90_23,  s_90_24,  s_90_25,  s_90_26;
wire  s_90_27,  s_90_28,  s_90_29,  s_90_30,  s_90_31,  s_90_32;
wire  s_90_33,  s_90_34,  s_90_35,  s_90_36,  s_90_37,  s_90_38;
wire  s_90_39,  s_90_40,  s_90_41,  s_90_42,  s_90_43,  s_90_44;
wire  s_90_45,  s_90_46,   s_91_0,   s_91_1,   s_91_2,   s_91_3;
wire   s_91_4,   s_91_5,   s_91_6,   s_91_7,   s_91_8,   s_91_9;
wire  s_91_10,  s_91_11,  s_91_12,  s_91_13,  s_91_14,  s_91_15;
wire  s_91_16,  s_91_17,  s_91_18,  s_91_19,  s_91_20,  s_91_21;
wire  s_91_22,  s_91_23,  s_91_24,  s_91_25,  s_91_26,  s_91_27;
wire  s_91_28,  s_91_29,  s_91_30,  s_91_31,  s_91_32,  s_91_33;
wire  s_91_34,  s_91_35,  s_91_36,  s_91_37,  s_91_38,  s_91_39;
wire  s_91_40,  s_91_41,  s_91_42,  s_91_43,  s_91_44,  s_91_45;
wire   s_92_0,   s_92_1,   s_92_2,   s_92_3,   s_92_4,   s_92_5;
wire   s_92_6,   s_92_7,   s_92_8,   s_92_9,  s_92_10,  s_92_11;
wire  s_92_12,  s_92_13,  s_92_14,  s_92_15,  s_92_16,  s_92_17;
wire  s_92_18,  s_92_19,  s_92_20,  s_92_21,  s_92_22,  s_92_23;
wire  s_92_24,  s_92_25,  s_92_26,  s_92_27,  s_92_28,  s_92_29;
wire  s_92_30,  s_92_31,  s_92_32,  s_92_33,  s_92_34,  s_92_35;
wire  s_92_36,  s_92_37,  s_92_38,  s_92_39,  s_92_40,  s_92_41;
wire  s_92_42,  s_92_43,  s_92_44,  s_92_45,  s_92_46,  s_92_47;
wire   s_93_0,   s_93_1,   s_93_2,   s_93_3,   s_93_4,   s_93_5;
wire   s_93_6,   s_93_7,   s_93_8,   s_93_9,  s_93_10,  s_93_11;
wire  s_93_12,  s_93_13,  s_93_14,  s_93_15,  s_93_16,  s_93_17;
wire  s_93_18,  s_93_19,  s_93_20,  s_93_21,  s_93_22,  s_93_23;
wire  s_93_24,  s_93_25,  s_93_26,  s_93_27,  s_93_28,  s_93_29;
wire  s_93_30,  s_93_31,  s_93_32,  s_93_33,  s_93_34,  s_93_35;
wire  s_93_36,  s_93_37,  s_93_38,  s_93_39,  s_93_40,  s_93_41;
wire  s_93_42,  s_93_43,  s_93_44,  s_93_45,  s_93_46,   s_94_0;
wire   s_94_1,   s_94_2,   s_94_3,   s_94_4,   s_94_5,   s_94_6;
wire   s_94_7,   s_94_8,   s_94_9,  s_94_10,  s_94_11,  s_94_12;
wire  s_94_13,  s_94_14,  s_94_15,  s_94_16,  s_94_17,  s_94_18;
wire  s_94_19,  s_94_20,  s_94_21,  s_94_22,  s_94_23,  s_94_24;
wire  s_94_25,  s_94_26,  s_94_27,  s_94_28,  s_94_29,  s_94_30;
wire  s_94_31,  s_94_32,  s_94_33,  s_94_34,  s_94_35,  s_94_36;
wire  s_94_37,  s_94_38,  s_94_39,  s_94_40,  s_94_41,  s_94_42;
wire  s_94_43,  s_94_44,  s_94_45,  s_94_46,  s_94_47,  s_94_48;
wire   s_95_0,   s_95_1,   s_95_2,   s_95_3,   s_95_4,   s_95_5;
wire   s_95_6,   s_95_7,   s_95_8,   s_95_9,  s_95_10,  s_95_11;
wire  s_95_12,  s_95_13,  s_95_14,  s_95_15,  s_95_16,  s_95_17;
wire  s_95_18,  s_95_19,  s_95_20,  s_95_21,  s_95_22,  s_95_23;
wire  s_95_24,  s_95_25,  s_95_26,  s_95_27,  s_95_28,  s_95_29;
wire  s_95_30,  s_95_31,  s_95_32,  s_95_33,  s_95_34,  s_95_35;
wire  s_95_36,  s_95_37,  s_95_38,  s_95_39,  s_95_40,  s_95_41;
wire  s_95_42,  s_95_43,  s_95_44,  s_95_45,  s_95_46,  s_95_47;
wire   s_96_0,   s_96_1,   s_96_2,   s_96_3,   s_96_4,   s_96_5;
wire   s_96_6,   s_96_7,   s_96_8,   s_96_9,  s_96_10,  s_96_11;
wire  s_96_12,  s_96_13,  s_96_14,  s_96_15,  s_96_16,  s_96_17;
wire  s_96_18,  s_96_19,  s_96_20,  s_96_21,  s_96_22,  s_96_23;
wire  s_96_24,  s_96_25,  s_96_26,  s_96_27,  s_96_28,  s_96_29;
wire  s_96_30,  s_96_31,  s_96_32,  s_96_33,  s_96_34,  s_96_35;
wire  s_96_36,  s_96_37,  s_96_38,  s_96_39,  s_96_40,  s_96_41;
wire  s_96_42,  s_96_43,  s_96_44,  s_96_45,  s_96_46,  s_96_47;
wire  s_96_48,  s_96_49,   s_97_0,   s_97_1,   s_97_2,   s_97_3;
wire   s_97_4,   s_97_5,   s_97_6,   s_97_7,   s_97_8,   s_97_9;
wire  s_97_10,  s_97_11,  s_97_12,  s_97_13,  s_97_14,  s_97_15;
wire  s_97_16,  s_97_17,  s_97_18,  s_97_19,  s_97_20,  s_97_21;
wire  s_97_22,  s_97_23,  s_97_24,  s_97_25,  s_97_26,  s_97_27;
wire  s_97_28,  s_97_29,  s_97_30,  s_97_31,  s_97_32,  s_97_33;
wire  s_97_34,  s_97_35,  s_97_36,  s_97_37,  s_97_38,  s_97_39;
wire  s_97_40,  s_97_41,  s_97_42,  s_97_43,  s_97_44,  s_97_45;
wire  s_97_46,  s_97_47,  s_97_48,   s_98_0,   s_98_1,   s_98_2;
wire   s_98_3,   s_98_4,   s_98_5,   s_98_6,   s_98_7,   s_98_8;
wire   s_98_9,  s_98_10,  s_98_11,  s_98_12,  s_98_13,  s_98_14;
wire  s_98_15,  s_98_16,  s_98_17,  s_98_18,  s_98_19,  s_98_20;
wire  s_98_21,  s_98_22,  s_98_23,  s_98_24,  s_98_25,  s_98_26;
wire  s_98_27,  s_98_28,  s_98_29,  s_98_30,  s_98_31,  s_98_32;
wire  s_98_33,  s_98_34,  s_98_35,  s_98_36,  s_98_37,  s_98_38;
wire  s_98_39,  s_98_40,  s_98_41,  s_98_42,  s_98_43,  s_98_44;
wire  s_98_45,  s_98_46,  s_98_47,  s_98_48,  s_98_49,  s_98_50;
wire   s_99_0,   s_99_1,   s_99_2,   s_99_3,   s_99_4,   s_99_5;
wire   s_99_6,   s_99_7,   s_99_8,   s_99_9,  s_99_10,  s_99_11;
wire  s_99_12,  s_99_13,  s_99_14,  s_99_15,  s_99_16,  s_99_17;
wire  s_99_18,  s_99_19,  s_99_20,  s_99_21,  s_99_22,  s_99_23;
wire  s_99_24,  s_99_25,  s_99_26,  s_99_27,  s_99_28,  s_99_29;
wire  s_99_30,  s_99_31,  s_99_32,  s_99_33,  s_99_34,  s_99_35;
wire  s_99_36,  s_99_37,  s_99_38,  s_99_39,  s_99_40,  s_99_41;
wire  s_99_42,  s_99_43,  s_99_44,  s_99_45,  s_99_46,  s_99_47;
wire  s_99_48,  s_99_49,  s_100_0,  s_100_1,  s_100_2,  s_100_3;
wire  s_100_4,  s_100_5,  s_100_6,  s_100_7,  s_100_8,  s_100_9;
wire s_100_10, s_100_11, s_100_12, s_100_13, s_100_14, s_100_15;
wire s_100_16, s_100_17, s_100_18, s_100_19, s_100_20, s_100_21;
wire s_100_22, s_100_23, s_100_24, s_100_25, s_100_26, s_100_27;
wire s_100_28, s_100_29, s_100_30, s_100_31, s_100_32, s_100_33;
wire s_100_34, s_100_35, s_100_36, s_100_37, s_100_38, s_100_39;
wire s_100_40, s_100_41, s_100_42, s_100_43, s_100_44, s_100_45;
wire s_100_46, s_100_47, s_100_48, s_100_49, s_100_50, s_100_51;
wire  s_101_0,  s_101_1,  s_101_2,  s_101_3,  s_101_4,  s_101_5;
wire  s_101_6,  s_101_7,  s_101_8,  s_101_9, s_101_10, s_101_11;
wire s_101_12, s_101_13, s_101_14, s_101_15, s_101_16, s_101_17;
wire s_101_18, s_101_19, s_101_20, s_101_21, s_101_22, s_101_23;
wire s_101_24, s_101_25, s_101_26, s_101_27, s_101_28, s_101_29;
wire s_101_30, s_101_31, s_101_32, s_101_33, s_101_34, s_101_35;
wire s_101_36, s_101_37, s_101_38, s_101_39, s_101_40, s_101_41;
wire s_101_42, s_101_43, s_101_44, s_101_45, s_101_46, s_101_47;
wire s_101_48, s_101_49, s_101_50,  s_102_0,  s_102_1,  s_102_2;
wire  s_102_3,  s_102_4,  s_102_5,  s_102_6,  s_102_7,  s_102_8;
wire  s_102_9, s_102_10, s_102_11, s_102_12, s_102_13, s_102_14;
wire s_102_15, s_102_16, s_102_17, s_102_18, s_102_19, s_102_20;
wire s_102_21, s_102_22, s_102_23, s_102_24, s_102_25, s_102_26;
wire s_102_27, s_102_28, s_102_29, s_102_30, s_102_31, s_102_32;
wire s_102_33, s_102_34, s_102_35, s_102_36, s_102_37, s_102_38;
wire s_102_39, s_102_40, s_102_41, s_102_42, s_102_43, s_102_44;
wire s_102_45, s_102_46, s_102_47, s_102_48, s_102_49, s_102_50;
wire s_102_51, s_102_52,  s_103_0,  s_103_1,  s_103_2,  s_103_3;
wire  s_103_4,  s_103_5,  s_103_6,  s_103_7,  s_103_8,  s_103_9;
wire s_103_10, s_103_11, s_103_12, s_103_13, s_103_14, s_103_15;
wire s_103_16, s_103_17, s_103_18, s_103_19, s_103_20, s_103_21;
wire s_103_22, s_103_23, s_103_24, s_103_25, s_103_26, s_103_27;
wire s_103_28, s_103_29, s_103_30, s_103_31, s_103_32, s_103_33;
wire s_103_34, s_103_35, s_103_36, s_103_37, s_103_38, s_103_39;
wire s_103_40, s_103_41, s_103_42, s_103_43, s_103_44, s_103_45;
wire s_103_46, s_103_47, s_103_48, s_103_49, s_103_50, s_103_51;
wire  s_104_0,  s_104_1,  s_104_2,  s_104_3,  s_104_4,  s_104_5;
wire  s_104_6,  s_104_7,  s_104_8,  s_104_9, s_104_10, s_104_11;
wire s_104_12, s_104_13, s_104_14, s_104_15, s_104_16, s_104_17;
wire s_104_18, s_104_19, s_104_20, s_104_21, s_104_22, s_104_23;
wire s_104_24, s_104_25, s_104_26, s_104_27, s_104_28, s_104_29;
wire s_104_30, s_104_31, s_104_32, s_104_33, s_104_34, s_104_35;
wire s_104_36, s_104_37, s_104_38, s_104_39, s_104_40, s_104_41;
wire s_104_42, s_104_43, s_104_44, s_104_45, s_104_46, s_104_47;
wire s_104_48, s_104_49, s_104_50, s_104_51, s_104_52, s_104_53;
wire  s_105_0,  s_105_1,  s_105_2,  s_105_3,  s_105_4,  s_105_5;
wire  s_105_6,  s_105_7,  s_105_8,  s_105_9, s_105_10, s_105_11;
wire s_105_12, s_105_13, s_105_14, s_105_15, s_105_16, s_105_17;
wire s_105_18, s_105_19, s_105_20, s_105_21, s_105_22, s_105_23;
wire s_105_24, s_105_25, s_105_26, s_105_27, s_105_28, s_105_29;
wire s_105_30, s_105_31, s_105_32, s_105_33, s_105_34, s_105_35;
wire s_105_36, s_105_37, s_105_38, s_105_39, s_105_40, s_105_41;
wire s_105_42, s_105_43, s_105_44, s_105_45, s_105_46, s_105_47;
wire s_105_48, s_105_49, s_105_50, s_105_51, s_105_52,  s_106_0;
wire  s_106_1,  s_106_2,  s_106_3,  s_106_4,  s_106_5,  s_106_6;
wire  s_106_7,  s_106_8,  s_106_9, s_106_10, s_106_11, s_106_12;
wire s_106_13, s_106_14, s_106_15, s_106_16, s_106_17, s_106_18;
wire s_106_19, s_106_20, s_106_21, s_106_22, s_106_23, s_106_24;
wire s_106_25, s_106_26, s_106_27, s_106_28, s_106_29, s_106_30;
wire s_106_31, s_106_32, s_106_33, s_106_34, s_106_35, s_106_36;
wire s_106_37, s_106_38, s_106_39, s_106_40, s_106_41, s_106_42;
wire s_106_43, s_106_44, s_106_45, s_106_46, s_106_47, s_106_48;
wire s_106_49, s_106_50, s_106_51, s_106_52, s_106_53, s_106_54;
wire  s_107_0,  s_107_1,  s_107_2,  s_107_3,  s_107_4,  s_107_5;
wire  s_107_6,  s_107_7,  s_107_8,  s_107_9, s_107_10, s_107_11;
wire s_107_12, s_107_13, s_107_14, s_107_15, s_107_16, s_107_17;
wire s_107_18, s_107_19, s_107_20, s_107_21, s_107_22, s_107_23;
wire s_107_24, s_107_25, s_107_26, s_107_27, s_107_28, s_107_29;
wire s_107_30, s_107_31, s_107_32, s_107_33, s_107_34, s_107_35;
wire s_107_36, s_107_37, s_107_38, s_107_39, s_107_40, s_107_41;
wire s_107_42, s_107_43, s_107_44, s_107_45, s_107_46, s_107_47;
wire s_107_48, s_107_49, s_107_50, s_107_51, s_107_52, s_107_53;
wire  s_108_0,  s_108_1,  s_108_2,  s_108_3,  s_108_4,  s_108_5;
wire  s_108_6,  s_108_7,  s_108_8,  s_108_9, s_108_10, s_108_11;
wire s_108_12, s_108_13, s_108_14, s_108_15, s_108_16, s_108_17;
wire s_108_18, s_108_19, s_108_20, s_108_21, s_108_22, s_108_23;
wire s_108_24, s_108_25, s_108_26, s_108_27, s_108_28, s_108_29;
wire s_108_30, s_108_31, s_108_32, s_108_33, s_108_34, s_108_35;
wire s_108_36, s_108_37, s_108_38, s_108_39, s_108_40, s_108_41;
wire s_108_42, s_108_43, s_108_44, s_108_45, s_108_46, s_108_47;
wire s_108_48, s_108_49, s_108_50, s_108_51, s_108_52, s_108_53;
wire s_108_54, s_108_55,  s_109_0,  s_109_1,  s_109_2,  s_109_3;
wire  s_109_4,  s_109_5,  s_109_6,  s_109_7,  s_109_8,  s_109_9;
wire s_109_10, s_109_11, s_109_12, s_109_13, s_109_14, s_109_15;
wire s_109_16, s_109_17, s_109_18, s_109_19, s_109_20, s_109_21;
wire s_109_22, s_109_23, s_109_24, s_109_25, s_109_26, s_109_27;
wire s_109_28, s_109_29, s_109_30, s_109_31, s_109_32, s_109_33;
wire s_109_34, s_109_35, s_109_36, s_109_37, s_109_38, s_109_39;
wire s_109_40, s_109_41, s_109_42, s_109_43, s_109_44, s_109_45;
wire s_109_46, s_109_47, s_109_48, s_109_49, s_109_50, s_109_51;
wire s_109_52, s_109_53, s_109_54,  s_110_0,  s_110_1,  s_110_2;
wire  s_110_3,  s_110_4,  s_110_5,  s_110_6,  s_110_7,  s_110_8;
wire  s_110_9, s_110_10, s_110_11, s_110_12, s_110_13, s_110_14;
wire s_110_15, s_110_16, s_110_17, s_110_18, s_110_19, s_110_20;
wire s_110_21, s_110_22, s_110_23, s_110_24, s_110_25, s_110_26;
wire s_110_27, s_110_28, s_110_29, s_110_30, s_110_31, s_110_32;
wire s_110_33, s_110_34, s_110_35, s_110_36, s_110_37, s_110_38;
wire s_110_39, s_110_40, s_110_41, s_110_42, s_110_43, s_110_44;
wire s_110_45, s_110_46, s_110_47, s_110_48, s_110_49, s_110_50;
wire s_110_51, s_110_52, s_110_53, s_110_54, s_110_55, s_110_56;
wire  s_111_0,  s_111_1,  s_111_2,  s_111_3,  s_111_4,  s_111_5;
wire  s_111_6,  s_111_7,  s_111_8,  s_111_9, s_111_10, s_111_11;
wire s_111_12, s_111_13, s_111_14, s_111_15, s_111_16, s_111_17;
wire s_111_18, s_111_19, s_111_20, s_111_21, s_111_22, s_111_23;
wire s_111_24, s_111_25, s_111_26, s_111_27, s_111_28, s_111_29;
wire s_111_30, s_111_31, s_111_32, s_111_33, s_111_34, s_111_35;
wire s_111_36, s_111_37, s_111_38, s_111_39, s_111_40, s_111_41;
wire s_111_42, s_111_43, s_111_44, s_111_45, s_111_46, s_111_47;
wire s_111_48, s_111_49, s_111_50, s_111_51, s_111_52, s_111_53;
wire s_111_54, s_111_55,  s_112_0,  s_112_1,  s_112_2,  s_112_3;
wire  s_112_4,  s_112_5,  s_112_6,  s_112_7,  s_112_8,  s_112_9;
wire s_112_10, s_112_11, s_112_12, s_112_13, s_112_14, s_112_15;
wire s_112_16, s_112_17, s_112_18, s_112_19, s_112_20, s_112_21;
wire s_112_22, s_112_23, s_112_24, s_112_25, s_112_26, s_112_27;
wire s_112_28, s_112_29, s_112_30, s_112_31, s_112_32, s_112_33;
wire s_112_34, s_112_35, s_112_36, s_112_37, s_112_38, s_112_39;
wire s_112_40, s_112_41, s_112_42, s_112_43, s_112_44, s_112_45;
wire s_112_46, s_112_47, s_112_48, s_112_49, s_112_50, s_112_51;
wire s_112_52, s_112_53, s_112_54, s_112_55, s_112_56, s_112_57;
wire  s_113_0,  s_113_1,  s_113_2,  s_113_3,  s_113_4,  s_113_5;
wire  s_113_6,  s_113_7,  s_113_8,  s_113_9, s_113_10, s_113_11;
wire s_113_12, s_113_13, s_113_14, s_113_15, s_113_16, s_113_17;
wire s_113_18, s_113_19, s_113_20, s_113_21, s_113_22, s_113_23;
wire s_113_24, s_113_25, s_113_26, s_113_27, s_113_28, s_113_29;
wire s_113_30, s_113_31, s_113_32, s_113_33, s_113_34, s_113_35;
wire s_113_36, s_113_37, s_113_38, s_113_39, s_113_40, s_113_41;
wire s_113_42, s_113_43, s_113_44, s_113_45, s_113_46, s_113_47;
wire s_113_48, s_113_49, s_113_50, s_113_51, s_113_52, s_113_53;
wire s_113_54, s_113_55, s_113_56,  s_114_0,  s_114_1,  s_114_2;
wire  s_114_3,  s_114_4,  s_114_5,  s_114_6,  s_114_7,  s_114_8;
wire  s_114_9, s_114_10, s_114_11, s_114_12, s_114_13, s_114_14;
wire s_114_15, s_114_16, s_114_17, s_114_18, s_114_19, s_114_20;
wire s_114_21, s_114_22, s_114_23, s_114_24, s_114_25, s_114_26;
wire s_114_27, s_114_28, s_114_29, s_114_30, s_114_31, s_114_32;
wire s_114_33, s_114_34, s_114_35, s_114_36, s_114_37, s_114_38;
wire s_114_39, s_114_40, s_114_41, s_114_42, s_114_43, s_114_44;
wire s_114_45, s_114_46, s_114_47, s_114_48, s_114_49, s_114_50;
wire s_114_51, s_114_52, s_114_53, s_114_54, s_114_55, s_114_56;
wire s_114_57, s_114_58,  s_115_0,  s_115_1,  s_115_2,  s_115_3;
wire  s_115_4,  s_115_5,  s_115_6,  s_115_7,  s_115_8,  s_115_9;
wire s_115_10, s_115_11, s_115_12, s_115_13, s_115_14, s_115_15;
wire s_115_16, s_115_17, s_115_18, s_115_19, s_115_20, s_115_21;
wire s_115_22, s_115_23, s_115_24, s_115_25, s_115_26, s_115_27;
wire s_115_28, s_115_29, s_115_30, s_115_31, s_115_32, s_115_33;
wire s_115_34, s_115_35, s_115_36, s_115_37, s_115_38, s_115_39;
wire s_115_40, s_115_41, s_115_42, s_115_43, s_115_44, s_115_45;
wire s_115_46, s_115_47, s_115_48, s_115_49, s_115_50, s_115_51;
wire s_115_52, s_115_53, s_115_54, s_115_55, s_115_56, s_115_57;
wire  s_116_0,  s_116_1,  s_116_2,  s_116_3,  s_116_4,  s_116_5;
wire  s_116_6,  s_116_7,  s_116_8,  s_116_9, s_116_10, s_116_11;
wire s_116_12, s_116_13, s_116_14, s_116_15, s_116_16, s_116_17;
wire s_116_18, s_116_19, s_116_20, s_116_21, s_116_22, s_116_23;
wire s_116_24, s_116_25, s_116_26, s_116_27, s_116_28, s_116_29;
wire s_116_30, s_116_31, s_116_32, s_116_33, s_116_34, s_116_35;
wire s_116_36, s_116_37, s_116_38, s_116_39, s_116_40, s_116_41;
wire s_116_42, s_116_43, s_116_44, s_116_45, s_116_46, s_116_47;
wire s_116_48, s_116_49, s_116_50, s_116_51, s_116_52, s_116_53;
wire s_116_54, s_116_55, s_116_56, s_116_57, s_116_58, s_116_59;
wire  s_117_0,  s_117_1,  s_117_2,  s_117_3,  s_117_4,  s_117_5;
wire  s_117_6,  s_117_7,  s_117_8,  s_117_9, s_117_10, s_117_11;
wire s_117_12, s_117_13, s_117_14, s_117_15, s_117_16, s_117_17;
wire s_117_18, s_117_19, s_117_20, s_117_21, s_117_22, s_117_23;
wire s_117_24, s_117_25, s_117_26, s_117_27, s_117_28, s_117_29;
wire s_117_30, s_117_31, s_117_32, s_117_33, s_117_34, s_117_35;
wire s_117_36, s_117_37, s_117_38, s_117_39, s_117_40, s_117_41;
wire s_117_42, s_117_43, s_117_44, s_117_45, s_117_46, s_117_47;
wire s_117_48, s_117_49, s_117_50, s_117_51, s_117_52, s_117_53;
wire s_117_54, s_117_55, s_117_56, s_117_57, s_117_58,  s_118_0;
wire  s_118_1,  s_118_2,  s_118_3,  s_118_4,  s_118_5,  s_118_6;
wire  s_118_7,  s_118_8,  s_118_9, s_118_10, s_118_11, s_118_12;
wire s_118_13, s_118_14, s_118_15, s_118_16, s_118_17, s_118_18;
wire s_118_19, s_118_20, s_118_21, s_118_22, s_118_23, s_118_24;
wire s_118_25, s_118_26, s_118_27, s_118_28, s_118_29, s_118_30;
wire s_118_31, s_118_32, s_118_33, s_118_34, s_118_35, s_118_36;
wire s_118_37, s_118_38, s_118_39, s_118_40, s_118_41, s_118_42;
wire s_118_43, s_118_44, s_118_45, s_118_46, s_118_47, s_118_48;
wire s_118_49, s_118_50, s_118_51, s_118_52, s_118_53, s_118_54;
wire s_118_55, s_118_56, s_118_57, s_118_58, s_118_59, s_118_60;
wire  s_119_0,  s_119_1,  s_119_2,  s_119_3,  s_119_4,  s_119_5;
wire  s_119_6,  s_119_7,  s_119_8,  s_119_9, s_119_10, s_119_11;
wire s_119_12, s_119_13, s_119_14, s_119_15, s_119_16, s_119_17;
wire s_119_18, s_119_19, s_119_20, s_119_21, s_119_22, s_119_23;
wire s_119_24, s_119_25, s_119_26, s_119_27, s_119_28, s_119_29;
wire s_119_30, s_119_31, s_119_32, s_119_33, s_119_34, s_119_35;
wire s_119_36, s_119_37, s_119_38, s_119_39, s_119_40, s_119_41;
wire s_119_42, s_119_43, s_119_44, s_119_45, s_119_46, s_119_47;
wire s_119_48, s_119_49, s_119_50, s_119_51, s_119_52, s_119_53;
wire s_119_54, s_119_55, s_119_56, s_119_57, s_119_58, s_119_59;
wire  s_120_0,  s_120_1,  s_120_2,  s_120_3,  s_120_4,  s_120_5;
wire  s_120_6,  s_120_7,  s_120_8,  s_120_9, s_120_10, s_120_11;
wire s_120_12, s_120_13, s_120_14, s_120_15, s_120_16, s_120_17;
wire s_120_18, s_120_19, s_120_20, s_120_21, s_120_22, s_120_23;
wire s_120_24, s_120_25, s_120_26, s_120_27, s_120_28, s_120_29;
wire s_120_30, s_120_31, s_120_32, s_120_33, s_120_34, s_120_35;
wire s_120_36, s_120_37, s_120_38, s_120_39, s_120_40, s_120_41;
wire s_120_42, s_120_43, s_120_44, s_120_45, s_120_46, s_120_47;
wire s_120_48, s_120_49, s_120_50, s_120_51, s_120_52, s_120_53;
wire s_120_54, s_120_55, s_120_56, s_120_57, s_120_58, s_120_59;
wire s_120_60, s_120_61,  s_121_0,  s_121_1,  s_121_2,  s_121_3;
wire  s_121_4,  s_121_5,  s_121_6,  s_121_7,  s_121_8,  s_121_9;
wire s_121_10, s_121_11, s_121_12, s_121_13, s_121_14, s_121_15;
wire s_121_16, s_121_17, s_121_18, s_121_19, s_121_20, s_121_21;
wire s_121_22, s_121_23, s_121_24, s_121_25, s_121_26, s_121_27;
wire s_121_28, s_121_29, s_121_30, s_121_31, s_121_32, s_121_33;
wire s_121_34, s_121_35, s_121_36, s_121_37, s_121_38, s_121_39;
wire s_121_40, s_121_41, s_121_42, s_121_43, s_121_44, s_121_45;
wire s_121_46, s_121_47, s_121_48, s_121_49, s_121_50, s_121_51;
wire s_121_52, s_121_53, s_121_54, s_121_55, s_121_56, s_121_57;
wire s_121_58, s_121_59, s_121_60,  s_122_0,  s_122_1,  s_122_2;
wire  s_122_3,  s_122_4,  s_122_5,  s_122_6,  s_122_7,  s_122_8;
wire  s_122_9, s_122_10, s_122_11, s_122_12, s_122_13, s_122_14;
wire s_122_15, s_122_16, s_122_17, s_122_18, s_122_19, s_122_20;
wire s_122_21, s_122_22, s_122_23, s_122_24, s_122_25, s_122_26;
wire s_122_27, s_122_28, s_122_29, s_122_30, s_122_31, s_122_32;
wire s_122_33, s_122_34, s_122_35, s_122_36, s_122_37, s_122_38;
wire s_122_39, s_122_40, s_122_41, s_122_42, s_122_43, s_122_44;
wire s_122_45, s_122_46, s_122_47, s_122_48, s_122_49, s_122_50;
wire s_122_51, s_122_52, s_122_53, s_122_54, s_122_55, s_122_56;
wire s_122_57, s_122_58, s_122_59, s_122_60, s_122_61, s_122_62;
wire  s_123_0,  s_123_1,  s_123_2,  s_123_3,  s_123_4,  s_123_5;
wire  s_123_6,  s_123_7,  s_123_8,  s_123_9, s_123_10, s_123_11;
wire s_123_12, s_123_13, s_123_14, s_123_15, s_123_16, s_123_17;
wire s_123_18, s_123_19, s_123_20, s_123_21, s_123_22, s_123_23;
wire s_123_24, s_123_25, s_123_26, s_123_27, s_123_28, s_123_29;
wire s_123_30, s_123_31, s_123_32, s_123_33, s_123_34, s_123_35;
wire s_123_36, s_123_37, s_123_38, s_123_39, s_123_40, s_123_41;
wire s_123_42, s_123_43, s_123_44, s_123_45, s_123_46, s_123_47;
wire s_123_48, s_123_49, s_123_50, s_123_51, s_123_52, s_123_53;
wire s_123_54, s_123_55, s_123_56, s_123_57, s_123_58, s_123_59;
wire s_123_60, s_123_61,  s_124_0,  s_124_1,  s_124_2,  s_124_3;
wire  s_124_4,  s_124_5,  s_124_6,  s_124_7,  s_124_8,  s_124_9;
wire s_124_10, s_124_11, s_124_12, s_124_13, s_124_14, s_124_15;
wire s_124_16, s_124_17, s_124_18, s_124_19, s_124_20, s_124_21;
wire s_124_22, s_124_23, s_124_24, s_124_25, s_124_26, s_124_27;
wire s_124_28, s_124_29, s_124_30, s_124_31, s_124_32, s_124_33;
wire s_124_34, s_124_35, s_124_36, s_124_37, s_124_38, s_124_39;
wire s_124_40, s_124_41, s_124_42, s_124_43, s_124_44, s_124_45;
wire s_124_46, s_124_47, s_124_48, s_124_49, s_124_50, s_124_51;
wire s_124_52, s_124_53, s_124_54, s_124_55, s_124_56, s_124_57;
wire s_124_58, s_124_59, s_124_60, s_124_61, s_124_62, s_124_63;
wire  s_125_0,  s_125_1,  s_125_2,  s_125_3,  s_125_4,  s_125_5;
wire  s_125_6,  s_125_7,  s_125_8,  s_125_9, s_125_10, s_125_11;
wire s_125_12, s_125_13, s_125_14, s_125_15, s_125_16, s_125_17;
wire s_125_18, s_125_19, s_125_20, s_125_21, s_125_22, s_125_23;
wire s_125_24, s_125_25, s_125_26, s_125_27, s_125_28, s_125_29;
wire s_125_30, s_125_31, s_125_32, s_125_33, s_125_34, s_125_35;
wire s_125_36, s_125_37, s_125_38, s_125_39, s_125_40, s_125_41;
wire s_125_42, s_125_43, s_125_44, s_125_45, s_125_46, s_125_47;
wire s_125_48, s_125_49, s_125_50, s_125_51, s_125_52, s_125_53;
wire s_125_54, s_125_55, s_125_56, s_125_57, s_125_58, s_125_59;
wire s_125_60, s_125_61, s_125_62,  s_126_0,  s_126_1,  s_126_2;
wire  s_126_3,  s_126_4,  s_126_5,  s_126_6,  s_126_7,  s_126_8;
wire  s_126_9, s_126_10, s_126_11, s_126_12, s_126_13, s_126_14;
wire s_126_15, s_126_16, s_126_17, s_126_18, s_126_19, s_126_20;
wire s_126_21, s_126_22, s_126_23, s_126_24, s_126_25, s_126_26;
wire s_126_27, s_126_28, s_126_29, s_126_30, s_126_31, s_126_32;
wire s_126_33, s_126_34, s_126_35, s_126_36, s_126_37, s_126_38;
wire s_126_39, s_126_40, s_126_41, s_126_42, s_126_43, s_126_44;
wire s_126_45, s_126_46, s_126_47, s_126_48, s_126_49, s_126_50;
wire s_126_51, s_126_52, s_126_53, s_126_54, s_126_55, s_126_56;
wire s_126_57, s_126_58, s_126_59, s_126_60, s_126_61, s_126_62;
wire s_126_63, s_126_64,  s_127_0,  s_127_1,  s_127_2,  s_127_3;
wire  s_127_4,  s_127_5,  s_127_6,  s_127_7,  s_127_8,  s_127_9;
wire s_127_10, s_127_11, s_127_12, s_127_13, s_127_14, s_127_15;
wire s_127_16, s_127_17, s_127_18, s_127_19, s_127_20, s_127_21;
wire s_127_22, s_127_23, s_127_24, s_127_25, s_127_26, s_127_27;
wire s_127_28, s_127_29, s_127_30, s_127_31, s_127_32, s_127_33;
wire s_127_34, s_127_35, s_127_36, s_127_37, s_127_38, s_127_39;
wire s_127_40, s_127_41, s_127_42, s_127_43, s_127_44, s_127_45;
wire s_127_46, s_127_47, s_127_48, s_127_49, s_127_50, s_127_51;
wire s_127_52, s_127_53, s_127_54, s_127_55, s_127_56, s_127_57;
wire s_127_58, s_127_59, s_127_60, s_127_61, s_127_62, s_127_63;
wire  s_128_0,  s_128_1,  s_128_2,  s_128_3,  s_128_4,  s_128_5;
wire  s_128_6,  s_128_7,  s_128_8,  s_128_9, s_128_10, s_128_11;
wire s_128_12, s_128_13, s_128_14, s_128_15, s_128_16, s_128_17;
wire s_128_18, s_128_19, s_128_20, s_128_21, s_128_22, s_128_23;
wire s_128_24, s_128_25, s_128_26, s_128_27, s_128_28, s_128_29;
wire s_128_30, s_128_31, s_128_32, s_128_33, s_128_34, s_128_35;
wire s_128_36, s_128_37, s_128_38, s_128_39, s_128_40, s_128_41;
wire s_128_42, s_128_43, s_128_44, s_128_45, s_128_46, s_128_47;
wire s_128_48, s_128_49, s_128_50, s_128_51, s_128_52, s_128_53;
wire s_128_54, s_128_55, s_128_56, s_128_57, s_128_58, s_128_59;
wire s_128_60, s_128_61, s_128_62, s_128_63, s_128_64,  s_129_0;
wire  s_129_1,  s_129_2,  s_129_3,  s_129_4,  s_129_5,  s_129_6;
wire  s_129_7,  s_129_8,  s_129_9, s_129_10, s_129_11, s_129_12;
wire s_129_13, s_129_14, s_129_15, s_129_16, s_129_17, s_129_18;
wire s_129_19, s_129_20, s_129_21, s_129_22, s_129_23, s_129_24;
wire s_129_25, s_129_26, s_129_27, s_129_28, s_129_29, s_129_30;
wire s_129_31, s_129_32, s_129_33, s_129_34, s_129_35, s_129_36;
wire s_129_37, s_129_38, s_129_39, s_129_40, s_129_41, s_129_42;
wire s_129_43, s_129_44, s_129_45, s_129_46, s_129_47, s_129_48;
wire s_129_49, s_129_50, s_129_51, s_129_52, s_129_53, s_129_54;
wire s_129_55, s_129_56, s_129_57, s_129_58, s_129_59, s_129_60;
wire s_129_61, s_129_62, s_129_63, s_129_64,  s_130_0,  s_130_1;
wire  s_130_2,  s_130_3,  s_130_4,  s_130_5,  s_130_6,  s_130_7;
wire  s_130_8,  s_130_9, s_130_10, s_130_11, s_130_12, s_130_13;
wire s_130_14, s_130_15, s_130_16, s_130_17, s_130_18, s_130_19;
wire s_130_20, s_130_21, s_130_22, s_130_23, s_130_24, s_130_25;
wire s_130_26, s_130_27, s_130_28, s_130_29, s_130_30, s_130_31;
wire s_130_32, s_130_33, s_130_34, s_130_35, s_130_36, s_130_37;
wire s_130_38, s_130_39, s_130_40, s_130_41, s_130_42, s_130_43;
wire s_130_44, s_130_45, s_130_46, s_130_47, s_130_48, s_130_49;
wire s_130_50, s_130_51, s_130_52, s_130_53, s_130_54, s_130_55;
wire s_130_56, s_130_57, s_130_58, s_130_59, s_130_60, s_130_61;
wire s_130_62, s_130_63,  s_131_0,  s_131_1,  s_131_2,  s_131_3;
wire  s_131_4,  s_131_5,  s_131_6,  s_131_7,  s_131_8,  s_131_9;
wire s_131_10, s_131_11, s_131_12, s_131_13, s_131_14, s_131_15;
wire s_131_16, s_131_17, s_131_18, s_131_19, s_131_20, s_131_21;
wire s_131_22, s_131_23, s_131_24, s_131_25, s_131_26, s_131_27;
wire s_131_28, s_131_29, s_131_30, s_131_31, s_131_32, s_131_33;
wire s_131_34, s_131_35, s_131_36, s_131_37, s_131_38, s_131_39;
wire s_131_40, s_131_41, s_131_42, s_131_43, s_131_44, s_131_45;
wire s_131_46, s_131_47, s_131_48, s_131_49, s_131_50, s_131_51;
wire s_131_52, s_131_53, s_131_54, s_131_55, s_131_56, s_131_57;
wire s_131_58, s_131_59, s_131_60, s_131_61, s_131_62, s_131_63;
wire  s_132_0,  s_132_1,  s_132_2,  s_132_3,  s_132_4,  s_132_5;
wire  s_132_6,  s_132_7,  s_132_8,  s_132_9, s_132_10, s_132_11;
wire s_132_12, s_132_13, s_132_14, s_132_15, s_132_16, s_132_17;
wire s_132_18, s_132_19, s_132_20, s_132_21, s_132_22, s_132_23;
wire s_132_24, s_132_25, s_132_26, s_132_27, s_132_28, s_132_29;
wire s_132_30, s_132_31, s_132_32, s_132_33, s_132_34, s_132_35;
wire s_132_36, s_132_37, s_132_38, s_132_39, s_132_40, s_132_41;
wire s_132_42, s_132_43, s_132_44, s_132_45, s_132_46, s_132_47;
wire s_132_48, s_132_49, s_132_50, s_132_51, s_132_52, s_132_53;
wire s_132_54, s_132_55, s_132_56, s_132_57, s_132_58, s_132_59;
wire s_132_60, s_132_61, s_132_62,  s_133_0,  s_133_1,  s_133_2;
wire  s_133_3,  s_133_4,  s_133_5,  s_133_6,  s_133_7,  s_133_8;
wire  s_133_9, s_133_10, s_133_11, s_133_12, s_133_13, s_133_14;
wire s_133_15, s_133_16, s_133_17, s_133_18, s_133_19, s_133_20;
wire s_133_21, s_133_22, s_133_23, s_133_24, s_133_25, s_133_26;
wire s_133_27, s_133_28, s_133_29, s_133_30, s_133_31, s_133_32;
wire s_133_33, s_133_34, s_133_35, s_133_36, s_133_37, s_133_38;
wire s_133_39, s_133_40, s_133_41, s_133_42, s_133_43, s_133_44;
wire s_133_45, s_133_46, s_133_47, s_133_48, s_133_49, s_133_50;
wire s_133_51, s_133_52, s_133_53, s_133_54, s_133_55, s_133_56;
wire s_133_57, s_133_58, s_133_59, s_133_60, s_133_61, s_133_62;
wire  s_134_0,  s_134_1,  s_134_2,  s_134_3,  s_134_4,  s_134_5;
wire  s_134_6,  s_134_7,  s_134_8,  s_134_9, s_134_10, s_134_11;
wire s_134_12, s_134_13, s_134_14, s_134_15, s_134_16, s_134_17;
wire s_134_18, s_134_19, s_134_20, s_134_21, s_134_22, s_134_23;
wire s_134_24, s_134_25, s_134_26, s_134_27, s_134_28, s_134_29;
wire s_134_30, s_134_31, s_134_32, s_134_33, s_134_34, s_134_35;
wire s_134_36, s_134_37, s_134_38, s_134_39, s_134_40, s_134_41;
wire s_134_42, s_134_43, s_134_44, s_134_45, s_134_46, s_134_47;
wire s_134_48, s_134_49, s_134_50, s_134_51, s_134_52, s_134_53;
wire s_134_54, s_134_55, s_134_56, s_134_57, s_134_58, s_134_59;
wire s_134_60, s_134_61,  s_135_0,  s_135_1,  s_135_2,  s_135_3;
wire  s_135_4,  s_135_5,  s_135_6,  s_135_7,  s_135_8,  s_135_9;
wire s_135_10, s_135_11, s_135_12, s_135_13, s_135_14, s_135_15;
wire s_135_16, s_135_17, s_135_18, s_135_19, s_135_20, s_135_21;
wire s_135_22, s_135_23, s_135_24, s_135_25, s_135_26, s_135_27;
wire s_135_28, s_135_29, s_135_30, s_135_31, s_135_32, s_135_33;
wire s_135_34, s_135_35, s_135_36, s_135_37, s_135_38, s_135_39;
wire s_135_40, s_135_41, s_135_42, s_135_43, s_135_44, s_135_45;
wire s_135_46, s_135_47, s_135_48, s_135_49, s_135_50, s_135_51;
wire s_135_52, s_135_53, s_135_54, s_135_55, s_135_56, s_135_57;
wire s_135_58, s_135_59, s_135_60, s_135_61,  s_136_0,  s_136_1;
wire  s_136_2,  s_136_3,  s_136_4,  s_136_5,  s_136_6,  s_136_7;
wire  s_136_8,  s_136_9, s_136_10, s_136_11, s_136_12, s_136_13;
wire s_136_14, s_136_15, s_136_16, s_136_17, s_136_18, s_136_19;
wire s_136_20, s_136_21, s_136_22, s_136_23, s_136_24, s_136_25;
wire s_136_26, s_136_27, s_136_28, s_136_29, s_136_30, s_136_31;
wire s_136_32, s_136_33, s_136_34, s_136_35, s_136_36, s_136_37;
wire s_136_38, s_136_39, s_136_40, s_136_41, s_136_42, s_136_43;
wire s_136_44, s_136_45, s_136_46, s_136_47, s_136_48, s_136_49;
wire s_136_50, s_136_51, s_136_52, s_136_53, s_136_54, s_136_55;
wire s_136_56, s_136_57, s_136_58, s_136_59, s_136_60,  s_137_0;
wire  s_137_1,  s_137_2,  s_137_3,  s_137_4,  s_137_5,  s_137_6;
wire  s_137_7,  s_137_8,  s_137_9, s_137_10, s_137_11, s_137_12;
wire s_137_13, s_137_14, s_137_15, s_137_16, s_137_17, s_137_18;
wire s_137_19, s_137_20, s_137_21, s_137_22, s_137_23, s_137_24;
wire s_137_25, s_137_26, s_137_27, s_137_28, s_137_29, s_137_30;
wire s_137_31, s_137_32, s_137_33, s_137_34, s_137_35, s_137_36;
wire s_137_37, s_137_38, s_137_39, s_137_40, s_137_41, s_137_42;
wire s_137_43, s_137_44, s_137_45, s_137_46, s_137_47, s_137_48;
wire s_137_49, s_137_50, s_137_51, s_137_52, s_137_53, s_137_54;
wire s_137_55, s_137_56, s_137_57, s_137_58, s_137_59, s_137_60;
wire  s_138_0,  s_138_1,  s_138_2,  s_138_3,  s_138_4,  s_138_5;
wire  s_138_6,  s_138_7,  s_138_8,  s_138_9, s_138_10, s_138_11;
wire s_138_12, s_138_13, s_138_14, s_138_15, s_138_16, s_138_17;
wire s_138_18, s_138_19, s_138_20, s_138_21, s_138_22, s_138_23;
wire s_138_24, s_138_25, s_138_26, s_138_27, s_138_28, s_138_29;
wire s_138_30, s_138_31, s_138_32, s_138_33, s_138_34, s_138_35;
wire s_138_36, s_138_37, s_138_38, s_138_39, s_138_40, s_138_41;
wire s_138_42, s_138_43, s_138_44, s_138_45, s_138_46, s_138_47;
wire s_138_48, s_138_49, s_138_50, s_138_51, s_138_52, s_138_53;
wire s_138_54, s_138_55, s_138_56, s_138_57, s_138_58, s_138_59;
wire  s_139_0,  s_139_1,  s_139_2,  s_139_3,  s_139_4,  s_139_5;
wire  s_139_6,  s_139_7,  s_139_8,  s_139_9, s_139_10, s_139_11;
wire s_139_12, s_139_13, s_139_14, s_139_15, s_139_16, s_139_17;
wire s_139_18, s_139_19, s_139_20, s_139_21, s_139_22, s_139_23;
wire s_139_24, s_139_25, s_139_26, s_139_27, s_139_28, s_139_29;
wire s_139_30, s_139_31, s_139_32, s_139_33, s_139_34, s_139_35;
wire s_139_36, s_139_37, s_139_38, s_139_39, s_139_40, s_139_41;
wire s_139_42, s_139_43, s_139_44, s_139_45, s_139_46, s_139_47;
wire s_139_48, s_139_49, s_139_50, s_139_51, s_139_52, s_139_53;
wire s_139_54, s_139_55, s_139_56, s_139_57, s_139_58, s_139_59;
wire  s_140_0,  s_140_1,  s_140_2,  s_140_3,  s_140_4,  s_140_5;
wire  s_140_6,  s_140_7,  s_140_8,  s_140_9, s_140_10, s_140_11;
wire s_140_12, s_140_13, s_140_14, s_140_15, s_140_16, s_140_17;
wire s_140_18, s_140_19, s_140_20, s_140_21, s_140_22, s_140_23;
wire s_140_24, s_140_25, s_140_26, s_140_27, s_140_28, s_140_29;
wire s_140_30, s_140_31, s_140_32, s_140_33, s_140_34, s_140_35;
wire s_140_36, s_140_37, s_140_38, s_140_39, s_140_40, s_140_41;
wire s_140_42, s_140_43, s_140_44, s_140_45, s_140_46, s_140_47;
wire s_140_48, s_140_49, s_140_50, s_140_51, s_140_52, s_140_53;
wire s_140_54, s_140_55, s_140_56, s_140_57, s_140_58,  s_141_0;
wire  s_141_1,  s_141_2,  s_141_3,  s_141_4,  s_141_5,  s_141_6;
wire  s_141_7,  s_141_8,  s_141_9, s_141_10, s_141_11, s_141_12;
wire s_141_13, s_141_14, s_141_15, s_141_16, s_141_17, s_141_18;
wire s_141_19, s_141_20, s_141_21, s_141_22, s_141_23, s_141_24;
wire s_141_25, s_141_26, s_141_27, s_141_28, s_141_29, s_141_30;
wire s_141_31, s_141_32, s_141_33, s_141_34, s_141_35, s_141_36;
wire s_141_37, s_141_38, s_141_39, s_141_40, s_141_41, s_141_42;
wire s_141_43, s_141_44, s_141_45, s_141_46, s_141_47, s_141_48;
wire s_141_49, s_141_50, s_141_51, s_141_52, s_141_53, s_141_54;
wire s_141_55, s_141_56, s_141_57, s_141_58,  s_142_0,  s_142_1;
wire  s_142_2,  s_142_3,  s_142_4,  s_142_5,  s_142_6,  s_142_7;
wire  s_142_8,  s_142_9, s_142_10, s_142_11, s_142_12, s_142_13;
wire s_142_14, s_142_15, s_142_16, s_142_17, s_142_18, s_142_19;
wire s_142_20, s_142_21, s_142_22, s_142_23, s_142_24, s_142_25;
wire s_142_26, s_142_27, s_142_28, s_142_29, s_142_30, s_142_31;
wire s_142_32, s_142_33, s_142_34, s_142_35, s_142_36, s_142_37;
wire s_142_38, s_142_39, s_142_40, s_142_41, s_142_42, s_142_43;
wire s_142_44, s_142_45, s_142_46, s_142_47, s_142_48, s_142_49;
wire s_142_50, s_142_51, s_142_52, s_142_53, s_142_54, s_142_55;
wire s_142_56, s_142_57,  s_143_0,  s_143_1,  s_143_2,  s_143_3;
wire  s_143_4,  s_143_5,  s_143_6,  s_143_7,  s_143_8,  s_143_9;
wire s_143_10, s_143_11, s_143_12, s_143_13, s_143_14, s_143_15;
wire s_143_16, s_143_17, s_143_18, s_143_19, s_143_20, s_143_21;
wire s_143_22, s_143_23, s_143_24, s_143_25, s_143_26, s_143_27;
wire s_143_28, s_143_29, s_143_30, s_143_31, s_143_32, s_143_33;
wire s_143_34, s_143_35, s_143_36, s_143_37, s_143_38, s_143_39;
wire s_143_40, s_143_41, s_143_42, s_143_43, s_143_44, s_143_45;
wire s_143_46, s_143_47, s_143_48, s_143_49, s_143_50, s_143_51;
wire s_143_52, s_143_53, s_143_54, s_143_55, s_143_56, s_143_57;
wire  s_144_0,  s_144_1,  s_144_2,  s_144_3,  s_144_4,  s_144_5;
wire  s_144_6,  s_144_7,  s_144_8,  s_144_9, s_144_10, s_144_11;
wire s_144_12, s_144_13, s_144_14, s_144_15, s_144_16, s_144_17;
wire s_144_18, s_144_19, s_144_20, s_144_21, s_144_22, s_144_23;
wire s_144_24, s_144_25, s_144_26, s_144_27, s_144_28, s_144_29;
wire s_144_30, s_144_31, s_144_32, s_144_33, s_144_34, s_144_35;
wire s_144_36, s_144_37, s_144_38, s_144_39, s_144_40, s_144_41;
wire s_144_42, s_144_43, s_144_44, s_144_45, s_144_46, s_144_47;
wire s_144_48, s_144_49, s_144_50, s_144_51, s_144_52, s_144_53;
wire s_144_54, s_144_55, s_144_56,  s_145_0,  s_145_1,  s_145_2;
wire  s_145_3,  s_145_4,  s_145_5,  s_145_6,  s_145_7,  s_145_8;
wire  s_145_9, s_145_10, s_145_11, s_145_12, s_145_13, s_145_14;
wire s_145_15, s_145_16, s_145_17, s_145_18, s_145_19, s_145_20;
wire s_145_21, s_145_22, s_145_23, s_145_24, s_145_25, s_145_26;
wire s_145_27, s_145_28, s_145_29, s_145_30, s_145_31, s_145_32;
wire s_145_33, s_145_34, s_145_35, s_145_36, s_145_37, s_145_38;
wire s_145_39, s_145_40, s_145_41, s_145_42, s_145_43, s_145_44;
wire s_145_45, s_145_46, s_145_47, s_145_48, s_145_49, s_145_50;
wire s_145_51, s_145_52, s_145_53, s_145_54, s_145_55, s_145_56;
wire  s_146_0,  s_146_1,  s_146_2,  s_146_3,  s_146_4,  s_146_5;
wire  s_146_6,  s_146_7,  s_146_8,  s_146_9, s_146_10, s_146_11;
wire s_146_12, s_146_13, s_146_14, s_146_15, s_146_16, s_146_17;
wire s_146_18, s_146_19, s_146_20, s_146_21, s_146_22, s_146_23;
wire s_146_24, s_146_25, s_146_26, s_146_27, s_146_28, s_146_29;
wire s_146_30, s_146_31, s_146_32, s_146_33, s_146_34, s_146_35;
wire s_146_36, s_146_37, s_146_38, s_146_39, s_146_40, s_146_41;
wire s_146_42, s_146_43, s_146_44, s_146_45, s_146_46, s_146_47;
wire s_146_48, s_146_49, s_146_50, s_146_51, s_146_52, s_146_53;
wire s_146_54, s_146_55,  s_147_0,  s_147_1,  s_147_2,  s_147_3;
wire  s_147_4,  s_147_5,  s_147_6,  s_147_7,  s_147_8,  s_147_9;
wire s_147_10, s_147_11, s_147_12, s_147_13, s_147_14, s_147_15;
wire s_147_16, s_147_17, s_147_18, s_147_19, s_147_20, s_147_21;
wire s_147_22, s_147_23, s_147_24, s_147_25, s_147_26, s_147_27;
wire s_147_28, s_147_29, s_147_30, s_147_31, s_147_32, s_147_33;
wire s_147_34, s_147_35, s_147_36, s_147_37, s_147_38, s_147_39;
wire s_147_40, s_147_41, s_147_42, s_147_43, s_147_44, s_147_45;
wire s_147_46, s_147_47, s_147_48, s_147_49, s_147_50, s_147_51;
wire s_147_52, s_147_53, s_147_54, s_147_55,  s_148_0,  s_148_1;
wire  s_148_2,  s_148_3,  s_148_4,  s_148_5,  s_148_6,  s_148_7;
wire  s_148_8,  s_148_9, s_148_10, s_148_11, s_148_12, s_148_13;
wire s_148_14, s_148_15, s_148_16, s_148_17, s_148_18, s_148_19;
wire s_148_20, s_148_21, s_148_22, s_148_23, s_148_24, s_148_25;
wire s_148_26, s_148_27, s_148_28, s_148_29, s_148_30, s_148_31;
wire s_148_32, s_148_33, s_148_34, s_148_35, s_148_36, s_148_37;
wire s_148_38, s_148_39, s_148_40, s_148_41, s_148_42, s_148_43;
wire s_148_44, s_148_45, s_148_46, s_148_47, s_148_48, s_148_49;
wire s_148_50, s_148_51, s_148_52, s_148_53, s_148_54,  s_149_0;
wire  s_149_1,  s_149_2,  s_149_3,  s_149_4,  s_149_5,  s_149_6;
wire  s_149_7,  s_149_8,  s_149_9, s_149_10, s_149_11, s_149_12;
wire s_149_13, s_149_14, s_149_15, s_149_16, s_149_17, s_149_18;
wire s_149_19, s_149_20, s_149_21, s_149_22, s_149_23, s_149_24;
wire s_149_25, s_149_26, s_149_27, s_149_28, s_149_29, s_149_30;
wire s_149_31, s_149_32, s_149_33, s_149_34, s_149_35, s_149_36;
wire s_149_37, s_149_38, s_149_39, s_149_40, s_149_41, s_149_42;
wire s_149_43, s_149_44, s_149_45, s_149_46, s_149_47, s_149_48;
wire s_149_49, s_149_50, s_149_51, s_149_52, s_149_53, s_149_54;
wire  s_150_0,  s_150_1,  s_150_2,  s_150_3,  s_150_4,  s_150_5;
wire  s_150_6,  s_150_7,  s_150_8,  s_150_9, s_150_10, s_150_11;
wire s_150_12, s_150_13, s_150_14, s_150_15, s_150_16, s_150_17;
wire s_150_18, s_150_19, s_150_20, s_150_21, s_150_22, s_150_23;
wire s_150_24, s_150_25, s_150_26, s_150_27, s_150_28, s_150_29;
wire s_150_30, s_150_31, s_150_32, s_150_33, s_150_34, s_150_35;
wire s_150_36, s_150_37, s_150_38, s_150_39, s_150_40, s_150_41;
wire s_150_42, s_150_43, s_150_44, s_150_45, s_150_46, s_150_47;
wire s_150_48, s_150_49, s_150_50, s_150_51, s_150_52, s_150_53;
wire  s_151_0,  s_151_1,  s_151_2,  s_151_3,  s_151_4,  s_151_5;
wire  s_151_6,  s_151_7,  s_151_8,  s_151_9, s_151_10, s_151_11;
wire s_151_12, s_151_13, s_151_14, s_151_15, s_151_16, s_151_17;
wire s_151_18, s_151_19, s_151_20, s_151_21, s_151_22, s_151_23;
wire s_151_24, s_151_25, s_151_26, s_151_27, s_151_28, s_151_29;
wire s_151_30, s_151_31, s_151_32, s_151_33, s_151_34, s_151_35;
wire s_151_36, s_151_37, s_151_38, s_151_39, s_151_40, s_151_41;
wire s_151_42, s_151_43, s_151_44, s_151_45, s_151_46, s_151_47;
wire s_151_48, s_151_49, s_151_50, s_151_51, s_151_52, s_151_53;
wire  s_152_0,  s_152_1,  s_152_2,  s_152_3,  s_152_4,  s_152_5;
wire  s_152_6,  s_152_7,  s_152_8,  s_152_9, s_152_10, s_152_11;
wire s_152_12, s_152_13, s_152_14, s_152_15, s_152_16, s_152_17;
wire s_152_18, s_152_19, s_152_20, s_152_21, s_152_22, s_152_23;
wire s_152_24, s_152_25, s_152_26, s_152_27, s_152_28, s_152_29;
wire s_152_30, s_152_31, s_152_32, s_152_33, s_152_34, s_152_35;
wire s_152_36, s_152_37, s_152_38, s_152_39, s_152_40, s_152_41;
wire s_152_42, s_152_43, s_152_44, s_152_45, s_152_46, s_152_47;
wire s_152_48, s_152_49, s_152_50, s_152_51, s_152_52,  s_153_0;
wire  s_153_1,  s_153_2,  s_153_3,  s_153_4,  s_153_5,  s_153_6;
wire  s_153_7,  s_153_8,  s_153_9, s_153_10, s_153_11, s_153_12;
wire s_153_13, s_153_14, s_153_15, s_153_16, s_153_17, s_153_18;
wire s_153_19, s_153_20, s_153_21, s_153_22, s_153_23, s_153_24;
wire s_153_25, s_153_26, s_153_27, s_153_28, s_153_29, s_153_30;
wire s_153_31, s_153_32, s_153_33, s_153_34, s_153_35, s_153_36;
wire s_153_37, s_153_38, s_153_39, s_153_40, s_153_41, s_153_42;
wire s_153_43, s_153_44, s_153_45, s_153_46, s_153_47, s_153_48;
wire s_153_49, s_153_50, s_153_51, s_153_52,  s_154_0,  s_154_1;
wire  s_154_2,  s_154_3,  s_154_4,  s_154_5,  s_154_6,  s_154_7;
wire  s_154_8,  s_154_9, s_154_10, s_154_11, s_154_12, s_154_13;
wire s_154_14, s_154_15, s_154_16, s_154_17, s_154_18, s_154_19;
wire s_154_20, s_154_21, s_154_22, s_154_23, s_154_24, s_154_25;
wire s_154_26, s_154_27, s_154_28, s_154_29, s_154_30, s_154_31;
wire s_154_32, s_154_33, s_154_34, s_154_35, s_154_36, s_154_37;
wire s_154_38, s_154_39, s_154_40, s_154_41, s_154_42, s_154_43;
wire s_154_44, s_154_45, s_154_46, s_154_47, s_154_48, s_154_49;
wire s_154_50, s_154_51,  s_155_0,  s_155_1,  s_155_2,  s_155_3;
wire  s_155_4,  s_155_5,  s_155_6,  s_155_7,  s_155_8,  s_155_9;
wire s_155_10, s_155_11, s_155_12, s_155_13, s_155_14, s_155_15;
wire s_155_16, s_155_17, s_155_18, s_155_19, s_155_20, s_155_21;
wire s_155_22, s_155_23, s_155_24, s_155_25, s_155_26, s_155_27;
wire s_155_28, s_155_29, s_155_30, s_155_31, s_155_32, s_155_33;
wire s_155_34, s_155_35, s_155_36, s_155_37, s_155_38, s_155_39;
wire s_155_40, s_155_41, s_155_42, s_155_43, s_155_44, s_155_45;
wire s_155_46, s_155_47, s_155_48, s_155_49, s_155_50, s_155_51;
wire  s_156_0,  s_156_1,  s_156_2,  s_156_3,  s_156_4,  s_156_5;
wire  s_156_6,  s_156_7,  s_156_8,  s_156_9, s_156_10, s_156_11;
wire s_156_12, s_156_13, s_156_14, s_156_15, s_156_16, s_156_17;
wire s_156_18, s_156_19, s_156_20, s_156_21, s_156_22, s_156_23;
wire s_156_24, s_156_25, s_156_26, s_156_27, s_156_28, s_156_29;
wire s_156_30, s_156_31, s_156_32, s_156_33, s_156_34, s_156_35;
wire s_156_36, s_156_37, s_156_38, s_156_39, s_156_40, s_156_41;
wire s_156_42, s_156_43, s_156_44, s_156_45, s_156_46, s_156_47;
wire s_156_48, s_156_49, s_156_50,  s_157_0,  s_157_1,  s_157_2;
wire  s_157_3,  s_157_4,  s_157_5,  s_157_6,  s_157_7,  s_157_8;
wire  s_157_9, s_157_10, s_157_11, s_157_12, s_157_13, s_157_14;
wire s_157_15, s_157_16, s_157_17, s_157_18, s_157_19, s_157_20;
wire s_157_21, s_157_22, s_157_23, s_157_24, s_157_25, s_157_26;
wire s_157_27, s_157_28, s_157_29, s_157_30, s_157_31, s_157_32;
wire s_157_33, s_157_34, s_157_35, s_157_36, s_157_37, s_157_38;
wire s_157_39, s_157_40, s_157_41, s_157_42, s_157_43, s_157_44;
wire s_157_45, s_157_46, s_157_47, s_157_48, s_157_49, s_157_50;
wire  s_158_0,  s_158_1,  s_158_2,  s_158_3,  s_158_4,  s_158_5;
wire  s_158_6,  s_158_7,  s_158_8,  s_158_9, s_158_10, s_158_11;
wire s_158_12, s_158_13, s_158_14, s_158_15, s_158_16, s_158_17;
wire s_158_18, s_158_19, s_158_20, s_158_21, s_158_22, s_158_23;
wire s_158_24, s_158_25, s_158_26, s_158_27, s_158_28, s_158_29;
wire s_158_30, s_158_31, s_158_32, s_158_33, s_158_34, s_158_35;
wire s_158_36, s_158_37, s_158_38, s_158_39, s_158_40, s_158_41;
wire s_158_42, s_158_43, s_158_44, s_158_45, s_158_46, s_158_47;
wire s_158_48, s_158_49,  s_159_0,  s_159_1,  s_159_2,  s_159_3;
wire  s_159_4,  s_159_5,  s_159_6,  s_159_7,  s_159_8,  s_159_9;
wire s_159_10, s_159_11, s_159_12, s_159_13, s_159_14, s_159_15;
wire s_159_16, s_159_17, s_159_18, s_159_19, s_159_20, s_159_21;
wire s_159_22, s_159_23, s_159_24, s_159_25, s_159_26, s_159_27;
wire s_159_28, s_159_29, s_159_30, s_159_31, s_159_32, s_159_33;
wire s_159_34, s_159_35, s_159_36, s_159_37, s_159_38, s_159_39;
wire s_159_40, s_159_41, s_159_42, s_159_43, s_159_44, s_159_45;
wire s_159_46, s_159_47, s_159_48, s_159_49,  s_160_0,  s_160_1;
wire  s_160_2,  s_160_3,  s_160_4,  s_160_5,  s_160_6,  s_160_7;
wire  s_160_8,  s_160_9, s_160_10, s_160_11, s_160_12, s_160_13;
wire s_160_14, s_160_15, s_160_16, s_160_17, s_160_18, s_160_19;
wire s_160_20, s_160_21, s_160_22, s_160_23, s_160_24, s_160_25;
wire s_160_26, s_160_27, s_160_28, s_160_29, s_160_30, s_160_31;
wire s_160_32, s_160_33, s_160_34, s_160_35, s_160_36, s_160_37;
wire s_160_38, s_160_39, s_160_40, s_160_41, s_160_42, s_160_43;
wire s_160_44, s_160_45, s_160_46, s_160_47, s_160_48,  s_161_0;
wire  s_161_1,  s_161_2,  s_161_3,  s_161_4,  s_161_5,  s_161_6;
wire  s_161_7,  s_161_8,  s_161_9, s_161_10, s_161_11, s_161_12;
wire s_161_13, s_161_14, s_161_15, s_161_16, s_161_17, s_161_18;
wire s_161_19, s_161_20, s_161_21, s_161_22, s_161_23, s_161_24;
wire s_161_25, s_161_26, s_161_27, s_161_28, s_161_29, s_161_30;
wire s_161_31, s_161_32, s_161_33, s_161_34, s_161_35, s_161_36;
wire s_161_37, s_161_38, s_161_39, s_161_40, s_161_41, s_161_42;
wire s_161_43, s_161_44, s_161_45, s_161_46, s_161_47, s_161_48;
wire  s_162_0,  s_162_1,  s_162_2,  s_162_3,  s_162_4,  s_162_5;
wire  s_162_6,  s_162_7,  s_162_8,  s_162_9, s_162_10, s_162_11;
wire s_162_12, s_162_13, s_162_14, s_162_15, s_162_16, s_162_17;
wire s_162_18, s_162_19, s_162_20, s_162_21, s_162_22, s_162_23;
wire s_162_24, s_162_25, s_162_26, s_162_27, s_162_28, s_162_29;
wire s_162_30, s_162_31, s_162_32, s_162_33, s_162_34, s_162_35;
wire s_162_36, s_162_37, s_162_38, s_162_39, s_162_40, s_162_41;
wire s_162_42, s_162_43, s_162_44, s_162_45, s_162_46, s_162_47;
wire  s_163_0,  s_163_1,  s_163_2,  s_163_3,  s_163_4,  s_163_5;
wire  s_163_6,  s_163_7,  s_163_8,  s_163_9, s_163_10, s_163_11;
wire s_163_12, s_163_13, s_163_14, s_163_15, s_163_16, s_163_17;
wire s_163_18, s_163_19, s_163_20, s_163_21, s_163_22, s_163_23;
wire s_163_24, s_163_25, s_163_26, s_163_27, s_163_28, s_163_29;
wire s_163_30, s_163_31, s_163_32, s_163_33, s_163_34, s_163_35;
wire s_163_36, s_163_37, s_163_38, s_163_39, s_163_40, s_163_41;
wire s_163_42, s_163_43, s_163_44, s_163_45, s_163_46, s_163_47;
wire  s_164_0,  s_164_1,  s_164_2,  s_164_3,  s_164_4,  s_164_5;
wire  s_164_6,  s_164_7,  s_164_8,  s_164_9, s_164_10, s_164_11;
wire s_164_12, s_164_13, s_164_14, s_164_15, s_164_16, s_164_17;
wire s_164_18, s_164_19, s_164_20, s_164_21, s_164_22, s_164_23;
wire s_164_24, s_164_25, s_164_26, s_164_27, s_164_28, s_164_29;
wire s_164_30, s_164_31, s_164_32, s_164_33, s_164_34, s_164_35;
wire s_164_36, s_164_37, s_164_38, s_164_39, s_164_40, s_164_41;
wire s_164_42, s_164_43, s_164_44, s_164_45, s_164_46,  s_165_0;
wire  s_165_1,  s_165_2,  s_165_3,  s_165_4,  s_165_5,  s_165_6;
wire  s_165_7,  s_165_8,  s_165_9, s_165_10, s_165_11, s_165_12;
wire s_165_13, s_165_14, s_165_15, s_165_16, s_165_17, s_165_18;
wire s_165_19, s_165_20, s_165_21, s_165_22, s_165_23, s_165_24;
wire s_165_25, s_165_26, s_165_27, s_165_28, s_165_29, s_165_30;
wire s_165_31, s_165_32, s_165_33, s_165_34, s_165_35, s_165_36;
wire s_165_37, s_165_38, s_165_39, s_165_40, s_165_41, s_165_42;
wire s_165_43, s_165_44, s_165_45, s_165_46,  s_166_0,  s_166_1;
wire  s_166_2,  s_166_3,  s_166_4,  s_166_5,  s_166_6,  s_166_7;
wire  s_166_8,  s_166_9, s_166_10, s_166_11, s_166_12, s_166_13;
wire s_166_14, s_166_15, s_166_16, s_166_17, s_166_18, s_166_19;
wire s_166_20, s_166_21, s_166_22, s_166_23, s_166_24, s_166_25;
wire s_166_26, s_166_27, s_166_28, s_166_29, s_166_30, s_166_31;
wire s_166_32, s_166_33, s_166_34, s_166_35, s_166_36, s_166_37;
wire s_166_38, s_166_39, s_166_40, s_166_41, s_166_42, s_166_43;
wire s_166_44, s_166_45,  s_167_0,  s_167_1,  s_167_2,  s_167_3;
wire  s_167_4,  s_167_5,  s_167_6,  s_167_7,  s_167_8,  s_167_9;
wire s_167_10, s_167_11, s_167_12, s_167_13, s_167_14, s_167_15;
wire s_167_16, s_167_17, s_167_18, s_167_19, s_167_20, s_167_21;
wire s_167_22, s_167_23, s_167_24, s_167_25, s_167_26, s_167_27;
wire s_167_28, s_167_29, s_167_30, s_167_31, s_167_32, s_167_33;
wire s_167_34, s_167_35, s_167_36, s_167_37, s_167_38, s_167_39;
wire s_167_40, s_167_41, s_167_42, s_167_43, s_167_44, s_167_45;
wire  s_168_0,  s_168_1,  s_168_2,  s_168_3,  s_168_4,  s_168_5;
wire  s_168_6,  s_168_7,  s_168_8,  s_168_9, s_168_10, s_168_11;
wire s_168_12, s_168_13, s_168_14, s_168_15, s_168_16, s_168_17;
wire s_168_18, s_168_19, s_168_20, s_168_21, s_168_22, s_168_23;
wire s_168_24, s_168_25, s_168_26, s_168_27, s_168_28, s_168_29;
wire s_168_30, s_168_31, s_168_32, s_168_33, s_168_34, s_168_35;
wire s_168_36, s_168_37, s_168_38, s_168_39, s_168_40, s_168_41;
wire s_168_42, s_168_43, s_168_44,  s_169_0,  s_169_1,  s_169_2;
wire  s_169_3,  s_169_4,  s_169_5,  s_169_6,  s_169_7,  s_169_8;
wire  s_169_9, s_169_10, s_169_11, s_169_12, s_169_13, s_169_14;
wire s_169_15, s_169_16, s_169_17, s_169_18, s_169_19, s_169_20;
wire s_169_21, s_169_22, s_169_23, s_169_24, s_169_25, s_169_26;
wire s_169_27, s_169_28, s_169_29, s_169_30, s_169_31, s_169_32;
wire s_169_33, s_169_34, s_169_35, s_169_36, s_169_37, s_169_38;
wire s_169_39, s_169_40, s_169_41, s_169_42, s_169_43, s_169_44;
wire  s_170_0,  s_170_1,  s_170_2,  s_170_3,  s_170_4,  s_170_5;
wire  s_170_6,  s_170_7,  s_170_8,  s_170_9, s_170_10, s_170_11;
wire s_170_12, s_170_13, s_170_14, s_170_15, s_170_16, s_170_17;
wire s_170_18, s_170_19, s_170_20, s_170_21, s_170_22, s_170_23;
wire s_170_24, s_170_25, s_170_26, s_170_27, s_170_28, s_170_29;
wire s_170_30, s_170_31, s_170_32, s_170_33, s_170_34, s_170_35;
wire s_170_36, s_170_37, s_170_38, s_170_39, s_170_40, s_170_41;
wire s_170_42, s_170_43,  s_171_0,  s_171_1,  s_171_2,  s_171_3;
wire  s_171_4,  s_171_5,  s_171_6,  s_171_7,  s_171_8,  s_171_9;
wire s_171_10, s_171_11, s_171_12, s_171_13, s_171_14, s_171_15;
wire s_171_16, s_171_17, s_171_18, s_171_19, s_171_20, s_171_21;
wire s_171_22, s_171_23, s_171_24, s_171_25, s_171_26, s_171_27;
wire s_171_28, s_171_29, s_171_30, s_171_31, s_171_32, s_171_33;
wire s_171_34, s_171_35, s_171_36, s_171_37, s_171_38, s_171_39;
wire s_171_40, s_171_41, s_171_42, s_171_43,  s_172_0,  s_172_1;
wire  s_172_2,  s_172_3,  s_172_4,  s_172_5,  s_172_6,  s_172_7;
wire  s_172_8,  s_172_9, s_172_10, s_172_11, s_172_12, s_172_13;
wire s_172_14, s_172_15, s_172_16, s_172_17, s_172_18, s_172_19;
wire s_172_20, s_172_21, s_172_22, s_172_23, s_172_24, s_172_25;
wire s_172_26, s_172_27, s_172_28, s_172_29, s_172_30, s_172_31;
wire s_172_32, s_172_33, s_172_34, s_172_35, s_172_36, s_172_37;
wire s_172_38, s_172_39, s_172_40, s_172_41, s_172_42,  s_173_0;
wire  s_173_1,  s_173_2,  s_173_3,  s_173_4,  s_173_5,  s_173_6;
wire  s_173_7,  s_173_8,  s_173_9, s_173_10, s_173_11, s_173_12;
wire s_173_13, s_173_14, s_173_15, s_173_16, s_173_17, s_173_18;
wire s_173_19, s_173_20, s_173_21, s_173_22, s_173_23, s_173_24;
wire s_173_25, s_173_26, s_173_27, s_173_28, s_173_29, s_173_30;
wire s_173_31, s_173_32, s_173_33, s_173_34, s_173_35, s_173_36;
wire s_173_37, s_173_38, s_173_39, s_173_40, s_173_41, s_173_42;
wire  s_174_0,  s_174_1,  s_174_2,  s_174_3,  s_174_4,  s_174_5;
wire  s_174_6,  s_174_7,  s_174_8,  s_174_9, s_174_10, s_174_11;
wire s_174_12, s_174_13, s_174_14, s_174_15, s_174_16, s_174_17;
wire s_174_18, s_174_19, s_174_20, s_174_21, s_174_22, s_174_23;
wire s_174_24, s_174_25, s_174_26, s_174_27, s_174_28, s_174_29;
wire s_174_30, s_174_31, s_174_32, s_174_33, s_174_34, s_174_35;
wire s_174_36, s_174_37, s_174_38, s_174_39, s_174_40, s_174_41;
wire  s_175_0,  s_175_1,  s_175_2,  s_175_3,  s_175_4,  s_175_5;
wire  s_175_6,  s_175_7,  s_175_8,  s_175_9, s_175_10, s_175_11;
wire s_175_12, s_175_13, s_175_14, s_175_15, s_175_16, s_175_17;
wire s_175_18, s_175_19, s_175_20, s_175_21, s_175_22, s_175_23;
wire s_175_24, s_175_25, s_175_26, s_175_27, s_175_28, s_175_29;
wire s_175_30, s_175_31, s_175_32, s_175_33, s_175_34, s_175_35;
wire s_175_36, s_175_37, s_175_38, s_175_39, s_175_40, s_175_41;
wire  s_176_0,  s_176_1,  s_176_2,  s_176_3,  s_176_4,  s_176_5;
wire  s_176_6,  s_176_7,  s_176_8,  s_176_9, s_176_10, s_176_11;
wire s_176_12, s_176_13, s_176_14, s_176_15, s_176_16, s_176_17;
wire s_176_18, s_176_19, s_176_20, s_176_21, s_176_22, s_176_23;
wire s_176_24, s_176_25, s_176_26, s_176_27, s_176_28, s_176_29;
wire s_176_30, s_176_31, s_176_32, s_176_33, s_176_34, s_176_35;
wire s_176_36, s_176_37, s_176_38, s_176_39, s_176_40,  s_177_0;
wire  s_177_1,  s_177_2,  s_177_3,  s_177_4,  s_177_5,  s_177_6;
wire  s_177_7,  s_177_8,  s_177_9, s_177_10, s_177_11, s_177_12;
wire s_177_13, s_177_14, s_177_15, s_177_16, s_177_17, s_177_18;
wire s_177_19, s_177_20, s_177_21, s_177_22, s_177_23, s_177_24;
wire s_177_25, s_177_26, s_177_27, s_177_28, s_177_29, s_177_30;
wire s_177_31, s_177_32, s_177_33, s_177_34, s_177_35, s_177_36;
wire s_177_37, s_177_38, s_177_39, s_177_40,  s_178_0,  s_178_1;
wire  s_178_2,  s_178_3,  s_178_4,  s_178_5,  s_178_6,  s_178_7;
wire  s_178_8,  s_178_9, s_178_10, s_178_11, s_178_12, s_178_13;
wire s_178_14, s_178_15, s_178_16, s_178_17, s_178_18, s_178_19;
wire s_178_20, s_178_21, s_178_22, s_178_23, s_178_24, s_178_25;
wire s_178_26, s_178_27, s_178_28, s_178_29, s_178_30, s_178_31;
wire s_178_32, s_178_33, s_178_34, s_178_35, s_178_36, s_178_37;
wire s_178_38, s_178_39,  s_179_0,  s_179_1,  s_179_2,  s_179_3;
wire  s_179_4,  s_179_5,  s_179_6,  s_179_7,  s_179_8,  s_179_9;
wire s_179_10, s_179_11, s_179_12, s_179_13, s_179_14, s_179_15;
wire s_179_16, s_179_17, s_179_18, s_179_19, s_179_20, s_179_21;
wire s_179_22, s_179_23, s_179_24, s_179_25, s_179_26, s_179_27;
wire s_179_28, s_179_29, s_179_30, s_179_31, s_179_32, s_179_33;
wire s_179_34, s_179_35, s_179_36, s_179_37, s_179_38, s_179_39;
wire  s_180_0,  s_180_1,  s_180_2,  s_180_3,  s_180_4,  s_180_5;
wire  s_180_6,  s_180_7,  s_180_8,  s_180_9, s_180_10, s_180_11;
wire s_180_12, s_180_13, s_180_14, s_180_15, s_180_16, s_180_17;
wire s_180_18, s_180_19, s_180_20, s_180_21, s_180_22, s_180_23;
wire s_180_24, s_180_25, s_180_26, s_180_27, s_180_28, s_180_29;
wire s_180_30, s_180_31, s_180_32, s_180_33, s_180_34, s_180_35;
wire s_180_36, s_180_37, s_180_38,  s_181_0,  s_181_1,  s_181_2;
wire  s_181_3,  s_181_4,  s_181_5,  s_181_6,  s_181_7,  s_181_8;
wire  s_181_9, s_181_10, s_181_11, s_181_12, s_181_13, s_181_14;
wire s_181_15, s_181_16, s_181_17, s_181_18, s_181_19, s_181_20;
wire s_181_21, s_181_22, s_181_23, s_181_24, s_181_25, s_181_26;
wire s_181_27, s_181_28, s_181_29, s_181_30, s_181_31, s_181_32;
wire s_181_33, s_181_34, s_181_35, s_181_36, s_181_37, s_181_38;
wire  s_182_0,  s_182_1,  s_182_2,  s_182_3,  s_182_4,  s_182_5;
wire  s_182_6,  s_182_7,  s_182_8,  s_182_9, s_182_10, s_182_11;
wire s_182_12, s_182_13, s_182_14, s_182_15, s_182_16, s_182_17;
wire s_182_18, s_182_19, s_182_20, s_182_21, s_182_22, s_182_23;
wire s_182_24, s_182_25, s_182_26, s_182_27, s_182_28, s_182_29;
wire s_182_30, s_182_31, s_182_32, s_182_33, s_182_34, s_182_35;
wire s_182_36, s_182_37,  s_183_0,  s_183_1,  s_183_2,  s_183_3;
wire  s_183_4,  s_183_5,  s_183_6,  s_183_7,  s_183_8,  s_183_9;
wire s_183_10, s_183_11, s_183_12, s_183_13, s_183_14, s_183_15;
wire s_183_16, s_183_17, s_183_18, s_183_19, s_183_20, s_183_21;
wire s_183_22, s_183_23, s_183_24, s_183_25, s_183_26, s_183_27;
wire s_183_28, s_183_29, s_183_30, s_183_31, s_183_32, s_183_33;
wire s_183_34, s_183_35, s_183_36, s_183_37,  s_184_0,  s_184_1;
wire  s_184_2,  s_184_3,  s_184_4,  s_184_5,  s_184_6,  s_184_7;
wire  s_184_8,  s_184_9, s_184_10, s_184_11, s_184_12, s_184_13;
wire s_184_14, s_184_15, s_184_16, s_184_17, s_184_18, s_184_19;
wire s_184_20, s_184_21, s_184_22, s_184_23, s_184_24, s_184_25;
wire s_184_26, s_184_27, s_184_28, s_184_29, s_184_30, s_184_31;
wire s_184_32, s_184_33, s_184_34, s_184_35, s_184_36,  s_185_0;
wire  s_185_1,  s_185_2,  s_185_3,  s_185_4,  s_185_5,  s_185_6;
wire  s_185_7,  s_185_8,  s_185_9, s_185_10, s_185_11, s_185_12;
wire s_185_13, s_185_14, s_185_15, s_185_16, s_185_17, s_185_18;
wire s_185_19, s_185_20, s_185_21, s_185_22, s_185_23, s_185_24;
wire s_185_25, s_185_26, s_185_27, s_185_28, s_185_29, s_185_30;
wire s_185_31, s_185_32, s_185_33, s_185_34, s_185_35, s_185_36;
wire  s_186_0,  s_186_1,  s_186_2,  s_186_3,  s_186_4,  s_186_5;
wire  s_186_6,  s_186_7,  s_186_8,  s_186_9, s_186_10, s_186_11;
wire s_186_12, s_186_13, s_186_14, s_186_15, s_186_16, s_186_17;
wire s_186_18, s_186_19, s_186_20, s_186_21, s_186_22, s_186_23;
wire s_186_24, s_186_25, s_186_26, s_186_27, s_186_28, s_186_29;
wire s_186_30, s_186_31, s_186_32, s_186_33, s_186_34, s_186_35;
wire  s_187_0,  s_187_1,  s_187_2,  s_187_3,  s_187_4,  s_187_5;
wire  s_187_6,  s_187_7,  s_187_8,  s_187_9, s_187_10, s_187_11;
wire s_187_12, s_187_13, s_187_14, s_187_15, s_187_16, s_187_17;
wire s_187_18, s_187_19, s_187_20, s_187_21, s_187_22, s_187_23;
wire s_187_24, s_187_25, s_187_26, s_187_27, s_187_28, s_187_29;
wire s_187_30, s_187_31, s_187_32, s_187_33, s_187_34, s_187_35;
wire  s_188_0,  s_188_1,  s_188_2,  s_188_3,  s_188_4,  s_188_5;
wire  s_188_6,  s_188_7,  s_188_8,  s_188_9, s_188_10, s_188_11;
wire s_188_12, s_188_13, s_188_14, s_188_15, s_188_16, s_188_17;
wire s_188_18, s_188_19, s_188_20, s_188_21, s_188_22, s_188_23;
wire s_188_24, s_188_25, s_188_26, s_188_27, s_188_28, s_188_29;
wire s_188_30, s_188_31, s_188_32, s_188_33, s_188_34,  s_189_0;
wire  s_189_1,  s_189_2,  s_189_3,  s_189_4,  s_189_5,  s_189_6;
wire  s_189_7,  s_189_8,  s_189_9, s_189_10, s_189_11, s_189_12;
wire s_189_13, s_189_14, s_189_15, s_189_16, s_189_17, s_189_18;
wire s_189_19, s_189_20, s_189_21, s_189_22, s_189_23, s_189_24;
wire s_189_25, s_189_26, s_189_27, s_189_28, s_189_29, s_189_30;
wire s_189_31, s_189_32, s_189_33, s_189_34,  s_190_0,  s_190_1;
wire  s_190_2,  s_190_3,  s_190_4,  s_190_5,  s_190_6,  s_190_7;
wire  s_190_8,  s_190_9, s_190_10, s_190_11, s_190_12, s_190_13;
wire s_190_14, s_190_15, s_190_16, s_190_17, s_190_18, s_190_19;
wire s_190_20, s_190_21, s_190_22, s_190_23, s_190_24, s_190_25;
wire s_190_26, s_190_27, s_190_28, s_190_29, s_190_30, s_190_31;
wire s_190_32, s_190_33,  s_191_0,  s_191_1,  s_191_2,  s_191_3;
wire  s_191_4,  s_191_5,  s_191_6,  s_191_7,  s_191_8,  s_191_9;
wire s_191_10, s_191_11, s_191_12, s_191_13, s_191_14, s_191_15;
wire s_191_16, s_191_17, s_191_18, s_191_19, s_191_20, s_191_21;
wire s_191_22, s_191_23, s_191_24, s_191_25, s_191_26, s_191_27;
wire s_191_28, s_191_29, s_191_30, s_191_31, s_191_32, s_191_33;
wire  s_192_0,  s_192_1,  s_192_2,  s_192_3,  s_192_4,  s_192_5;
wire  s_192_6,  s_192_7,  s_192_8,  s_192_9, s_192_10, s_192_11;
wire s_192_12, s_192_13, s_192_14, s_192_15, s_192_16, s_192_17;
wire s_192_18, s_192_19, s_192_20, s_192_21, s_192_22, s_192_23;
wire s_192_24, s_192_25, s_192_26, s_192_27, s_192_28, s_192_29;
wire s_192_30, s_192_31, s_192_32,  s_193_0,  s_193_1,  s_193_2;
wire  s_193_3,  s_193_4,  s_193_5,  s_193_6,  s_193_7,  s_193_8;
wire  s_193_9, s_193_10, s_193_11, s_193_12, s_193_13, s_193_14;
wire s_193_15, s_193_16, s_193_17, s_193_18, s_193_19, s_193_20;
wire s_193_21, s_193_22, s_193_23, s_193_24, s_193_25, s_193_26;
wire s_193_27, s_193_28, s_193_29, s_193_30, s_193_31, s_193_32;
wire  s_194_0,  s_194_1,  s_194_2,  s_194_3,  s_194_4,  s_194_5;
wire  s_194_6,  s_194_7,  s_194_8,  s_194_9, s_194_10, s_194_11;
wire s_194_12, s_194_13, s_194_14, s_194_15, s_194_16, s_194_17;
wire s_194_18, s_194_19, s_194_20, s_194_21, s_194_22, s_194_23;
wire s_194_24, s_194_25, s_194_26, s_194_27, s_194_28, s_194_29;
wire s_194_30, s_194_31,  s_195_0,  s_195_1,  s_195_2,  s_195_3;
wire  s_195_4,  s_195_5,  s_195_6,  s_195_7,  s_195_8,  s_195_9;
wire s_195_10, s_195_11, s_195_12, s_195_13, s_195_14, s_195_15;
wire s_195_16, s_195_17, s_195_18, s_195_19, s_195_20, s_195_21;
wire s_195_22, s_195_23, s_195_24, s_195_25, s_195_26, s_195_27;
wire s_195_28, s_195_29, s_195_30, s_195_31,  s_196_0,  s_196_1;
wire  s_196_2,  s_196_3,  s_196_4,  s_196_5,  s_196_6,  s_196_7;
wire  s_196_8,  s_196_9, s_196_10, s_196_11, s_196_12, s_196_13;
wire s_196_14, s_196_15, s_196_16, s_196_17, s_196_18, s_196_19;
wire s_196_20, s_196_21, s_196_22, s_196_23, s_196_24, s_196_25;
wire s_196_26, s_196_27, s_196_28, s_196_29, s_196_30,  s_197_0;
wire  s_197_1,  s_197_2,  s_197_3,  s_197_4,  s_197_5,  s_197_6;
wire  s_197_7,  s_197_8,  s_197_9, s_197_10, s_197_11, s_197_12;
wire s_197_13, s_197_14, s_197_15, s_197_16, s_197_17, s_197_18;
wire s_197_19, s_197_20, s_197_21, s_197_22, s_197_23, s_197_24;
wire s_197_25, s_197_26, s_197_27, s_197_28, s_197_29, s_197_30;
wire  s_198_0,  s_198_1,  s_198_2,  s_198_3,  s_198_4,  s_198_5;
wire  s_198_6,  s_198_7,  s_198_8,  s_198_9, s_198_10, s_198_11;
wire s_198_12, s_198_13, s_198_14, s_198_15, s_198_16, s_198_17;
wire s_198_18, s_198_19, s_198_20, s_198_21, s_198_22, s_198_23;
wire s_198_24, s_198_25, s_198_26, s_198_27, s_198_28, s_198_29;
wire  s_199_0,  s_199_1,  s_199_2,  s_199_3,  s_199_4,  s_199_5;
wire  s_199_6,  s_199_7,  s_199_8,  s_199_9, s_199_10, s_199_11;
wire s_199_12, s_199_13, s_199_14, s_199_15, s_199_16, s_199_17;
wire s_199_18, s_199_19, s_199_20, s_199_21, s_199_22, s_199_23;
wire s_199_24, s_199_25, s_199_26, s_199_27, s_199_28, s_199_29;
wire  s_200_0,  s_200_1,  s_200_2,  s_200_3,  s_200_4,  s_200_5;
wire  s_200_6,  s_200_7,  s_200_8,  s_200_9, s_200_10, s_200_11;
wire s_200_12, s_200_13, s_200_14, s_200_15, s_200_16, s_200_17;
wire s_200_18, s_200_19, s_200_20, s_200_21, s_200_22, s_200_23;
wire s_200_24, s_200_25, s_200_26, s_200_27, s_200_28,  s_201_0;
wire  s_201_1,  s_201_2,  s_201_3,  s_201_4,  s_201_5,  s_201_6;
wire  s_201_7,  s_201_8,  s_201_9, s_201_10, s_201_11, s_201_12;
wire s_201_13, s_201_14, s_201_15, s_201_16, s_201_17, s_201_18;
wire s_201_19, s_201_20, s_201_21, s_201_22, s_201_23, s_201_24;
wire s_201_25, s_201_26, s_201_27, s_201_28,  s_202_0,  s_202_1;
wire  s_202_2,  s_202_3,  s_202_4,  s_202_5,  s_202_6,  s_202_7;
wire  s_202_8,  s_202_9, s_202_10, s_202_11, s_202_12, s_202_13;
wire s_202_14, s_202_15, s_202_16, s_202_17, s_202_18, s_202_19;
wire s_202_20, s_202_21, s_202_22, s_202_23, s_202_24, s_202_25;
wire s_202_26, s_202_27,  s_203_0,  s_203_1,  s_203_2,  s_203_3;
wire  s_203_4,  s_203_5,  s_203_6,  s_203_7,  s_203_8,  s_203_9;
wire s_203_10, s_203_11, s_203_12, s_203_13, s_203_14, s_203_15;
wire s_203_16, s_203_17, s_203_18, s_203_19, s_203_20, s_203_21;
wire s_203_22, s_203_23, s_203_24, s_203_25, s_203_26, s_203_27;
wire  s_204_0,  s_204_1,  s_204_2,  s_204_3,  s_204_4,  s_204_5;
wire  s_204_6,  s_204_7,  s_204_8,  s_204_9, s_204_10, s_204_11;
wire s_204_12, s_204_13, s_204_14, s_204_15, s_204_16, s_204_17;
wire s_204_18, s_204_19, s_204_20, s_204_21, s_204_22, s_204_23;
wire s_204_24, s_204_25, s_204_26,  s_205_0,  s_205_1,  s_205_2;
wire  s_205_3,  s_205_4,  s_205_5,  s_205_6,  s_205_7,  s_205_8;
wire  s_205_9, s_205_10, s_205_11, s_205_12, s_205_13, s_205_14;
wire s_205_15, s_205_16, s_205_17, s_205_18, s_205_19, s_205_20;
wire s_205_21, s_205_22, s_205_23, s_205_24, s_205_25, s_205_26;
wire  s_206_0,  s_206_1,  s_206_2,  s_206_3,  s_206_4,  s_206_5;
wire  s_206_6,  s_206_7,  s_206_8,  s_206_9, s_206_10, s_206_11;
wire s_206_12, s_206_13, s_206_14, s_206_15, s_206_16, s_206_17;
wire s_206_18, s_206_19, s_206_20, s_206_21, s_206_22, s_206_23;
wire s_206_24, s_206_25,  s_207_0,  s_207_1,  s_207_2,  s_207_3;
wire  s_207_4,  s_207_5,  s_207_6,  s_207_7,  s_207_8,  s_207_9;
wire s_207_10, s_207_11, s_207_12, s_207_13, s_207_14, s_207_15;
wire s_207_16, s_207_17, s_207_18, s_207_19, s_207_20, s_207_21;
wire s_207_22, s_207_23, s_207_24, s_207_25,  s_208_0,  s_208_1;
wire  s_208_2,  s_208_3,  s_208_4,  s_208_5,  s_208_6,  s_208_7;
wire  s_208_8,  s_208_9, s_208_10, s_208_11, s_208_12, s_208_13;
wire s_208_14, s_208_15, s_208_16, s_208_17, s_208_18, s_208_19;
wire s_208_20, s_208_21, s_208_22, s_208_23, s_208_24,  s_209_0;
wire  s_209_1,  s_209_2,  s_209_3,  s_209_4,  s_209_5,  s_209_6;
wire  s_209_7,  s_209_8,  s_209_9, s_209_10, s_209_11, s_209_12;
wire s_209_13, s_209_14, s_209_15, s_209_16, s_209_17, s_209_18;
wire s_209_19, s_209_20, s_209_21, s_209_22, s_209_23, s_209_24;
wire  s_210_0,  s_210_1,  s_210_2,  s_210_3,  s_210_4,  s_210_5;
wire  s_210_6,  s_210_7,  s_210_8,  s_210_9, s_210_10, s_210_11;
wire s_210_12, s_210_13, s_210_14, s_210_15, s_210_16, s_210_17;
wire s_210_18, s_210_19, s_210_20, s_210_21, s_210_22, s_210_23;
wire  s_211_0,  s_211_1,  s_211_2,  s_211_3,  s_211_4,  s_211_5;
wire  s_211_6,  s_211_7,  s_211_8,  s_211_9, s_211_10, s_211_11;
wire s_211_12, s_211_13, s_211_14, s_211_15, s_211_16, s_211_17;
wire s_211_18, s_211_19, s_211_20, s_211_21, s_211_22, s_211_23;
wire  s_212_0,  s_212_1,  s_212_2,  s_212_3,  s_212_4,  s_212_5;
wire  s_212_6,  s_212_7,  s_212_8,  s_212_9, s_212_10, s_212_11;
wire s_212_12, s_212_13, s_212_14, s_212_15, s_212_16, s_212_17;
wire s_212_18, s_212_19, s_212_20, s_212_21, s_212_22,  s_213_0;
wire  s_213_1,  s_213_2,  s_213_3,  s_213_4,  s_213_5,  s_213_6;
wire  s_213_7,  s_213_8,  s_213_9, s_213_10, s_213_11, s_213_12;
wire s_213_13, s_213_14, s_213_15, s_213_16, s_213_17, s_213_18;
wire s_213_19, s_213_20, s_213_21, s_213_22,  s_214_0,  s_214_1;
wire  s_214_2,  s_214_3,  s_214_4,  s_214_5,  s_214_6,  s_214_7;
wire  s_214_8,  s_214_9, s_214_10, s_214_11, s_214_12, s_214_13;
wire s_214_14, s_214_15, s_214_16, s_214_17, s_214_18, s_214_19;
wire s_214_20, s_214_21,  s_215_0,  s_215_1,  s_215_2,  s_215_3;
wire  s_215_4,  s_215_5,  s_215_6,  s_215_7,  s_215_8,  s_215_9;
wire s_215_10, s_215_11, s_215_12, s_215_13, s_215_14, s_215_15;
wire s_215_16, s_215_17, s_215_18, s_215_19, s_215_20, s_215_21;
wire  s_216_0,  s_216_1,  s_216_2,  s_216_3,  s_216_4,  s_216_5;
wire  s_216_6,  s_216_7,  s_216_8,  s_216_9, s_216_10, s_216_11;
wire s_216_12, s_216_13, s_216_14, s_216_15, s_216_16, s_216_17;
wire s_216_18, s_216_19, s_216_20,  s_217_0,  s_217_1,  s_217_2;
wire  s_217_3,  s_217_4,  s_217_5,  s_217_6,  s_217_7,  s_217_8;
wire  s_217_9, s_217_10, s_217_11, s_217_12, s_217_13, s_217_14;
wire s_217_15, s_217_16, s_217_17, s_217_18, s_217_19, s_217_20;
wire  s_218_0,  s_218_1,  s_218_2,  s_218_3,  s_218_4,  s_218_5;
wire  s_218_6,  s_218_7,  s_218_8,  s_218_9, s_218_10, s_218_11;
wire s_218_12, s_218_13, s_218_14, s_218_15, s_218_16, s_218_17;
wire s_218_18, s_218_19,  s_219_0,  s_219_1,  s_219_2,  s_219_3;
wire  s_219_4,  s_219_5,  s_219_6,  s_219_7,  s_219_8,  s_219_9;
wire s_219_10, s_219_11, s_219_12, s_219_13, s_219_14, s_219_15;
wire s_219_16, s_219_17, s_219_18, s_219_19,  s_220_0,  s_220_1;
wire  s_220_2,  s_220_3,  s_220_4,  s_220_5,  s_220_6,  s_220_7;
wire  s_220_8,  s_220_9, s_220_10, s_220_11, s_220_12, s_220_13;
wire s_220_14, s_220_15, s_220_16, s_220_17, s_220_18,  s_221_0;
wire  s_221_1,  s_221_2,  s_221_3,  s_221_4,  s_221_5,  s_221_6;
wire  s_221_7,  s_221_8,  s_221_9, s_221_10, s_221_11, s_221_12;
wire s_221_13, s_221_14, s_221_15, s_221_16, s_221_17, s_221_18;
wire  s_222_0,  s_222_1,  s_222_2,  s_222_3,  s_222_4,  s_222_5;
wire  s_222_6,  s_222_7,  s_222_8,  s_222_9, s_222_10, s_222_11;
wire s_222_12, s_222_13, s_222_14, s_222_15, s_222_16, s_222_17;
wire  s_223_0,  s_223_1,  s_223_2,  s_223_3,  s_223_4,  s_223_5;
wire  s_223_6,  s_223_7,  s_223_8,  s_223_9, s_223_10, s_223_11;
wire s_223_12, s_223_13, s_223_14, s_223_15, s_223_16, s_223_17;
wire  s_224_0,  s_224_1,  s_224_2,  s_224_3,  s_224_4,  s_224_5;
wire  s_224_6,  s_224_7,  s_224_8,  s_224_9, s_224_10, s_224_11;
wire s_224_12, s_224_13, s_224_14, s_224_15, s_224_16,  s_225_0;
wire  s_225_1,  s_225_2,  s_225_3,  s_225_4,  s_225_5,  s_225_6;
wire  s_225_7,  s_225_8,  s_225_9, s_225_10, s_225_11, s_225_12;
wire s_225_13, s_225_14, s_225_15, s_225_16,  s_226_0,  s_226_1;
wire  s_226_2,  s_226_3,  s_226_4,  s_226_5,  s_226_6,  s_226_7;
wire  s_226_8,  s_226_9, s_226_10, s_226_11, s_226_12, s_226_13;
wire s_226_14, s_226_15,  s_227_0,  s_227_1,  s_227_2,  s_227_3;
wire  s_227_4,  s_227_5,  s_227_6,  s_227_7,  s_227_8,  s_227_9;
wire s_227_10, s_227_11, s_227_12, s_227_13, s_227_14, s_227_15;
wire  s_228_0,  s_228_1,  s_228_2,  s_228_3,  s_228_4,  s_228_5;
wire  s_228_6,  s_228_7,  s_228_8,  s_228_9, s_228_10, s_228_11;
wire s_228_12, s_228_13, s_228_14,  s_229_0,  s_229_1,  s_229_2;
wire  s_229_3,  s_229_4,  s_229_5,  s_229_6,  s_229_7,  s_229_8;
wire  s_229_9, s_229_10, s_229_11, s_229_12, s_229_13, s_229_14;
wire  s_230_0,  s_230_1,  s_230_2,  s_230_3,  s_230_4,  s_230_5;
wire  s_230_6,  s_230_7,  s_230_8,  s_230_9, s_230_10, s_230_11;
wire s_230_12, s_230_13,  s_231_0,  s_231_1,  s_231_2,  s_231_3;
wire  s_231_4,  s_231_5,  s_231_6,  s_231_7,  s_231_8,  s_231_9;
wire s_231_10, s_231_11, s_231_12, s_231_13,  s_232_0,  s_232_1;
wire  s_232_2,  s_232_3,  s_232_4,  s_232_5,  s_232_6,  s_232_7;
wire  s_232_8,  s_232_9, s_232_10, s_232_11, s_232_12,  s_233_0;
wire  s_233_1,  s_233_2,  s_233_3,  s_233_4,  s_233_5,  s_233_6;
wire  s_233_7,  s_233_8,  s_233_9, s_233_10, s_233_11, s_233_12;
wire  s_234_0,  s_234_1,  s_234_2,  s_234_3,  s_234_4,  s_234_5;
wire  s_234_6,  s_234_7,  s_234_8,  s_234_9, s_234_10, s_234_11;
wire  s_235_0,  s_235_1,  s_235_2,  s_235_3,  s_235_4,  s_235_5;
wire  s_235_6,  s_235_7,  s_235_8,  s_235_9, s_235_10, s_235_11;
wire  s_236_0,  s_236_1,  s_236_2,  s_236_3,  s_236_4,  s_236_5;
wire  s_236_6,  s_236_7,  s_236_8,  s_236_9, s_236_10,  s_237_0;
wire  s_237_1,  s_237_2,  s_237_3,  s_237_4,  s_237_5,  s_237_6;
wire  s_237_7,  s_237_8,  s_237_9, s_237_10,  s_238_0,  s_238_1;
wire  s_238_2,  s_238_3,  s_238_4,  s_238_5,  s_238_6,  s_238_7;
wire  s_238_8,  s_238_9,  s_239_0,  s_239_1,  s_239_2,  s_239_3;
wire  s_239_4,  s_239_5,  s_239_6,  s_239_7,  s_239_8,  s_239_9;
wire  s_240_0,  s_240_1,  s_240_2,  s_240_3,  s_240_4,  s_240_5;
wire  s_240_6,  s_240_7,  s_240_8,  s_241_0,  s_241_1,  s_241_2;
wire  s_241_3,  s_241_4,  s_241_5,  s_241_6,  s_241_7,  s_241_8;
wire  s_242_0,  s_242_1,  s_242_2,  s_242_3,  s_242_4,  s_242_5;
wire  s_242_6,  s_242_7,  s_243_0,  s_243_1,  s_243_2,  s_243_3;
wire  s_243_4,  s_243_5,  s_243_6,  s_243_7,  s_244_0,  s_244_1;
wire  s_244_2,  s_244_3,  s_244_4,  s_244_5,  s_244_6,  s_245_0;
wire  s_245_1,  s_245_2,  s_245_3,  s_245_4,  s_245_5,  s_245_6;
wire  s_246_0,  s_246_1,  s_246_2,  s_246_3,  s_246_4,  s_246_5;
wire  s_247_0,  s_247_1,  s_247_2,  s_247_3,  s_247_4,  s_247_5;
wire  s_248_0,  s_248_1,  s_248_2,  s_248_3,  s_248_4,  s_249_0;
wire  s_249_1,  s_249_2,  s_249_3,  s_249_4,  s_250_0,  s_250_1;
wire  s_250_2,  s_250_3,  s_251_0,  s_251_1,  s_251_2,  s_251_3;
wire  s_252_0,  s_252_1,  s_252_2,  s_253_0,  s_253_1,  s_253_2;
wire  s_254_0,  s_254_1,  s_255_0,  s_255_1;

assign {
s_126_64, s_124_63, s_122_62, s_120_61, s_118_60, s_116_59, 
s_114_58, s_112_57, s_110_56, s_108_55, s_106_54, s_104_53, 
s_102_52, s_100_51,  s_98_50,  s_96_49,  s_94_48,  s_92_47, 
 s_90_46,  s_88_45,  s_86_44,  s_84_43,  s_82_42,  s_80_41, 
 s_78_40,  s_76_39,  s_74_38,  s_72_37,  s_70_36,  s_68_35, 
 s_66_34,  s_64_33,  s_62_32,  s_60_31,  s_58_30,  s_56_29, 
 s_54_28,  s_52_27,  s_50_26,  s_48_25,  s_46_24,  s_44_23, 
 s_42_22,  s_40_21,  s_38_20,  s_36_19,  s_34_18,  s_32_17, 
 s_30_16,  s_28_15,  s_26_14,  s_24_13,  s_22_12,  s_20_11, 
 s_18_10,   s_16_9,   s_14_8,   s_12_7,   s_10_6,    s_8_5, 
   s_6_4,    s_4_3,    s_2_2,    s_0_1
} = carry;

assign {
 s_129_0,  s_128_0,  s_127_0,  s_126_0,  s_125_0,  s_124_0, 
 s_123_0,  s_122_0,  s_121_0,  s_120_0,  s_119_0,  s_118_0, 
 s_117_0,  s_116_0,  s_115_0,  s_114_0,  s_113_0,  s_112_0, 
 s_111_0,  s_110_0,  s_109_0,  s_108_0,  s_107_0,  s_106_0, 
 s_105_0,  s_104_0,  s_103_0,  s_102_0,  s_101_0,  s_100_0, 
  s_99_0,   s_98_0,   s_97_0,   s_96_0,   s_95_0,   s_94_0, 
  s_93_0,   s_92_0,   s_91_0,   s_90_0,   s_89_0,   s_88_0, 
  s_87_0,   s_86_0,   s_85_0,   s_84_0,   s_83_0,   s_82_0, 
  s_81_0,   s_80_0,   s_79_0,   s_78_0,   s_77_0,   s_76_0, 
  s_75_0,   s_74_0,   s_73_0,   s_72_0,   s_71_0,   s_70_0, 
  s_69_0,   s_68_0,   s_67_0,   s_66_0,   s_65_0,   s_64_0, 
  s_63_0,   s_62_0,   s_61_0,   s_60_0,   s_59_0,   s_58_0, 
  s_57_0,   s_56_0,   s_55_0,   s_54_0,   s_53_0,   s_52_0, 
  s_51_0,   s_50_0,   s_49_0,   s_48_0,   s_47_0,   s_46_0, 
  s_45_0,   s_44_0,   s_43_0,   s_42_0,   s_41_0,   s_40_0, 
  s_39_0,   s_38_0,   s_37_0,   s_36_0,   s_35_0,   s_34_0, 
  s_33_0,   s_32_0,   s_31_0,   s_30_0,   s_29_0,   s_28_0, 
  s_27_0,   s_26_0,   s_25_0,   s_24_0,   s_23_0,   s_22_0, 
  s_21_0,   s_20_0,   s_19_0,   s_18_0,   s_17_0,   s_16_0, 
  s_15_0,   s_14_0,   s_13_0,   s_12_0,   s_11_0,   s_10_0, 
   s_9_0,    s_8_0,    s_7_0,    s_6_0,    s_5_0,    s_4_0, 
   s_3_0,    s_2_0,    s_1_0,    s_0_0
} = partial_products[(width+2)*(0+1)-1:(width+2)*0];

assign {
 s_131_0,  s_130_0,  s_129_1,  s_128_1,  s_127_1,  s_126_1, 
 s_125_1,  s_124_1,  s_123_1,  s_122_1,  s_121_1,  s_120_1, 
 s_119_1,  s_118_1,  s_117_1,  s_116_1,  s_115_1,  s_114_1, 
 s_113_1,  s_112_1,  s_111_1,  s_110_1,  s_109_1,  s_108_1, 
 s_107_1,  s_106_1,  s_105_1,  s_104_1,  s_103_1,  s_102_1, 
 s_101_1,  s_100_1,   s_99_1,   s_98_1,   s_97_1,   s_96_1, 
  s_95_1,   s_94_1,   s_93_1,   s_92_1,   s_91_1,   s_90_1, 
  s_89_1,   s_88_1,   s_87_1,   s_86_1,   s_85_1,   s_84_1, 
  s_83_1,   s_82_1,   s_81_1,   s_80_1,   s_79_1,   s_78_1, 
  s_77_1,   s_76_1,   s_75_1,   s_74_1,   s_73_1,   s_72_1, 
  s_71_1,   s_70_1,   s_69_1,   s_68_1,   s_67_1,   s_66_1, 
  s_65_1,   s_64_1,   s_63_1,   s_62_1,   s_61_1,   s_60_1, 
  s_59_1,   s_58_1,   s_57_1,   s_56_1,   s_55_1,   s_54_1, 
  s_53_1,   s_52_1,   s_51_1,   s_50_1,   s_49_1,   s_48_1, 
  s_47_1,   s_46_1,   s_45_1,   s_44_1,   s_43_1,   s_42_1, 
  s_41_1,   s_40_1,   s_39_1,   s_38_1,   s_37_1,   s_36_1, 
  s_35_1,   s_34_1,   s_33_1,   s_32_1,   s_31_1,   s_30_1, 
  s_29_1,   s_28_1,   s_27_1,   s_26_1,   s_25_1,   s_24_1, 
  s_23_1,   s_22_1,   s_21_1,   s_20_1,   s_19_1,   s_18_1, 
  s_17_1,   s_16_1,   s_15_1,   s_14_1,   s_13_1,   s_12_1, 
  s_11_1,   s_10_1,    s_9_1,    s_8_1,    s_7_1,    s_6_1, 
   s_5_1,    s_4_1,    s_3_1,    s_2_1
} = partial_products[(width+2)*(1+1)-1:(width+2)*1];

assign {
 s_133_0,  s_132_0,  s_131_1,  s_130_1,  s_129_2,  s_128_2, 
 s_127_2,  s_126_2,  s_125_2,  s_124_2,  s_123_2,  s_122_2, 
 s_121_2,  s_120_2,  s_119_2,  s_118_2,  s_117_2,  s_116_2, 
 s_115_2,  s_114_2,  s_113_2,  s_112_2,  s_111_2,  s_110_2, 
 s_109_2,  s_108_2,  s_107_2,  s_106_2,  s_105_2,  s_104_2, 
 s_103_2,  s_102_2,  s_101_2,  s_100_2,   s_99_2,   s_98_2, 
  s_97_2,   s_96_2,   s_95_2,   s_94_2,   s_93_2,   s_92_2, 
  s_91_2,   s_90_2,   s_89_2,   s_88_2,   s_87_2,   s_86_2, 
  s_85_2,   s_84_2,   s_83_2,   s_82_2,   s_81_2,   s_80_2, 
  s_79_2,   s_78_2,   s_77_2,   s_76_2,   s_75_2,   s_74_2, 
  s_73_2,   s_72_2,   s_71_2,   s_70_2,   s_69_2,   s_68_2, 
  s_67_2,   s_66_2,   s_65_2,   s_64_2,   s_63_2,   s_62_2, 
  s_61_2,   s_60_2,   s_59_2,   s_58_2,   s_57_2,   s_56_2, 
  s_55_2,   s_54_2,   s_53_2,   s_52_2,   s_51_2,   s_50_2, 
  s_49_2,   s_48_2,   s_47_2,   s_46_2,   s_45_2,   s_44_2, 
  s_43_2,   s_42_2,   s_41_2,   s_40_2,   s_39_2,   s_38_2, 
  s_37_2,   s_36_2,   s_35_2,   s_34_2,   s_33_2,   s_32_2, 
  s_31_2,   s_30_2,   s_29_2,   s_28_2,   s_27_2,   s_26_2, 
  s_25_2,   s_24_2,   s_23_2,   s_22_2,   s_21_2,   s_20_2, 
  s_19_2,   s_18_2,   s_17_2,   s_16_2,   s_15_2,   s_14_2, 
  s_13_2,   s_12_2,   s_11_2,   s_10_2,    s_9_2,    s_8_2, 
   s_7_2,    s_6_2,    s_5_2,    s_4_2
} = partial_products[(width+2)*(2+1)-1:(width+2)*2];

assign {
 s_135_0,  s_134_0,  s_133_1,  s_132_1,  s_131_2,  s_130_2, 
 s_129_3,  s_128_3,  s_127_3,  s_126_3,  s_125_3,  s_124_3, 
 s_123_3,  s_122_3,  s_121_3,  s_120_3,  s_119_3,  s_118_3, 
 s_117_3,  s_116_3,  s_115_3,  s_114_3,  s_113_3,  s_112_3, 
 s_111_3,  s_110_3,  s_109_3,  s_108_3,  s_107_3,  s_106_3, 
 s_105_3,  s_104_3,  s_103_3,  s_102_3,  s_101_3,  s_100_3, 
  s_99_3,   s_98_3,   s_97_3,   s_96_3,   s_95_3,   s_94_3, 
  s_93_3,   s_92_3,   s_91_3,   s_90_3,   s_89_3,   s_88_3, 
  s_87_3,   s_86_3,   s_85_3,   s_84_3,   s_83_3,   s_82_3, 
  s_81_3,   s_80_3,   s_79_3,   s_78_3,   s_77_3,   s_76_3, 
  s_75_3,   s_74_3,   s_73_3,   s_72_3,   s_71_3,   s_70_3, 
  s_69_3,   s_68_3,   s_67_3,   s_66_3,   s_65_3,   s_64_3, 
  s_63_3,   s_62_3,   s_61_3,   s_60_3,   s_59_3,   s_58_3, 
  s_57_3,   s_56_3,   s_55_3,   s_54_3,   s_53_3,   s_52_3, 
  s_51_3,   s_50_3,   s_49_3,   s_48_3,   s_47_3,   s_46_3, 
  s_45_3,   s_44_3,   s_43_3,   s_42_3,   s_41_3,   s_40_3, 
  s_39_3,   s_38_3,   s_37_3,   s_36_3,   s_35_3,   s_34_3, 
  s_33_3,   s_32_3,   s_31_3,   s_30_3,   s_29_3,   s_28_3, 
  s_27_3,   s_26_3,   s_25_3,   s_24_3,   s_23_3,   s_22_3, 
  s_21_3,   s_20_3,   s_19_3,   s_18_3,   s_17_3,   s_16_3, 
  s_15_3,   s_14_3,   s_13_3,   s_12_3,   s_11_3,   s_10_3, 
   s_9_3,    s_8_3,    s_7_3,    s_6_3
} = partial_products[(width+2)*(3+1)-1:(width+2)*3];

assign {
 s_137_0,  s_136_0,  s_135_1,  s_134_1,  s_133_2,  s_132_2, 
 s_131_3,  s_130_3,  s_129_4,  s_128_4,  s_127_4,  s_126_4, 
 s_125_4,  s_124_4,  s_123_4,  s_122_4,  s_121_4,  s_120_4, 
 s_119_4,  s_118_4,  s_117_4,  s_116_4,  s_115_4,  s_114_4, 
 s_113_4,  s_112_4,  s_111_4,  s_110_4,  s_109_4,  s_108_4, 
 s_107_4,  s_106_4,  s_105_4,  s_104_4,  s_103_4,  s_102_4, 
 s_101_4,  s_100_4,   s_99_4,   s_98_4,   s_97_4,   s_96_4, 
  s_95_4,   s_94_4,   s_93_4,   s_92_4,   s_91_4,   s_90_4, 
  s_89_4,   s_88_4,   s_87_4,   s_86_4,   s_85_4,   s_84_4, 
  s_83_4,   s_82_4,   s_81_4,   s_80_4,   s_79_4,   s_78_4, 
  s_77_4,   s_76_4,   s_75_4,   s_74_4,   s_73_4,   s_72_4, 
  s_71_4,   s_70_4,   s_69_4,   s_68_4,   s_67_4,   s_66_4, 
  s_65_4,   s_64_4,   s_63_4,   s_62_4,   s_61_4,   s_60_4, 
  s_59_4,   s_58_4,   s_57_4,   s_56_4,   s_55_4,   s_54_4, 
  s_53_4,   s_52_4,   s_51_4,   s_50_4,   s_49_4,   s_48_4, 
  s_47_4,   s_46_4,   s_45_4,   s_44_4,   s_43_4,   s_42_4, 
  s_41_4,   s_40_4,   s_39_4,   s_38_4,   s_37_4,   s_36_4, 
  s_35_4,   s_34_4,   s_33_4,   s_32_4,   s_31_4,   s_30_4, 
  s_29_4,   s_28_4,   s_27_4,   s_26_4,   s_25_4,   s_24_4, 
  s_23_4,   s_22_4,   s_21_4,   s_20_4,   s_19_4,   s_18_4, 
  s_17_4,   s_16_4,   s_15_4,   s_14_4,   s_13_4,   s_12_4, 
  s_11_4,   s_10_4,    s_9_4,    s_8_4
} = partial_products[(width+2)*(4+1)-1:(width+2)*4];

assign {
 s_139_0,  s_138_0,  s_137_1,  s_136_1,  s_135_2,  s_134_2, 
 s_133_3,  s_132_3,  s_131_4,  s_130_4,  s_129_5,  s_128_5, 
 s_127_5,  s_126_5,  s_125_5,  s_124_5,  s_123_5,  s_122_5, 
 s_121_5,  s_120_5,  s_119_5,  s_118_5,  s_117_5,  s_116_5, 
 s_115_5,  s_114_5,  s_113_5,  s_112_5,  s_111_5,  s_110_5, 
 s_109_5,  s_108_5,  s_107_5,  s_106_5,  s_105_5,  s_104_5, 
 s_103_5,  s_102_5,  s_101_5,  s_100_5,   s_99_5,   s_98_5, 
  s_97_5,   s_96_5,   s_95_5,   s_94_5,   s_93_5,   s_92_5, 
  s_91_5,   s_90_5,   s_89_5,   s_88_5,   s_87_5,   s_86_5, 
  s_85_5,   s_84_5,   s_83_5,   s_82_5,   s_81_5,   s_80_5, 
  s_79_5,   s_78_5,   s_77_5,   s_76_5,   s_75_5,   s_74_5, 
  s_73_5,   s_72_5,   s_71_5,   s_70_5,   s_69_5,   s_68_5, 
  s_67_5,   s_66_5,   s_65_5,   s_64_5,   s_63_5,   s_62_5, 
  s_61_5,   s_60_5,   s_59_5,   s_58_5,   s_57_5,   s_56_5, 
  s_55_5,   s_54_5,   s_53_5,   s_52_5,   s_51_5,   s_50_5, 
  s_49_5,   s_48_5,   s_47_5,   s_46_5,   s_45_5,   s_44_5, 
  s_43_5,   s_42_5,   s_41_5,   s_40_5,   s_39_5,   s_38_5, 
  s_37_5,   s_36_5,   s_35_5,   s_34_5,   s_33_5,   s_32_5, 
  s_31_5,   s_30_5,   s_29_5,   s_28_5,   s_27_5,   s_26_5, 
  s_25_5,   s_24_5,   s_23_5,   s_22_5,   s_21_5,   s_20_5, 
  s_19_5,   s_18_5,   s_17_5,   s_16_5,   s_15_5,   s_14_5, 
  s_13_5,   s_12_5,   s_11_5,   s_10_5
} = partial_products[(width+2)*(5+1)-1:(width+2)*5];

assign {
 s_141_0,  s_140_0,  s_139_1,  s_138_1,  s_137_2,  s_136_2, 
 s_135_3,  s_134_3,  s_133_4,  s_132_4,  s_131_5,  s_130_5, 
 s_129_6,  s_128_6,  s_127_6,  s_126_6,  s_125_6,  s_124_6, 
 s_123_6,  s_122_6,  s_121_6,  s_120_6,  s_119_6,  s_118_6, 
 s_117_6,  s_116_6,  s_115_6,  s_114_6,  s_113_6,  s_112_6, 
 s_111_6,  s_110_6,  s_109_6,  s_108_6,  s_107_6,  s_106_6, 
 s_105_6,  s_104_6,  s_103_6,  s_102_6,  s_101_6,  s_100_6, 
  s_99_6,   s_98_6,   s_97_6,   s_96_6,   s_95_6,   s_94_6, 
  s_93_6,   s_92_6,   s_91_6,   s_90_6,   s_89_6,   s_88_6, 
  s_87_6,   s_86_6,   s_85_6,   s_84_6,   s_83_6,   s_82_6, 
  s_81_6,   s_80_6,   s_79_6,   s_78_6,   s_77_6,   s_76_6, 
  s_75_6,   s_74_6,   s_73_6,   s_72_6,   s_71_6,   s_70_6, 
  s_69_6,   s_68_6,   s_67_6,   s_66_6,   s_65_6,   s_64_6, 
  s_63_6,   s_62_6,   s_61_6,   s_60_6,   s_59_6,   s_58_6, 
  s_57_6,   s_56_6,   s_55_6,   s_54_6,   s_53_6,   s_52_6, 
  s_51_6,   s_50_6,   s_49_6,   s_48_6,   s_47_6,   s_46_6, 
  s_45_6,   s_44_6,   s_43_6,   s_42_6,   s_41_6,   s_40_6, 
  s_39_6,   s_38_6,   s_37_6,   s_36_6,   s_35_6,   s_34_6, 
  s_33_6,   s_32_6,   s_31_6,   s_30_6,   s_29_6,   s_28_6, 
  s_27_6,   s_26_6,   s_25_6,   s_24_6,   s_23_6,   s_22_6, 
  s_21_6,   s_20_6,   s_19_6,   s_18_6,   s_17_6,   s_16_6, 
  s_15_6,   s_14_6,   s_13_6,   s_12_6
} = partial_products[(width+2)*(6+1)-1:(width+2)*6];

assign {
 s_143_0,  s_142_0,  s_141_1,  s_140_1,  s_139_2,  s_138_2, 
 s_137_3,  s_136_3,  s_135_4,  s_134_4,  s_133_5,  s_132_5, 
 s_131_6,  s_130_6,  s_129_7,  s_128_7,  s_127_7,  s_126_7, 
 s_125_7,  s_124_7,  s_123_7,  s_122_7,  s_121_7,  s_120_7, 
 s_119_7,  s_118_7,  s_117_7,  s_116_7,  s_115_7,  s_114_7, 
 s_113_7,  s_112_7,  s_111_7,  s_110_7,  s_109_7,  s_108_7, 
 s_107_7,  s_106_7,  s_105_7,  s_104_7,  s_103_7,  s_102_7, 
 s_101_7,  s_100_7,   s_99_7,   s_98_7,   s_97_7,   s_96_7, 
  s_95_7,   s_94_7,   s_93_7,   s_92_7,   s_91_7,   s_90_7, 
  s_89_7,   s_88_7,   s_87_7,   s_86_7,   s_85_7,   s_84_7, 
  s_83_7,   s_82_7,   s_81_7,   s_80_7,   s_79_7,   s_78_7, 
  s_77_7,   s_76_7,   s_75_7,   s_74_7,   s_73_7,   s_72_7, 
  s_71_7,   s_70_7,   s_69_7,   s_68_7,   s_67_7,   s_66_7, 
  s_65_7,   s_64_7,   s_63_7,   s_62_7,   s_61_7,   s_60_7, 
  s_59_7,   s_58_7,   s_57_7,   s_56_7,   s_55_7,   s_54_7, 
  s_53_7,   s_52_7,   s_51_7,   s_50_7,   s_49_7,   s_48_7, 
  s_47_7,   s_46_7,   s_45_7,   s_44_7,   s_43_7,   s_42_7, 
  s_41_7,   s_40_7,   s_39_7,   s_38_7,   s_37_7,   s_36_7, 
  s_35_7,   s_34_7,   s_33_7,   s_32_7,   s_31_7,   s_30_7, 
  s_29_7,   s_28_7,   s_27_7,   s_26_7,   s_25_7,   s_24_7, 
  s_23_7,   s_22_7,   s_21_7,   s_20_7,   s_19_7,   s_18_7, 
  s_17_7,   s_16_7,   s_15_7,   s_14_7
} = partial_products[(width+2)*(7+1)-1:(width+2)*7];

assign {
 s_145_0,  s_144_0,  s_143_1,  s_142_1,  s_141_2,  s_140_2, 
 s_139_3,  s_138_3,  s_137_4,  s_136_4,  s_135_5,  s_134_5, 
 s_133_6,  s_132_6,  s_131_7,  s_130_7,  s_129_8,  s_128_8, 
 s_127_8,  s_126_8,  s_125_8,  s_124_8,  s_123_8,  s_122_8, 
 s_121_8,  s_120_8,  s_119_8,  s_118_8,  s_117_8,  s_116_8, 
 s_115_8,  s_114_8,  s_113_8,  s_112_8,  s_111_8,  s_110_8, 
 s_109_8,  s_108_8,  s_107_8,  s_106_8,  s_105_8,  s_104_8, 
 s_103_8,  s_102_8,  s_101_8,  s_100_8,   s_99_8,   s_98_8, 
  s_97_8,   s_96_8,   s_95_8,   s_94_8,   s_93_8,   s_92_8, 
  s_91_8,   s_90_8,   s_89_8,   s_88_8,   s_87_8,   s_86_8, 
  s_85_8,   s_84_8,   s_83_8,   s_82_8,   s_81_8,   s_80_8, 
  s_79_8,   s_78_8,   s_77_8,   s_76_8,   s_75_8,   s_74_8, 
  s_73_8,   s_72_8,   s_71_8,   s_70_8,   s_69_8,   s_68_8, 
  s_67_8,   s_66_8,   s_65_8,   s_64_8,   s_63_8,   s_62_8, 
  s_61_8,   s_60_8,   s_59_8,   s_58_8,   s_57_8,   s_56_8, 
  s_55_8,   s_54_8,   s_53_8,   s_52_8,   s_51_8,   s_50_8, 
  s_49_8,   s_48_8,   s_47_8,   s_46_8,   s_45_8,   s_44_8, 
  s_43_8,   s_42_8,   s_41_8,   s_40_8,   s_39_8,   s_38_8, 
  s_37_8,   s_36_8,   s_35_8,   s_34_8,   s_33_8,   s_32_8, 
  s_31_8,   s_30_8,   s_29_8,   s_28_8,   s_27_8,   s_26_8, 
  s_25_8,   s_24_8,   s_23_8,   s_22_8,   s_21_8,   s_20_8, 
  s_19_8,   s_18_8,   s_17_8,   s_16_8
} = partial_products[(width+2)*(8+1)-1:(width+2)*8];

assign {
 s_147_0,  s_146_0,  s_145_1,  s_144_1,  s_143_2,  s_142_2, 
 s_141_3,  s_140_3,  s_139_4,  s_138_4,  s_137_5,  s_136_5, 
 s_135_6,  s_134_6,  s_133_7,  s_132_7,  s_131_8,  s_130_8, 
 s_129_9,  s_128_9,  s_127_9,  s_126_9,  s_125_9,  s_124_9, 
 s_123_9,  s_122_9,  s_121_9,  s_120_9,  s_119_9,  s_118_9, 
 s_117_9,  s_116_9,  s_115_9,  s_114_9,  s_113_9,  s_112_9, 
 s_111_9,  s_110_9,  s_109_9,  s_108_9,  s_107_9,  s_106_9, 
 s_105_9,  s_104_9,  s_103_9,  s_102_9,  s_101_9,  s_100_9, 
  s_99_9,   s_98_9,   s_97_9,   s_96_9,   s_95_9,   s_94_9, 
  s_93_9,   s_92_9,   s_91_9,   s_90_9,   s_89_9,   s_88_9, 
  s_87_9,   s_86_9,   s_85_9,   s_84_9,   s_83_9,   s_82_9, 
  s_81_9,   s_80_9,   s_79_9,   s_78_9,   s_77_9,   s_76_9, 
  s_75_9,   s_74_9,   s_73_9,   s_72_9,   s_71_9,   s_70_9, 
  s_69_9,   s_68_9,   s_67_9,   s_66_9,   s_65_9,   s_64_9, 
  s_63_9,   s_62_9,   s_61_9,   s_60_9,   s_59_9,   s_58_9, 
  s_57_9,   s_56_9,   s_55_9,   s_54_9,   s_53_9,   s_52_9, 
  s_51_9,   s_50_9,   s_49_9,   s_48_9,   s_47_9,   s_46_9, 
  s_45_9,   s_44_9,   s_43_9,   s_42_9,   s_41_9,   s_40_9, 
  s_39_9,   s_38_9,   s_37_9,   s_36_9,   s_35_9,   s_34_9, 
  s_33_9,   s_32_9,   s_31_9,   s_30_9,   s_29_9,   s_28_9, 
  s_27_9,   s_26_9,   s_25_9,   s_24_9,   s_23_9,   s_22_9, 
  s_21_9,   s_20_9,   s_19_9,   s_18_9
} = partial_products[(width+2)*(9+1)-1:(width+2)*9];

assign {
 s_149_0,  s_148_0,  s_147_1,  s_146_1,  s_145_2,  s_144_2, 
 s_143_3,  s_142_3,  s_141_4,  s_140_4,  s_139_5,  s_138_5, 
 s_137_6,  s_136_6,  s_135_7,  s_134_7,  s_133_8,  s_132_8, 
 s_131_9,  s_130_9, s_129_10, s_128_10, s_127_10, s_126_10, 
s_125_10, s_124_10, s_123_10, s_122_10, s_121_10, s_120_10, 
s_119_10, s_118_10, s_117_10, s_116_10, s_115_10, s_114_10, 
s_113_10, s_112_10, s_111_10, s_110_10, s_109_10, s_108_10, 
s_107_10, s_106_10, s_105_10, s_104_10, s_103_10, s_102_10, 
s_101_10, s_100_10,  s_99_10,  s_98_10,  s_97_10,  s_96_10, 
 s_95_10,  s_94_10,  s_93_10,  s_92_10,  s_91_10,  s_90_10, 
 s_89_10,  s_88_10,  s_87_10,  s_86_10,  s_85_10,  s_84_10, 
 s_83_10,  s_82_10,  s_81_10,  s_80_10,  s_79_10,  s_78_10, 
 s_77_10,  s_76_10,  s_75_10,  s_74_10,  s_73_10,  s_72_10, 
 s_71_10,  s_70_10,  s_69_10,  s_68_10,  s_67_10,  s_66_10, 
 s_65_10,  s_64_10,  s_63_10,  s_62_10,  s_61_10,  s_60_10, 
 s_59_10,  s_58_10,  s_57_10,  s_56_10,  s_55_10,  s_54_10, 
 s_53_10,  s_52_10,  s_51_10,  s_50_10,  s_49_10,  s_48_10, 
 s_47_10,  s_46_10,  s_45_10,  s_44_10,  s_43_10,  s_42_10, 
 s_41_10,  s_40_10,  s_39_10,  s_38_10,  s_37_10,  s_36_10, 
 s_35_10,  s_34_10,  s_33_10,  s_32_10,  s_31_10,  s_30_10, 
 s_29_10,  s_28_10,  s_27_10,  s_26_10,  s_25_10,  s_24_10, 
 s_23_10,  s_22_10,  s_21_10,  s_20_10
} = partial_products[(width+2)*(10+1)-1:(width+2)*10];

assign {
 s_151_0,  s_150_0,  s_149_1,  s_148_1,  s_147_2,  s_146_2, 
 s_145_3,  s_144_3,  s_143_4,  s_142_4,  s_141_5,  s_140_5, 
 s_139_6,  s_138_6,  s_137_7,  s_136_7,  s_135_8,  s_134_8, 
 s_133_9,  s_132_9, s_131_10, s_130_10, s_129_11, s_128_11, 
s_127_11, s_126_11, s_125_11, s_124_11, s_123_11, s_122_11, 
s_121_11, s_120_11, s_119_11, s_118_11, s_117_11, s_116_11, 
s_115_11, s_114_11, s_113_11, s_112_11, s_111_11, s_110_11, 
s_109_11, s_108_11, s_107_11, s_106_11, s_105_11, s_104_11, 
s_103_11, s_102_11, s_101_11, s_100_11,  s_99_11,  s_98_11, 
 s_97_11,  s_96_11,  s_95_11,  s_94_11,  s_93_11,  s_92_11, 
 s_91_11,  s_90_11,  s_89_11,  s_88_11,  s_87_11,  s_86_11, 
 s_85_11,  s_84_11,  s_83_11,  s_82_11,  s_81_11,  s_80_11, 
 s_79_11,  s_78_11,  s_77_11,  s_76_11,  s_75_11,  s_74_11, 
 s_73_11,  s_72_11,  s_71_11,  s_70_11,  s_69_11,  s_68_11, 
 s_67_11,  s_66_11,  s_65_11,  s_64_11,  s_63_11,  s_62_11, 
 s_61_11,  s_60_11,  s_59_11,  s_58_11,  s_57_11,  s_56_11, 
 s_55_11,  s_54_11,  s_53_11,  s_52_11,  s_51_11,  s_50_11, 
 s_49_11,  s_48_11,  s_47_11,  s_46_11,  s_45_11,  s_44_11, 
 s_43_11,  s_42_11,  s_41_11,  s_40_11,  s_39_11,  s_38_11, 
 s_37_11,  s_36_11,  s_35_11,  s_34_11,  s_33_11,  s_32_11, 
 s_31_11,  s_30_11,  s_29_11,  s_28_11,  s_27_11,  s_26_11, 
 s_25_11,  s_24_11,  s_23_11,  s_22_11
} = partial_products[(width+2)*(11+1)-1:(width+2)*11];

assign {
 s_153_0,  s_152_0,  s_151_1,  s_150_1,  s_149_2,  s_148_2, 
 s_147_3,  s_146_3,  s_145_4,  s_144_4,  s_143_5,  s_142_5, 
 s_141_6,  s_140_6,  s_139_7,  s_138_7,  s_137_8,  s_136_8, 
 s_135_9,  s_134_9, s_133_10, s_132_10, s_131_11, s_130_11, 
s_129_12, s_128_12, s_127_12, s_126_12, s_125_12, s_124_12, 
s_123_12, s_122_12, s_121_12, s_120_12, s_119_12, s_118_12, 
s_117_12, s_116_12, s_115_12, s_114_12, s_113_12, s_112_12, 
s_111_12, s_110_12, s_109_12, s_108_12, s_107_12, s_106_12, 
s_105_12, s_104_12, s_103_12, s_102_12, s_101_12, s_100_12, 
 s_99_12,  s_98_12,  s_97_12,  s_96_12,  s_95_12,  s_94_12, 
 s_93_12,  s_92_12,  s_91_12,  s_90_12,  s_89_12,  s_88_12, 
 s_87_12,  s_86_12,  s_85_12,  s_84_12,  s_83_12,  s_82_12, 
 s_81_12,  s_80_12,  s_79_12,  s_78_12,  s_77_12,  s_76_12, 
 s_75_12,  s_74_12,  s_73_12,  s_72_12,  s_71_12,  s_70_12, 
 s_69_12,  s_68_12,  s_67_12,  s_66_12,  s_65_12,  s_64_12, 
 s_63_12,  s_62_12,  s_61_12,  s_60_12,  s_59_12,  s_58_12, 
 s_57_12,  s_56_12,  s_55_12,  s_54_12,  s_53_12,  s_52_12, 
 s_51_12,  s_50_12,  s_49_12,  s_48_12,  s_47_12,  s_46_12, 
 s_45_12,  s_44_12,  s_43_12,  s_42_12,  s_41_12,  s_40_12, 
 s_39_12,  s_38_12,  s_37_12,  s_36_12,  s_35_12,  s_34_12, 
 s_33_12,  s_32_12,  s_31_12,  s_30_12,  s_29_12,  s_28_12, 
 s_27_12,  s_26_12,  s_25_12,  s_24_12
} = partial_products[(width+2)*(12+1)-1:(width+2)*12];

assign {
 s_155_0,  s_154_0,  s_153_1,  s_152_1,  s_151_2,  s_150_2, 
 s_149_3,  s_148_3,  s_147_4,  s_146_4,  s_145_5,  s_144_5, 
 s_143_6,  s_142_6,  s_141_7,  s_140_7,  s_139_8,  s_138_8, 
 s_137_9,  s_136_9, s_135_10, s_134_10, s_133_11, s_132_11, 
s_131_12, s_130_12, s_129_13, s_128_13, s_127_13, s_126_13, 
s_125_13, s_124_13, s_123_13, s_122_13, s_121_13, s_120_13, 
s_119_13, s_118_13, s_117_13, s_116_13, s_115_13, s_114_13, 
s_113_13, s_112_13, s_111_13, s_110_13, s_109_13, s_108_13, 
s_107_13, s_106_13, s_105_13, s_104_13, s_103_13, s_102_13, 
s_101_13, s_100_13,  s_99_13,  s_98_13,  s_97_13,  s_96_13, 
 s_95_13,  s_94_13,  s_93_13,  s_92_13,  s_91_13,  s_90_13, 
 s_89_13,  s_88_13,  s_87_13,  s_86_13,  s_85_13,  s_84_13, 
 s_83_13,  s_82_13,  s_81_13,  s_80_13,  s_79_13,  s_78_13, 
 s_77_13,  s_76_13,  s_75_13,  s_74_13,  s_73_13,  s_72_13, 
 s_71_13,  s_70_13,  s_69_13,  s_68_13,  s_67_13,  s_66_13, 
 s_65_13,  s_64_13,  s_63_13,  s_62_13,  s_61_13,  s_60_13, 
 s_59_13,  s_58_13,  s_57_13,  s_56_13,  s_55_13,  s_54_13, 
 s_53_13,  s_52_13,  s_51_13,  s_50_13,  s_49_13,  s_48_13, 
 s_47_13,  s_46_13,  s_45_13,  s_44_13,  s_43_13,  s_42_13, 
 s_41_13,  s_40_13,  s_39_13,  s_38_13,  s_37_13,  s_36_13, 
 s_35_13,  s_34_13,  s_33_13,  s_32_13,  s_31_13,  s_30_13, 
 s_29_13,  s_28_13,  s_27_13,  s_26_13
} = partial_products[(width+2)*(13+1)-1:(width+2)*13];

assign {
 s_157_0,  s_156_0,  s_155_1,  s_154_1,  s_153_2,  s_152_2, 
 s_151_3,  s_150_3,  s_149_4,  s_148_4,  s_147_5,  s_146_5, 
 s_145_6,  s_144_6,  s_143_7,  s_142_7,  s_141_8,  s_140_8, 
 s_139_9,  s_138_9, s_137_10, s_136_10, s_135_11, s_134_11, 
s_133_12, s_132_12, s_131_13, s_130_13, s_129_14, s_128_14, 
s_127_14, s_126_14, s_125_14, s_124_14, s_123_14, s_122_14, 
s_121_14, s_120_14, s_119_14, s_118_14, s_117_14, s_116_14, 
s_115_14, s_114_14, s_113_14, s_112_14, s_111_14, s_110_14, 
s_109_14, s_108_14, s_107_14, s_106_14, s_105_14, s_104_14, 
s_103_14, s_102_14, s_101_14, s_100_14,  s_99_14,  s_98_14, 
 s_97_14,  s_96_14,  s_95_14,  s_94_14,  s_93_14,  s_92_14, 
 s_91_14,  s_90_14,  s_89_14,  s_88_14,  s_87_14,  s_86_14, 
 s_85_14,  s_84_14,  s_83_14,  s_82_14,  s_81_14,  s_80_14, 
 s_79_14,  s_78_14,  s_77_14,  s_76_14,  s_75_14,  s_74_14, 
 s_73_14,  s_72_14,  s_71_14,  s_70_14,  s_69_14,  s_68_14, 
 s_67_14,  s_66_14,  s_65_14,  s_64_14,  s_63_14,  s_62_14, 
 s_61_14,  s_60_14,  s_59_14,  s_58_14,  s_57_14,  s_56_14, 
 s_55_14,  s_54_14,  s_53_14,  s_52_14,  s_51_14,  s_50_14, 
 s_49_14,  s_48_14,  s_47_14,  s_46_14,  s_45_14,  s_44_14, 
 s_43_14,  s_42_14,  s_41_14,  s_40_14,  s_39_14,  s_38_14, 
 s_37_14,  s_36_14,  s_35_14,  s_34_14,  s_33_14,  s_32_14, 
 s_31_14,  s_30_14,  s_29_14,  s_28_14
} = partial_products[(width+2)*(14+1)-1:(width+2)*14];

assign {
 s_159_0,  s_158_0,  s_157_1,  s_156_1,  s_155_2,  s_154_2, 
 s_153_3,  s_152_3,  s_151_4,  s_150_4,  s_149_5,  s_148_5, 
 s_147_6,  s_146_6,  s_145_7,  s_144_7,  s_143_8,  s_142_8, 
 s_141_9,  s_140_9, s_139_10, s_138_10, s_137_11, s_136_11, 
s_135_12, s_134_12, s_133_13, s_132_13, s_131_14, s_130_14, 
s_129_15, s_128_15, s_127_15, s_126_15, s_125_15, s_124_15, 
s_123_15, s_122_15, s_121_15, s_120_15, s_119_15, s_118_15, 
s_117_15, s_116_15, s_115_15, s_114_15, s_113_15, s_112_15, 
s_111_15, s_110_15, s_109_15, s_108_15, s_107_15, s_106_15, 
s_105_15, s_104_15, s_103_15, s_102_15, s_101_15, s_100_15, 
 s_99_15,  s_98_15,  s_97_15,  s_96_15,  s_95_15,  s_94_15, 
 s_93_15,  s_92_15,  s_91_15,  s_90_15,  s_89_15,  s_88_15, 
 s_87_15,  s_86_15,  s_85_15,  s_84_15,  s_83_15,  s_82_15, 
 s_81_15,  s_80_15,  s_79_15,  s_78_15,  s_77_15,  s_76_15, 
 s_75_15,  s_74_15,  s_73_15,  s_72_15,  s_71_15,  s_70_15, 
 s_69_15,  s_68_15,  s_67_15,  s_66_15,  s_65_15,  s_64_15, 
 s_63_15,  s_62_15,  s_61_15,  s_60_15,  s_59_15,  s_58_15, 
 s_57_15,  s_56_15,  s_55_15,  s_54_15,  s_53_15,  s_52_15, 
 s_51_15,  s_50_15,  s_49_15,  s_48_15,  s_47_15,  s_46_15, 
 s_45_15,  s_44_15,  s_43_15,  s_42_15,  s_41_15,  s_40_15, 
 s_39_15,  s_38_15,  s_37_15,  s_36_15,  s_35_15,  s_34_15, 
 s_33_15,  s_32_15,  s_31_15,  s_30_15
} = partial_products[(width+2)*(15+1)-1:(width+2)*15];

assign {
 s_161_0,  s_160_0,  s_159_1,  s_158_1,  s_157_2,  s_156_2, 
 s_155_3,  s_154_3,  s_153_4,  s_152_4,  s_151_5,  s_150_5, 
 s_149_6,  s_148_6,  s_147_7,  s_146_7,  s_145_8,  s_144_8, 
 s_143_9,  s_142_9, s_141_10, s_140_10, s_139_11, s_138_11, 
s_137_12, s_136_12, s_135_13, s_134_13, s_133_14, s_132_14, 
s_131_15, s_130_15, s_129_16, s_128_16, s_127_16, s_126_16, 
s_125_16, s_124_16, s_123_16, s_122_16, s_121_16, s_120_16, 
s_119_16, s_118_16, s_117_16, s_116_16, s_115_16, s_114_16, 
s_113_16, s_112_16, s_111_16, s_110_16, s_109_16, s_108_16, 
s_107_16, s_106_16, s_105_16, s_104_16, s_103_16, s_102_16, 
s_101_16, s_100_16,  s_99_16,  s_98_16,  s_97_16,  s_96_16, 
 s_95_16,  s_94_16,  s_93_16,  s_92_16,  s_91_16,  s_90_16, 
 s_89_16,  s_88_16,  s_87_16,  s_86_16,  s_85_16,  s_84_16, 
 s_83_16,  s_82_16,  s_81_16,  s_80_16,  s_79_16,  s_78_16, 
 s_77_16,  s_76_16,  s_75_16,  s_74_16,  s_73_16,  s_72_16, 
 s_71_16,  s_70_16,  s_69_16,  s_68_16,  s_67_16,  s_66_16, 
 s_65_16,  s_64_16,  s_63_16,  s_62_16,  s_61_16,  s_60_16, 
 s_59_16,  s_58_16,  s_57_16,  s_56_16,  s_55_16,  s_54_16, 
 s_53_16,  s_52_16,  s_51_16,  s_50_16,  s_49_16,  s_48_16, 
 s_47_16,  s_46_16,  s_45_16,  s_44_16,  s_43_16,  s_42_16, 
 s_41_16,  s_40_16,  s_39_16,  s_38_16,  s_37_16,  s_36_16, 
 s_35_16,  s_34_16,  s_33_16,  s_32_16
} = partial_products[(width+2)*(16+1)-1:(width+2)*16];

assign {
 s_163_0,  s_162_0,  s_161_1,  s_160_1,  s_159_2,  s_158_2, 
 s_157_3,  s_156_3,  s_155_4,  s_154_4,  s_153_5,  s_152_5, 
 s_151_6,  s_150_6,  s_149_7,  s_148_7,  s_147_8,  s_146_8, 
 s_145_9,  s_144_9, s_143_10, s_142_10, s_141_11, s_140_11, 
s_139_12, s_138_12, s_137_13, s_136_13, s_135_14, s_134_14, 
s_133_15, s_132_15, s_131_16, s_130_16, s_129_17, s_128_17, 
s_127_17, s_126_17, s_125_17, s_124_17, s_123_17, s_122_17, 
s_121_17, s_120_17, s_119_17, s_118_17, s_117_17, s_116_17, 
s_115_17, s_114_17, s_113_17, s_112_17, s_111_17, s_110_17, 
s_109_17, s_108_17, s_107_17, s_106_17, s_105_17, s_104_17, 
s_103_17, s_102_17, s_101_17, s_100_17,  s_99_17,  s_98_17, 
 s_97_17,  s_96_17,  s_95_17,  s_94_17,  s_93_17,  s_92_17, 
 s_91_17,  s_90_17,  s_89_17,  s_88_17,  s_87_17,  s_86_17, 
 s_85_17,  s_84_17,  s_83_17,  s_82_17,  s_81_17,  s_80_17, 
 s_79_17,  s_78_17,  s_77_17,  s_76_17,  s_75_17,  s_74_17, 
 s_73_17,  s_72_17,  s_71_17,  s_70_17,  s_69_17,  s_68_17, 
 s_67_17,  s_66_17,  s_65_17,  s_64_17,  s_63_17,  s_62_17, 
 s_61_17,  s_60_17,  s_59_17,  s_58_17,  s_57_17,  s_56_17, 
 s_55_17,  s_54_17,  s_53_17,  s_52_17,  s_51_17,  s_50_17, 
 s_49_17,  s_48_17,  s_47_17,  s_46_17,  s_45_17,  s_44_17, 
 s_43_17,  s_42_17,  s_41_17,  s_40_17,  s_39_17,  s_38_17, 
 s_37_17,  s_36_17,  s_35_17,  s_34_17
} = partial_products[(width+2)*(17+1)-1:(width+2)*17];

assign {
 s_165_0,  s_164_0,  s_163_1,  s_162_1,  s_161_2,  s_160_2, 
 s_159_3,  s_158_3,  s_157_4,  s_156_4,  s_155_5,  s_154_5, 
 s_153_6,  s_152_6,  s_151_7,  s_150_7,  s_149_8,  s_148_8, 
 s_147_9,  s_146_9, s_145_10, s_144_10, s_143_11, s_142_11, 
s_141_12, s_140_12, s_139_13, s_138_13, s_137_14, s_136_14, 
s_135_15, s_134_15, s_133_16, s_132_16, s_131_17, s_130_17, 
s_129_18, s_128_18, s_127_18, s_126_18, s_125_18, s_124_18, 
s_123_18, s_122_18, s_121_18, s_120_18, s_119_18, s_118_18, 
s_117_18, s_116_18, s_115_18, s_114_18, s_113_18, s_112_18, 
s_111_18, s_110_18, s_109_18, s_108_18, s_107_18, s_106_18, 
s_105_18, s_104_18, s_103_18, s_102_18, s_101_18, s_100_18, 
 s_99_18,  s_98_18,  s_97_18,  s_96_18,  s_95_18,  s_94_18, 
 s_93_18,  s_92_18,  s_91_18,  s_90_18,  s_89_18,  s_88_18, 
 s_87_18,  s_86_18,  s_85_18,  s_84_18,  s_83_18,  s_82_18, 
 s_81_18,  s_80_18,  s_79_18,  s_78_18,  s_77_18,  s_76_18, 
 s_75_18,  s_74_18,  s_73_18,  s_72_18,  s_71_18,  s_70_18, 
 s_69_18,  s_68_18,  s_67_18,  s_66_18,  s_65_18,  s_64_18, 
 s_63_18,  s_62_18,  s_61_18,  s_60_18,  s_59_18,  s_58_18, 
 s_57_18,  s_56_18,  s_55_18,  s_54_18,  s_53_18,  s_52_18, 
 s_51_18,  s_50_18,  s_49_18,  s_48_18,  s_47_18,  s_46_18, 
 s_45_18,  s_44_18,  s_43_18,  s_42_18,  s_41_18,  s_40_18, 
 s_39_18,  s_38_18,  s_37_18,  s_36_18
} = partial_products[(width+2)*(18+1)-1:(width+2)*18];

assign {
 s_167_0,  s_166_0,  s_165_1,  s_164_1,  s_163_2,  s_162_2, 
 s_161_3,  s_160_3,  s_159_4,  s_158_4,  s_157_5,  s_156_5, 
 s_155_6,  s_154_6,  s_153_7,  s_152_7,  s_151_8,  s_150_8, 
 s_149_9,  s_148_9, s_147_10, s_146_10, s_145_11, s_144_11, 
s_143_12, s_142_12, s_141_13, s_140_13, s_139_14, s_138_14, 
s_137_15, s_136_15, s_135_16, s_134_16, s_133_17, s_132_17, 
s_131_18, s_130_18, s_129_19, s_128_19, s_127_19, s_126_19, 
s_125_19, s_124_19, s_123_19, s_122_19, s_121_19, s_120_19, 
s_119_19, s_118_19, s_117_19, s_116_19, s_115_19, s_114_19, 
s_113_19, s_112_19, s_111_19, s_110_19, s_109_19, s_108_19, 
s_107_19, s_106_19, s_105_19, s_104_19, s_103_19, s_102_19, 
s_101_19, s_100_19,  s_99_19,  s_98_19,  s_97_19,  s_96_19, 
 s_95_19,  s_94_19,  s_93_19,  s_92_19,  s_91_19,  s_90_19, 
 s_89_19,  s_88_19,  s_87_19,  s_86_19,  s_85_19,  s_84_19, 
 s_83_19,  s_82_19,  s_81_19,  s_80_19,  s_79_19,  s_78_19, 
 s_77_19,  s_76_19,  s_75_19,  s_74_19,  s_73_19,  s_72_19, 
 s_71_19,  s_70_19,  s_69_19,  s_68_19,  s_67_19,  s_66_19, 
 s_65_19,  s_64_19,  s_63_19,  s_62_19,  s_61_19,  s_60_19, 
 s_59_19,  s_58_19,  s_57_19,  s_56_19,  s_55_19,  s_54_19, 
 s_53_19,  s_52_19,  s_51_19,  s_50_19,  s_49_19,  s_48_19, 
 s_47_19,  s_46_19,  s_45_19,  s_44_19,  s_43_19,  s_42_19, 
 s_41_19,  s_40_19,  s_39_19,  s_38_19
} = partial_products[(width+2)*(19+1)-1:(width+2)*19];

assign {
 s_169_0,  s_168_0,  s_167_1,  s_166_1,  s_165_2,  s_164_2, 
 s_163_3,  s_162_3,  s_161_4,  s_160_4,  s_159_5,  s_158_5, 
 s_157_6,  s_156_6,  s_155_7,  s_154_7,  s_153_8,  s_152_8, 
 s_151_9,  s_150_9, s_149_10, s_148_10, s_147_11, s_146_11, 
s_145_12, s_144_12, s_143_13, s_142_13, s_141_14, s_140_14, 
s_139_15, s_138_15, s_137_16, s_136_16, s_135_17, s_134_17, 
s_133_18, s_132_18, s_131_19, s_130_19, s_129_20, s_128_20, 
s_127_20, s_126_20, s_125_20, s_124_20, s_123_20, s_122_20, 
s_121_20, s_120_20, s_119_20, s_118_20, s_117_20, s_116_20, 
s_115_20, s_114_20, s_113_20, s_112_20, s_111_20, s_110_20, 
s_109_20, s_108_20, s_107_20, s_106_20, s_105_20, s_104_20, 
s_103_20, s_102_20, s_101_20, s_100_20,  s_99_20,  s_98_20, 
 s_97_20,  s_96_20,  s_95_20,  s_94_20,  s_93_20,  s_92_20, 
 s_91_20,  s_90_20,  s_89_20,  s_88_20,  s_87_20,  s_86_20, 
 s_85_20,  s_84_20,  s_83_20,  s_82_20,  s_81_20,  s_80_20, 
 s_79_20,  s_78_20,  s_77_20,  s_76_20,  s_75_20,  s_74_20, 
 s_73_20,  s_72_20,  s_71_20,  s_70_20,  s_69_20,  s_68_20, 
 s_67_20,  s_66_20,  s_65_20,  s_64_20,  s_63_20,  s_62_20, 
 s_61_20,  s_60_20,  s_59_20,  s_58_20,  s_57_20,  s_56_20, 
 s_55_20,  s_54_20,  s_53_20,  s_52_20,  s_51_20,  s_50_20, 
 s_49_20,  s_48_20,  s_47_20,  s_46_20,  s_45_20,  s_44_20, 
 s_43_20,  s_42_20,  s_41_20,  s_40_20
} = partial_products[(width+2)*(20+1)-1:(width+2)*20];

assign {
 s_171_0,  s_170_0,  s_169_1,  s_168_1,  s_167_2,  s_166_2, 
 s_165_3,  s_164_3,  s_163_4,  s_162_4,  s_161_5,  s_160_5, 
 s_159_6,  s_158_6,  s_157_7,  s_156_7,  s_155_8,  s_154_8, 
 s_153_9,  s_152_9, s_151_10, s_150_10, s_149_11, s_148_11, 
s_147_12, s_146_12, s_145_13, s_144_13, s_143_14, s_142_14, 
s_141_15, s_140_15, s_139_16, s_138_16, s_137_17, s_136_17, 
s_135_18, s_134_18, s_133_19, s_132_19, s_131_20, s_130_20, 
s_129_21, s_128_21, s_127_21, s_126_21, s_125_21, s_124_21, 
s_123_21, s_122_21, s_121_21, s_120_21, s_119_21, s_118_21, 
s_117_21, s_116_21, s_115_21, s_114_21, s_113_21, s_112_21, 
s_111_21, s_110_21, s_109_21, s_108_21, s_107_21, s_106_21, 
s_105_21, s_104_21, s_103_21, s_102_21, s_101_21, s_100_21, 
 s_99_21,  s_98_21,  s_97_21,  s_96_21,  s_95_21,  s_94_21, 
 s_93_21,  s_92_21,  s_91_21,  s_90_21,  s_89_21,  s_88_21, 
 s_87_21,  s_86_21,  s_85_21,  s_84_21,  s_83_21,  s_82_21, 
 s_81_21,  s_80_21,  s_79_21,  s_78_21,  s_77_21,  s_76_21, 
 s_75_21,  s_74_21,  s_73_21,  s_72_21,  s_71_21,  s_70_21, 
 s_69_21,  s_68_21,  s_67_21,  s_66_21,  s_65_21,  s_64_21, 
 s_63_21,  s_62_21,  s_61_21,  s_60_21,  s_59_21,  s_58_21, 
 s_57_21,  s_56_21,  s_55_21,  s_54_21,  s_53_21,  s_52_21, 
 s_51_21,  s_50_21,  s_49_21,  s_48_21,  s_47_21,  s_46_21, 
 s_45_21,  s_44_21,  s_43_21,  s_42_21
} = partial_products[(width+2)*(21+1)-1:(width+2)*21];

assign {
 s_173_0,  s_172_0,  s_171_1,  s_170_1,  s_169_2,  s_168_2, 
 s_167_3,  s_166_3,  s_165_4,  s_164_4,  s_163_5,  s_162_5, 
 s_161_6,  s_160_6,  s_159_7,  s_158_7,  s_157_8,  s_156_8, 
 s_155_9,  s_154_9, s_153_10, s_152_10, s_151_11, s_150_11, 
s_149_12, s_148_12, s_147_13, s_146_13, s_145_14, s_144_14, 
s_143_15, s_142_15, s_141_16, s_140_16, s_139_17, s_138_17, 
s_137_18, s_136_18, s_135_19, s_134_19, s_133_20, s_132_20, 
s_131_21, s_130_21, s_129_22, s_128_22, s_127_22, s_126_22, 
s_125_22, s_124_22, s_123_22, s_122_22, s_121_22, s_120_22, 
s_119_22, s_118_22, s_117_22, s_116_22, s_115_22, s_114_22, 
s_113_22, s_112_22, s_111_22, s_110_22, s_109_22, s_108_22, 
s_107_22, s_106_22, s_105_22, s_104_22, s_103_22, s_102_22, 
s_101_22, s_100_22,  s_99_22,  s_98_22,  s_97_22,  s_96_22, 
 s_95_22,  s_94_22,  s_93_22,  s_92_22,  s_91_22,  s_90_22, 
 s_89_22,  s_88_22,  s_87_22,  s_86_22,  s_85_22,  s_84_22, 
 s_83_22,  s_82_22,  s_81_22,  s_80_22,  s_79_22,  s_78_22, 
 s_77_22,  s_76_22,  s_75_22,  s_74_22,  s_73_22,  s_72_22, 
 s_71_22,  s_70_22,  s_69_22,  s_68_22,  s_67_22,  s_66_22, 
 s_65_22,  s_64_22,  s_63_22,  s_62_22,  s_61_22,  s_60_22, 
 s_59_22,  s_58_22,  s_57_22,  s_56_22,  s_55_22,  s_54_22, 
 s_53_22,  s_52_22,  s_51_22,  s_50_22,  s_49_22,  s_48_22, 
 s_47_22,  s_46_22,  s_45_22,  s_44_22
} = partial_products[(width+2)*(22+1)-1:(width+2)*22];

assign {
 s_175_0,  s_174_0,  s_173_1,  s_172_1,  s_171_2,  s_170_2, 
 s_169_3,  s_168_3,  s_167_4,  s_166_4,  s_165_5,  s_164_5, 
 s_163_6,  s_162_6,  s_161_7,  s_160_7,  s_159_8,  s_158_8, 
 s_157_9,  s_156_9, s_155_10, s_154_10, s_153_11, s_152_11, 
s_151_12, s_150_12, s_149_13, s_148_13, s_147_14, s_146_14, 
s_145_15, s_144_15, s_143_16, s_142_16, s_141_17, s_140_17, 
s_139_18, s_138_18, s_137_19, s_136_19, s_135_20, s_134_20, 
s_133_21, s_132_21, s_131_22, s_130_22, s_129_23, s_128_23, 
s_127_23, s_126_23, s_125_23, s_124_23, s_123_23, s_122_23, 
s_121_23, s_120_23, s_119_23, s_118_23, s_117_23, s_116_23, 
s_115_23, s_114_23, s_113_23, s_112_23, s_111_23, s_110_23, 
s_109_23, s_108_23, s_107_23, s_106_23, s_105_23, s_104_23, 
s_103_23, s_102_23, s_101_23, s_100_23,  s_99_23,  s_98_23, 
 s_97_23,  s_96_23,  s_95_23,  s_94_23,  s_93_23,  s_92_23, 
 s_91_23,  s_90_23,  s_89_23,  s_88_23,  s_87_23,  s_86_23, 
 s_85_23,  s_84_23,  s_83_23,  s_82_23,  s_81_23,  s_80_23, 
 s_79_23,  s_78_23,  s_77_23,  s_76_23,  s_75_23,  s_74_23, 
 s_73_23,  s_72_23,  s_71_23,  s_70_23,  s_69_23,  s_68_23, 
 s_67_23,  s_66_23,  s_65_23,  s_64_23,  s_63_23,  s_62_23, 
 s_61_23,  s_60_23,  s_59_23,  s_58_23,  s_57_23,  s_56_23, 
 s_55_23,  s_54_23,  s_53_23,  s_52_23,  s_51_23,  s_50_23, 
 s_49_23,  s_48_23,  s_47_23,  s_46_23
} = partial_products[(width+2)*(23+1)-1:(width+2)*23];

assign {
 s_177_0,  s_176_0,  s_175_1,  s_174_1,  s_173_2,  s_172_2, 
 s_171_3,  s_170_3,  s_169_4,  s_168_4,  s_167_5,  s_166_5, 
 s_165_6,  s_164_6,  s_163_7,  s_162_7,  s_161_8,  s_160_8, 
 s_159_9,  s_158_9, s_157_10, s_156_10, s_155_11, s_154_11, 
s_153_12, s_152_12, s_151_13, s_150_13, s_149_14, s_148_14, 
s_147_15, s_146_15, s_145_16, s_144_16, s_143_17, s_142_17, 
s_141_18, s_140_18, s_139_19, s_138_19, s_137_20, s_136_20, 
s_135_21, s_134_21, s_133_22, s_132_22, s_131_23, s_130_23, 
s_129_24, s_128_24, s_127_24, s_126_24, s_125_24, s_124_24, 
s_123_24, s_122_24, s_121_24, s_120_24, s_119_24, s_118_24, 
s_117_24, s_116_24, s_115_24, s_114_24, s_113_24, s_112_24, 
s_111_24, s_110_24, s_109_24, s_108_24, s_107_24, s_106_24, 
s_105_24, s_104_24, s_103_24, s_102_24, s_101_24, s_100_24, 
 s_99_24,  s_98_24,  s_97_24,  s_96_24,  s_95_24,  s_94_24, 
 s_93_24,  s_92_24,  s_91_24,  s_90_24,  s_89_24,  s_88_24, 
 s_87_24,  s_86_24,  s_85_24,  s_84_24,  s_83_24,  s_82_24, 
 s_81_24,  s_80_24,  s_79_24,  s_78_24,  s_77_24,  s_76_24, 
 s_75_24,  s_74_24,  s_73_24,  s_72_24,  s_71_24,  s_70_24, 
 s_69_24,  s_68_24,  s_67_24,  s_66_24,  s_65_24,  s_64_24, 
 s_63_24,  s_62_24,  s_61_24,  s_60_24,  s_59_24,  s_58_24, 
 s_57_24,  s_56_24,  s_55_24,  s_54_24,  s_53_24,  s_52_24, 
 s_51_24,  s_50_24,  s_49_24,  s_48_24
} = partial_products[(width+2)*(24+1)-1:(width+2)*24];

assign {
 s_179_0,  s_178_0,  s_177_1,  s_176_1,  s_175_2,  s_174_2, 
 s_173_3,  s_172_3,  s_171_4,  s_170_4,  s_169_5,  s_168_5, 
 s_167_6,  s_166_6,  s_165_7,  s_164_7,  s_163_8,  s_162_8, 
 s_161_9,  s_160_9, s_159_10, s_158_10, s_157_11, s_156_11, 
s_155_12, s_154_12, s_153_13, s_152_13, s_151_14, s_150_14, 
s_149_15, s_148_15, s_147_16, s_146_16, s_145_17, s_144_17, 
s_143_18, s_142_18, s_141_19, s_140_19, s_139_20, s_138_20, 
s_137_21, s_136_21, s_135_22, s_134_22, s_133_23, s_132_23, 
s_131_24, s_130_24, s_129_25, s_128_25, s_127_25, s_126_25, 
s_125_25, s_124_25, s_123_25, s_122_25, s_121_25, s_120_25, 
s_119_25, s_118_25, s_117_25, s_116_25, s_115_25, s_114_25, 
s_113_25, s_112_25, s_111_25, s_110_25, s_109_25, s_108_25, 
s_107_25, s_106_25, s_105_25, s_104_25, s_103_25, s_102_25, 
s_101_25, s_100_25,  s_99_25,  s_98_25,  s_97_25,  s_96_25, 
 s_95_25,  s_94_25,  s_93_25,  s_92_25,  s_91_25,  s_90_25, 
 s_89_25,  s_88_25,  s_87_25,  s_86_25,  s_85_25,  s_84_25, 
 s_83_25,  s_82_25,  s_81_25,  s_80_25,  s_79_25,  s_78_25, 
 s_77_25,  s_76_25,  s_75_25,  s_74_25,  s_73_25,  s_72_25, 
 s_71_25,  s_70_25,  s_69_25,  s_68_25,  s_67_25,  s_66_25, 
 s_65_25,  s_64_25,  s_63_25,  s_62_25,  s_61_25,  s_60_25, 
 s_59_25,  s_58_25,  s_57_25,  s_56_25,  s_55_25,  s_54_25, 
 s_53_25,  s_52_25,  s_51_25,  s_50_25
} = partial_products[(width+2)*(25+1)-1:(width+2)*25];

assign {
 s_181_0,  s_180_0,  s_179_1,  s_178_1,  s_177_2,  s_176_2, 
 s_175_3,  s_174_3,  s_173_4,  s_172_4,  s_171_5,  s_170_5, 
 s_169_6,  s_168_6,  s_167_7,  s_166_7,  s_165_8,  s_164_8, 
 s_163_9,  s_162_9, s_161_10, s_160_10, s_159_11, s_158_11, 
s_157_12, s_156_12, s_155_13, s_154_13, s_153_14, s_152_14, 
s_151_15, s_150_15, s_149_16, s_148_16, s_147_17, s_146_17, 
s_145_18, s_144_18, s_143_19, s_142_19, s_141_20, s_140_20, 
s_139_21, s_138_21, s_137_22, s_136_22, s_135_23, s_134_23, 
s_133_24, s_132_24, s_131_25, s_130_25, s_129_26, s_128_26, 
s_127_26, s_126_26, s_125_26, s_124_26, s_123_26, s_122_26, 
s_121_26, s_120_26, s_119_26, s_118_26, s_117_26, s_116_26, 
s_115_26, s_114_26, s_113_26, s_112_26, s_111_26, s_110_26, 
s_109_26, s_108_26, s_107_26, s_106_26, s_105_26, s_104_26, 
s_103_26, s_102_26, s_101_26, s_100_26,  s_99_26,  s_98_26, 
 s_97_26,  s_96_26,  s_95_26,  s_94_26,  s_93_26,  s_92_26, 
 s_91_26,  s_90_26,  s_89_26,  s_88_26,  s_87_26,  s_86_26, 
 s_85_26,  s_84_26,  s_83_26,  s_82_26,  s_81_26,  s_80_26, 
 s_79_26,  s_78_26,  s_77_26,  s_76_26,  s_75_26,  s_74_26, 
 s_73_26,  s_72_26,  s_71_26,  s_70_26,  s_69_26,  s_68_26, 
 s_67_26,  s_66_26,  s_65_26,  s_64_26,  s_63_26,  s_62_26, 
 s_61_26,  s_60_26,  s_59_26,  s_58_26,  s_57_26,  s_56_26, 
 s_55_26,  s_54_26,  s_53_26,  s_52_26
} = partial_products[(width+2)*(26+1)-1:(width+2)*26];

assign {
 s_183_0,  s_182_0,  s_181_1,  s_180_1,  s_179_2,  s_178_2, 
 s_177_3,  s_176_3,  s_175_4,  s_174_4,  s_173_5,  s_172_5, 
 s_171_6,  s_170_6,  s_169_7,  s_168_7,  s_167_8,  s_166_8, 
 s_165_9,  s_164_9, s_163_10, s_162_10, s_161_11, s_160_11, 
s_159_12, s_158_12, s_157_13, s_156_13, s_155_14, s_154_14, 
s_153_15, s_152_15, s_151_16, s_150_16, s_149_17, s_148_17, 
s_147_18, s_146_18, s_145_19, s_144_19, s_143_20, s_142_20, 
s_141_21, s_140_21, s_139_22, s_138_22, s_137_23, s_136_23, 
s_135_24, s_134_24, s_133_25, s_132_25, s_131_26, s_130_26, 
s_129_27, s_128_27, s_127_27, s_126_27, s_125_27, s_124_27, 
s_123_27, s_122_27, s_121_27, s_120_27, s_119_27, s_118_27, 
s_117_27, s_116_27, s_115_27, s_114_27, s_113_27, s_112_27, 
s_111_27, s_110_27, s_109_27, s_108_27, s_107_27, s_106_27, 
s_105_27, s_104_27, s_103_27, s_102_27, s_101_27, s_100_27, 
 s_99_27,  s_98_27,  s_97_27,  s_96_27,  s_95_27,  s_94_27, 
 s_93_27,  s_92_27,  s_91_27,  s_90_27,  s_89_27,  s_88_27, 
 s_87_27,  s_86_27,  s_85_27,  s_84_27,  s_83_27,  s_82_27, 
 s_81_27,  s_80_27,  s_79_27,  s_78_27,  s_77_27,  s_76_27, 
 s_75_27,  s_74_27,  s_73_27,  s_72_27,  s_71_27,  s_70_27, 
 s_69_27,  s_68_27,  s_67_27,  s_66_27,  s_65_27,  s_64_27, 
 s_63_27,  s_62_27,  s_61_27,  s_60_27,  s_59_27,  s_58_27, 
 s_57_27,  s_56_27,  s_55_27,  s_54_27
} = partial_products[(width+2)*(27+1)-1:(width+2)*27];

assign {
 s_185_0,  s_184_0,  s_183_1,  s_182_1,  s_181_2,  s_180_2, 
 s_179_3,  s_178_3,  s_177_4,  s_176_4,  s_175_5,  s_174_5, 
 s_173_6,  s_172_6,  s_171_7,  s_170_7,  s_169_8,  s_168_8, 
 s_167_9,  s_166_9, s_165_10, s_164_10, s_163_11, s_162_11, 
s_161_12, s_160_12, s_159_13, s_158_13, s_157_14, s_156_14, 
s_155_15, s_154_15, s_153_16, s_152_16, s_151_17, s_150_17, 
s_149_18, s_148_18, s_147_19, s_146_19, s_145_20, s_144_20, 
s_143_21, s_142_21, s_141_22, s_140_22, s_139_23, s_138_23, 
s_137_24, s_136_24, s_135_25, s_134_25, s_133_26, s_132_26, 
s_131_27, s_130_27, s_129_28, s_128_28, s_127_28, s_126_28, 
s_125_28, s_124_28, s_123_28, s_122_28, s_121_28, s_120_28, 
s_119_28, s_118_28, s_117_28, s_116_28, s_115_28, s_114_28, 
s_113_28, s_112_28, s_111_28, s_110_28, s_109_28, s_108_28, 
s_107_28, s_106_28, s_105_28, s_104_28, s_103_28, s_102_28, 
s_101_28, s_100_28,  s_99_28,  s_98_28,  s_97_28,  s_96_28, 
 s_95_28,  s_94_28,  s_93_28,  s_92_28,  s_91_28,  s_90_28, 
 s_89_28,  s_88_28,  s_87_28,  s_86_28,  s_85_28,  s_84_28, 
 s_83_28,  s_82_28,  s_81_28,  s_80_28,  s_79_28,  s_78_28, 
 s_77_28,  s_76_28,  s_75_28,  s_74_28,  s_73_28,  s_72_28, 
 s_71_28,  s_70_28,  s_69_28,  s_68_28,  s_67_28,  s_66_28, 
 s_65_28,  s_64_28,  s_63_28,  s_62_28,  s_61_28,  s_60_28, 
 s_59_28,  s_58_28,  s_57_28,  s_56_28
} = partial_products[(width+2)*(28+1)-1:(width+2)*28];

assign {
 s_187_0,  s_186_0,  s_185_1,  s_184_1,  s_183_2,  s_182_2, 
 s_181_3,  s_180_3,  s_179_4,  s_178_4,  s_177_5,  s_176_5, 
 s_175_6,  s_174_6,  s_173_7,  s_172_7,  s_171_8,  s_170_8, 
 s_169_9,  s_168_9, s_167_10, s_166_10, s_165_11, s_164_11, 
s_163_12, s_162_12, s_161_13, s_160_13, s_159_14, s_158_14, 
s_157_15, s_156_15, s_155_16, s_154_16, s_153_17, s_152_17, 
s_151_18, s_150_18, s_149_19, s_148_19, s_147_20, s_146_20, 
s_145_21, s_144_21, s_143_22, s_142_22, s_141_23, s_140_23, 
s_139_24, s_138_24, s_137_25, s_136_25, s_135_26, s_134_26, 
s_133_27, s_132_27, s_131_28, s_130_28, s_129_29, s_128_29, 
s_127_29, s_126_29, s_125_29, s_124_29, s_123_29, s_122_29, 
s_121_29, s_120_29, s_119_29, s_118_29, s_117_29, s_116_29, 
s_115_29, s_114_29, s_113_29, s_112_29, s_111_29, s_110_29, 
s_109_29, s_108_29, s_107_29, s_106_29, s_105_29, s_104_29, 
s_103_29, s_102_29, s_101_29, s_100_29,  s_99_29,  s_98_29, 
 s_97_29,  s_96_29,  s_95_29,  s_94_29,  s_93_29,  s_92_29, 
 s_91_29,  s_90_29,  s_89_29,  s_88_29,  s_87_29,  s_86_29, 
 s_85_29,  s_84_29,  s_83_29,  s_82_29,  s_81_29,  s_80_29, 
 s_79_29,  s_78_29,  s_77_29,  s_76_29,  s_75_29,  s_74_29, 
 s_73_29,  s_72_29,  s_71_29,  s_70_29,  s_69_29,  s_68_29, 
 s_67_29,  s_66_29,  s_65_29,  s_64_29,  s_63_29,  s_62_29, 
 s_61_29,  s_60_29,  s_59_29,  s_58_29
} = partial_products[(width+2)*(29+1)-1:(width+2)*29];

assign {
 s_189_0,  s_188_0,  s_187_1,  s_186_1,  s_185_2,  s_184_2, 
 s_183_3,  s_182_3,  s_181_4,  s_180_4,  s_179_5,  s_178_5, 
 s_177_6,  s_176_6,  s_175_7,  s_174_7,  s_173_8,  s_172_8, 
 s_171_9,  s_170_9, s_169_10, s_168_10, s_167_11, s_166_11, 
s_165_12, s_164_12, s_163_13, s_162_13, s_161_14, s_160_14, 
s_159_15, s_158_15, s_157_16, s_156_16, s_155_17, s_154_17, 
s_153_18, s_152_18, s_151_19, s_150_19, s_149_20, s_148_20, 
s_147_21, s_146_21, s_145_22, s_144_22, s_143_23, s_142_23, 
s_141_24, s_140_24, s_139_25, s_138_25, s_137_26, s_136_26, 
s_135_27, s_134_27, s_133_28, s_132_28, s_131_29, s_130_29, 
s_129_30, s_128_30, s_127_30, s_126_30, s_125_30, s_124_30, 
s_123_30, s_122_30, s_121_30, s_120_30, s_119_30, s_118_30, 
s_117_30, s_116_30, s_115_30, s_114_30, s_113_30, s_112_30, 
s_111_30, s_110_30, s_109_30, s_108_30, s_107_30, s_106_30, 
s_105_30, s_104_30, s_103_30, s_102_30, s_101_30, s_100_30, 
 s_99_30,  s_98_30,  s_97_30,  s_96_30,  s_95_30,  s_94_30, 
 s_93_30,  s_92_30,  s_91_30,  s_90_30,  s_89_30,  s_88_30, 
 s_87_30,  s_86_30,  s_85_30,  s_84_30,  s_83_30,  s_82_30, 
 s_81_30,  s_80_30,  s_79_30,  s_78_30,  s_77_30,  s_76_30, 
 s_75_30,  s_74_30,  s_73_30,  s_72_30,  s_71_30,  s_70_30, 
 s_69_30,  s_68_30,  s_67_30,  s_66_30,  s_65_30,  s_64_30, 
 s_63_30,  s_62_30,  s_61_30,  s_60_30
} = partial_products[(width+2)*(30+1)-1:(width+2)*30];

assign {
 s_191_0,  s_190_0,  s_189_1,  s_188_1,  s_187_2,  s_186_2, 
 s_185_3,  s_184_3,  s_183_4,  s_182_4,  s_181_5,  s_180_5, 
 s_179_6,  s_178_6,  s_177_7,  s_176_7,  s_175_8,  s_174_8, 
 s_173_9,  s_172_9, s_171_10, s_170_10, s_169_11, s_168_11, 
s_167_12, s_166_12, s_165_13, s_164_13, s_163_14, s_162_14, 
s_161_15, s_160_15, s_159_16, s_158_16, s_157_17, s_156_17, 
s_155_18, s_154_18, s_153_19, s_152_19, s_151_20, s_150_20, 
s_149_21, s_148_21, s_147_22, s_146_22, s_145_23, s_144_23, 
s_143_24, s_142_24, s_141_25, s_140_25, s_139_26, s_138_26, 
s_137_27, s_136_27, s_135_28, s_134_28, s_133_29, s_132_29, 
s_131_30, s_130_30, s_129_31, s_128_31, s_127_31, s_126_31, 
s_125_31, s_124_31, s_123_31, s_122_31, s_121_31, s_120_31, 
s_119_31, s_118_31, s_117_31, s_116_31, s_115_31, s_114_31, 
s_113_31, s_112_31, s_111_31, s_110_31, s_109_31, s_108_31, 
s_107_31, s_106_31, s_105_31, s_104_31, s_103_31, s_102_31, 
s_101_31, s_100_31,  s_99_31,  s_98_31,  s_97_31,  s_96_31, 
 s_95_31,  s_94_31,  s_93_31,  s_92_31,  s_91_31,  s_90_31, 
 s_89_31,  s_88_31,  s_87_31,  s_86_31,  s_85_31,  s_84_31, 
 s_83_31,  s_82_31,  s_81_31,  s_80_31,  s_79_31,  s_78_31, 
 s_77_31,  s_76_31,  s_75_31,  s_74_31,  s_73_31,  s_72_31, 
 s_71_31,  s_70_31,  s_69_31,  s_68_31,  s_67_31,  s_66_31, 
 s_65_31,  s_64_31,  s_63_31,  s_62_31
} = partial_products[(width+2)*(31+1)-1:(width+2)*31];

assign {
 s_193_0,  s_192_0,  s_191_1,  s_190_1,  s_189_2,  s_188_2, 
 s_187_3,  s_186_3,  s_185_4,  s_184_4,  s_183_5,  s_182_5, 
 s_181_6,  s_180_6,  s_179_7,  s_178_7,  s_177_8,  s_176_8, 
 s_175_9,  s_174_9, s_173_10, s_172_10, s_171_11, s_170_11, 
s_169_12, s_168_12, s_167_13, s_166_13, s_165_14, s_164_14, 
s_163_15, s_162_15, s_161_16, s_160_16, s_159_17, s_158_17, 
s_157_18, s_156_18, s_155_19, s_154_19, s_153_20, s_152_20, 
s_151_21, s_150_21, s_149_22, s_148_22, s_147_23, s_146_23, 
s_145_24, s_144_24, s_143_25, s_142_25, s_141_26, s_140_26, 
s_139_27, s_138_27, s_137_28, s_136_28, s_135_29, s_134_29, 
s_133_30, s_132_30, s_131_31, s_130_31, s_129_32, s_128_32, 
s_127_32, s_126_32, s_125_32, s_124_32, s_123_32, s_122_32, 
s_121_32, s_120_32, s_119_32, s_118_32, s_117_32, s_116_32, 
s_115_32, s_114_32, s_113_32, s_112_32, s_111_32, s_110_32, 
s_109_32, s_108_32, s_107_32, s_106_32, s_105_32, s_104_32, 
s_103_32, s_102_32, s_101_32, s_100_32,  s_99_32,  s_98_32, 
 s_97_32,  s_96_32,  s_95_32,  s_94_32,  s_93_32,  s_92_32, 
 s_91_32,  s_90_32,  s_89_32,  s_88_32,  s_87_32,  s_86_32, 
 s_85_32,  s_84_32,  s_83_32,  s_82_32,  s_81_32,  s_80_32, 
 s_79_32,  s_78_32,  s_77_32,  s_76_32,  s_75_32,  s_74_32, 
 s_73_32,  s_72_32,  s_71_32,  s_70_32,  s_69_32,  s_68_32, 
 s_67_32,  s_66_32,  s_65_32,  s_64_32
} = partial_products[(width+2)*(32+1)-1:(width+2)*32];

assign {
 s_195_0,  s_194_0,  s_193_1,  s_192_1,  s_191_2,  s_190_2, 
 s_189_3,  s_188_3,  s_187_4,  s_186_4,  s_185_5,  s_184_5, 
 s_183_6,  s_182_6,  s_181_7,  s_180_7,  s_179_8,  s_178_8, 
 s_177_9,  s_176_9, s_175_10, s_174_10, s_173_11, s_172_11, 
s_171_12, s_170_12, s_169_13, s_168_13, s_167_14, s_166_14, 
s_165_15, s_164_15, s_163_16, s_162_16, s_161_17, s_160_17, 
s_159_18, s_158_18, s_157_19, s_156_19, s_155_20, s_154_20, 
s_153_21, s_152_21, s_151_22, s_150_22, s_149_23, s_148_23, 
s_147_24, s_146_24, s_145_25, s_144_25, s_143_26, s_142_26, 
s_141_27, s_140_27, s_139_28, s_138_28, s_137_29, s_136_29, 
s_135_30, s_134_30, s_133_31, s_132_31, s_131_32, s_130_32, 
s_129_33, s_128_33, s_127_33, s_126_33, s_125_33, s_124_33, 
s_123_33, s_122_33, s_121_33, s_120_33, s_119_33, s_118_33, 
s_117_33, s_116_33, s_115_33, s_114_33, s_113_33, s_112_33, 
s_111_33, s_110_33, s_109_33, s_108_33, s_107_33, s_106_33, 
s_105_33, s_104_33, s_103_33, s_102_33, s_101_33, s_100_33, 
 s_99_33,  s_98_33,  s_97_33,  s_96_33,  s_95_33,  s_94_33, 
 s_93_33,  s_92_33,  s_91_33,  s_90_33,  s_89_33,  s_88_33, 
 s_87_33,  s_86_33,  s_85_33,  s_84_33,  s_83_33,  s_82_33, 
 s_81_33,  s_80_33,  s_79_33,  s_78_33,  s_77_33,  s_76_33, 
 s_75_33,  s_74_33,  s_73_33,  s_72_33,  s_71_33,  s_70_33, 
 s_69_33,  s_68_33,  s_67_33,  s_66_33
} = partial_products[(width+2)*(33+1)-1:(width+2)*33];

assign {
 s_197_0,  s_196_0,  s_195_1,  s_194_1,  s_193_2,  s_192_2, 
 s_191_3,  s_190_3,  s_189_4,  s_188_4,  s_187_5,  s_186_5, 
 s_185_6,  s_184_6,  s_183_7,  s_182_7,  s_181_8,  s_180_8, 
 s_179_9,  s_178_9, s_177_10, s_176_10, s_175_11, s_174_11, 
s_173_12, s_172_12, s_171_13, s_170_13, s_169_14, s_168_14, 
s_167_15, s_166_15, s_165_16, s_164_16, s_163_17, s_162_17, 
s_161_18, s_160_18, s_159_19, s_158_19, s_157_20, s_156_20, 
s_155_21, s_154_21, s_153_22, s_152_22, s_151_23, s_150_23, 
s_149_24, s_148_24, s_147_25, s_146_25, s_145_26, s_144_26, 
s_143_27, s_142_27, s_141_28, s_140_28, s_139_29, s_138_29, 
s_137_30, s_136_30, s_135_31, s_134_31, s_133_32, s_132_32, 
s_131_33, s_130_33, s_129_34, s_128_34, s_127_34, s_126_34, 
s_125_34, s_124_34, s_123_34, s_122_34, s_121_34, s_120_34, 
s_119_34, s_118_34, s_117_34, s_116_34, s_115_34, s_114_34, 
s_113_34, s_112_34, s_111_34, s_110_34, s_109_34, s_108_34, 
s_107_34, s_106_34, s_105_34, s_104_34, s_103_34, s_102_34, 
s_101_34, s_100_34,  s_99_34,  s_98_34,  s_97_34,  s_96_34, 
 s_95_34,  s_94_34,  s_93_34,  s_92_34,  s_91_34,  s_90_34, 
 s_89_34,  s_88_34,  s_87_34,  s_86_34,  s_85_34,  s_84_34, 
 s_83_34,  s_82_34,  s_81_34,  s_80_34,  s_79_34,  s_78_34, 
 s_77_34,  s_76_34,  s_75_34,  s_74_34,  s_73_34,  s_72_34, 
 s_71_34,  s_70_34,  s_69_34,  s_68_34
} = partial_products[(width+2)*(34+1)-1:(width+2)*34];

assign {
 s_199_0,  s_198_0,  s_197_1,  s_196_1,  s_195_2,  s_194_2, 
 s_193_3,  s_192_3,  s_191_4,  s_190_4,  s_189_5,  s_188_5, 
 s_187_6,  s_186_6,  s_185_7,  s_184_7,  s_183_8,  s_182_8, 
 s_181_9,  s_180_9, s_179_10, s_178_10, s_177_11, s_176_11, 
s_175_12, s_174_12, s_173_13, s_172_13, s_171_14, s_170_14, 
s_169_15, s_168_15, s_167_16, s_166_16, s_165_17, s_164_17, 
s_163_18, s_162_18, s_161_19, s_160_19, s_159_20, s_158_20, 
s_157_21, s_156_21, s_155_22, s_154_22, s_153_23, s_152_23, 
s_151_24, s_150_24, s_149_25, s_148_25, s_147_26, s_146_26, 
s_145_27, s_144_27, s_143_28, s_142_28, s_141_29, s_140_29, 
s_139_30, s_138_30, s_137_31, s_136_31, s_135_32, s_134_32, 
s_133_33, s_132_33, s_131_34, s_130_34, s_129_35, s_128_35, 
s_127_35, s_126_35, s_125_35, s_124_35, s_123_35, s_122_35, 
s_121_35, s_120_35, s_119_35, s_118_35, s_117_35, s_116_35, 
s_115_35, s_114_35, s_113_35, s_112_35, s_111_35, s_110_35, 
s_109_35, s_108_35, s_107_35, s_106_35, s_105_35, s_104_35, 
s_103_35, s_102_35, s_101_35, s_100_35,  s_99_35,  s_98_35, 
 s_97_35,  s_96_35,  s_95_35,  s_94_35,  s_93_35,  s_92_35, 
 s_91_35,  s_90_35,  s_89_35,  s_88_35,  s_87_35,  s_86_35, 
 s_85_35,  s_84_35,  s_83_35,  s_82_35,  s_81_35,  s_80_35, 
 s_79_35,  s_78_35,  s_77_35,  s_76_35,  s_75_35,  s_74_35, 
 s_73_35,  s_72_35,  s_71_35,  s_70_35
} = partial_products[(width+2)*(35+1)-1:(width+2)*35];

assign {
 s_201_0,  s_200_0,  s_199_1,  s_198_1,  s_197_2,  s_196_2, 
 s_195_3,  s_194_3,  s_193_4,  s_192_4,  s_191_5,  s_190_5, 
 s_189_6,  s_188_6,  s_187_7,  s_186_7,  s_185_8,  s_184_8, 
 s_183_9,  s_182_9, s_181_10, s_180_10, s_179_11, s_178_11, 
s_177_12, s_176_12, s_175_13, s_174_13, s_173_14, s_172_14, 
s_171_15, s_170_15, s_169_16, s_168_16, s_167_17, s_166_17, 
s_165_18, s_164_18, s_163_19, s_162_19, s_161_20, s_160_20, 
s_159_21, s_158_21, s_157_22, s_156_22, s_155_23, s_154_23, 
s_153_24, s_152_24, s_151_25, s_150_25, s_149_26, s_148_26, 
s_147_27, s_146_27, s_145_28, s_144_28, s_143_29, s_142_29, 
s_141_30, s_140_30, s_139_31, s_138_31, s_137_32, s_136_32, 
s_135_33, s_134_33, s_133_34, s_132_34, s_131_35, s_130_35, 
s_129_36, s_128_36, s_127_36, s_126_36, s_125_36, s_124_36, 
s_123_36, s_122_36, s_121_36, s_120_36, s_119_36, s_118_36, 
s_117_36, s_116_36, s_115_36, s_114_36, s_113_36, s_112_36, 
s_111_36, s_110_36, s_109_36, s_108_36, s_107_36, s_106_36, 
s_105_36, s_104_36, s_103_36, s_102_36, s_101_36, s_100_36, 
 s_99_36,  s_98_36,  s_97_36,  s_96_36,  s_95_36,  s_94_36, 
 s_93_36,  s_92_36,  s_91_36,  s_90_36,  s_89_36,  s_88_36, 
 s_87_36,  s_86_36,  s_85_36,  s_84_36,  s_83_36,  s_82_36, 
 s_81_36,  s_80_36,  s_79_36,  s_78_36,  s_77_36,  s_76_36, 
 s_75_36,  s_74_36,  s_73_36,  s_72_36
} = partial_products[(width+2)*(36+1)-1:(width+2)*36];

assign {
 s_203_0,  s_202_0,  s_201_1,  s_200_1,  s_199_2,  s_198_2, 
 s_197_3,  s_196_3,  s_195_4,  s_194_4,  s_193_5,  s_192_5, 
 s_191_6,  s_190_6,  s_189_7,  s_188_7,  s_187_8,  s_186_8, 
 s_185_9,  s_184_9, s_183_10, s_182_10, s_181_11, s_180_11, 
s_179_12, s_178_12, s_177_13, s_176_13, s_175_14, s_174_14, 
s_173_15, s_172_15, s_171_16, s_170_16, s_169_17, s_168_17, 
s_167_18, s_166_18, s_165_19, s_164_19, s_163_20, s_162_20, 
s_161_21, s_160_21, s_159_22, s_158_22, s_157_23, s_156_23, 
s_155_24, s_154_24, s_153_25, s_152_25, s_151_26, s_150_26, 
s_149_27, s_148_27, s_147_28, s_146_28, s_145_29, s_144_29, 
s_143_30, s_142_30, s_141_31, s_140_31, s_139_32, s_138_32, 
s_137_33, s_136_33, s_135_34, s_134_34, s_133_35, s_132_35, 
s_131_36, s_130_36, s_129_37, s_128_37, s_127_37, s_126_37, 
s_125_37, s_124_37, s_123_37, s_122_37, s_121_37, s_120_37, 
s_119_37, s_118_37, s_117_37, s_116_37, s_115_37, s_114_37, 
s_113_37, s_112_37, s_111_37, s_110_37, s_109_37, s_108_37, 
s_107_37, s_106_37, s_105_37, s_104_37, s_103_37, s_102_37, 
s_101_37, s_100_37,  s_99_37,  s_98_37,  s_97_37,  s_96_37, 
 s_95_37,  s_94_37,  s_93_37,  s_92_37,  s_91_37,  s_90_37, 
 s_89_37,  s_88_37,  s_87_37,  s_86_37,  s_85_37,  s_84_37, 
 s_83_37,  s_82_37,  s_81_37,  s_80_37,  s_79_37,  s_78_37, 
 s_77_37,  s_76_37,  s_75_37,  s_74_37
} = partial_products[(width+2)*(37+1)-1:(width+2)*37];

assign {
 s_205_0,  s_204_0,  s_203_1,  s_202_1,  s_201_2,  s_200_2, 
 s_199_3,  s_198_3,  s_197_4,  s_196_4,  s_195_5,  s_194_5, 
 s_193_6,  s_192_6,  s_191_7,  s_190_7,  s_189_8,  s_188_8, 
 s_187_9,  s_186_9, s_185_10, s_184_10, s_183_11, s_182_11, 
s_181_12, s_180_12, s_179_13, s_178_13, s_177_14, s_176_14, 
s_175_15, s_174_15, s_173_16, s_172_16, s_171_17, s_170_17, 
s_169_18, s_168_18, s_167_19, s_166_19, s_165_20, s_164_20, 
s_163_21, s_162_21, s_161_22, s_160_22, s_159_23, s_158_23, 
s_157_24, s_156_24, s_155_25, s_154_25, s_153_26, s_152_26, 
s_151_27, s_150_27, s_149_28, s_148_28, s_147_29, s_146_29, 
s_145_30, s_144_30, s_143_31, s_142_31, s_141_32, s_140_32, 
s_139_33, s_138_33, s_137_34, s_136_34, s_135_35, s_134_35, 
s_133_36, s_132_36, s_131_37, s_130_37, s_129_38, s_128_38, 
s_127_38, s_126_38, s_125_38, s_124_38, s_123_38, s_122_38, 
s_121_38, s_120_38, s_119_38, s_118_38, s_117_38, s_116_38, 
s_115_38, s_114_38, s_113_38, s_112_38, s_111_38, s_110_38, 
s_109_38, s_108_38, s_107_38, s_106_38, s_105_38, s_104_38, 
s_103_38, s_102_38, s_101_38, s_100_38,  s_99_38,  s_98_38, 
 s_97_38,  s_96_38,  s_95_38,  s_94_38,  s_93_38,  s_92_38, 
 s_91_38,  s_90_38,  s_89_38,  s_88_38,  s_87_38,  s_86_38, 
 s_85_38,  s_84_38,  s_83_38,  s_82_38,  s_81_38,  s_80_38, 
 s_79_38,  s_78_38,  s_77_38,  s_76_38
} = partial_products[(width+2)*(38+1)-1:(width+2)*38];

assign {
 s_207_0,  s_206_0,  s_205_1,  s_204_1,  s_203_2,  s_202_2, 
 s_201_3,  s_200_3,  s_199_4,  s_198_4,  s_197_5,  s_196_5, 
 s_195_6,  s_194_6,  s_193_7,  s_192_7,  s_191_8,  s_190_8, 
 s_189_9,  s_188_9, s_187_10, s_186_10, s_185_11, s_184_11, 
s_183_12, s_182_12, s_181_13, s_180_13, s_179_14, s_178_14, 
s_177_15, s_176_15, s_175_16, s_174_16, s_173_17, s_172_17, 
s_171_18, s_170_18, s_169_19, s_168_19, s_167_20, s_166_20, 
s_165_21, s_164_21, s_163_22, s_162_22, s_161_23, s_160_23, 
s_159_24, s_158_24, s_157_25, s_156_25, s_155_26, s_154_26, 
s_153_27, s_152_27, s_151_28, s_150_28, s_149_29, s_148_29, 
s_147_30, s_146_30, s_145_31, s_144_31, s_143_32, s_142_32, 
s_141_33, s_140_33, s_139_34, s_138_34, s_137_35, s_136_35, 
s_135_36, s_134_36, s_133_37, s_132_37, s_131_38, s_130_38, 
s_129_39, s_128_39, s_127_39, s_126_39, s_125_39, s_124_39, 
s_123_39, s_122_39, s_121_39, s_120_39, s_119_39, s_118_39, 
s_117_39, s_116_39, s_115_39, s_114_39, s_113_39, s_112_39, 
s_111_39, s_110_39, s_109_39, s_108_39, s_107_39, s_106_39, 
s_105_39, s_104_39, s_103_39, s_102_39, s_101_39, s_100_39, 
 s_99_39,  s_98_39,  s_97_39,  s_96_39,  s_95_39,  s_94_39, 
 s_93_39,  s_92_39,  s_91_39,  s_90_39,  s_89_39,  s_88_39, 
 s_87_39,  s_86_39,  s_85_39,  s_84_39,  s_83_39,  s_82_39, 
 s_81_39,  s_80_39,  s_79_39,  s_78_39
} = partial_products[(width+2)*(39+1)-1:(width+2)*39];

assign {
 s_209_0,  s_208_0,  s_207_1,  s_206_1,  s_205_2,  s_204_2, 
 s_203_3,  s_202_3,  s_201_4,  s_200_4,  s_199_5,  s_198_5, 
 s_197_6,  s_196_6,  s_195_7,  s_194_7,  s_193_8,  s_192_8, 
 s_191_9,  s_190_9, s_189_10, s_188_10, s_187_11, s_186_11, 
s_185_12, s_184_12, s_183_13, s_182_13, s_181_14, s_180_14, 
s_179_15, s_178_15, s_177_16, s_176_16, s_175_17, s_174_17, 
s_173_18, s_172_18, s_171_19, s_170_19, s_169_20, s_168_20, 
s_167_21, s_166_21, s_165_22, s_164_22, s_163_23, s_162_23, 
s_161_24, s_160_24, s_159_25, s_158_25, s_157_26, s_156_26, 
s_155_27, s_154_27, s_153_28, s_152_28, s_151_29, s_150_29, 
s_149_30, s_148_30, s_147_31, s_146_31, s_145_32, s_144_32, 
s_143_33, s_142_33, s_141_34, s_140_34, s_139_35, s_138_35, 
s_137_36, s_136_36, s_135_37, s_134_37, s_133_38, s_132_38, 
s_131_39, s_130_39, s_129_40, s_128_40, s_127_40, s_126_40, 
s_125_40, s_124_40, s_123_40, s_122_40, s_121_40, s_120_40, 
s_119_40, s_118_40, s_117_40, s_116_40, s_115_40, s_114_40, 
s_113_40, s_112_40, s_111_40, s_110_40, s_109_40, s_108_40, 
s_107_40, s_106_40, s_105_40, s_104_40, s_103_40, s_102_40, 
s_101_40, s_100_40,  s_99_40,  s_98_40,  s_97_40,  s_96_40, 
 s_95_40,  s_94_40,  s_93_40,  s_92_40,  s_91_40,  s_90_40, 
 s_89_40,  s_88_40,  s_87_40,  s_86_40,  s_85_40,  s_84_40, 
 s_83_40,  s_82_40,  s_81_40,  s_80_40
} = partial_products[(width+2)*(40+1)-1:(width+2)*40];

assign {
 s_211_0,  s_210_0,  s_209_1,  s_208_1,  s_207_2,  s_206_2, 
 s_205_3,  s_204_3,  s_203_4,  s_202_4,  s_201_5,  s_200_5, 
 s_199_6,  s_198_6,  s_197_7,  s_196_7,  s_195_8,  s_194_8, 
 s_193_9,  s_192_9, s_191_10, s_190_10, s_189_11, s_188_11, 
s_187_12, s_186_12, s_185_13, s_184_13, s_183_14, s_182_14, 
s_181_15, s_180_15, s_179_16, s_178_16, s_177_17, s_176_17, 
s_175_18, s_174_18, s_173_19, s_172_19, s_171_20, s_170_20, 
s_169_21, s_168_21, s_167_22, s_166_22, s_165_23, s_164_23, 
s_163_24, s_162_24, s_161_25, s_160_25, s_159_26, s_158_26, 
s_157_27, s_156_27, s_155_28, s_154_28, s_153_29, s_152_29, 
s_151_30, s_150_30, s_149_31, s_148_31, s_147_32, s_146_32, 
s_145_33, s_144_33, s_143_34, s_142_34, s_141_35, s_140_35, 
s_139_36, s_138_36, s_137_37, s_136_37, s_135_38, s_134_38, 
s_133_39, s_132_39, s_131_40, s_130_40, s_129_41, s_128_41, 
s_127_41, s_126_41, s_125_41, s_124_41, s_123_41, s_122_41, 
s_121_41, s_120_41, s_119_41, s_118_41, s_117_41, s_116_41, 
s_115_41, s_114_41, s_113_41, s_112_41, s_111_41, s_110_41, 
s_109_41, s_108_41, s_107_41, s_106_41, s_105_41, s_104_41, 
s_103_41, s_102_41, s_101_41, s_100_41,  s_99_41,  s_98_41, 
 s_97_41,  s_96_41,  s_95_41,  s_94_41,  s_93_41,  s_92_41, 
 s_91_41,  s_90_41,  s_89_41,  s_88_41,  s_87_41,  s_86_41, 
 s_85_41,  s_84_41,  s_83_41,  s_82_41
} = partial_products[(width+2)*(41+1)-1:(width+2)*41];

assign {
 s_213_0,  s_212_0,  s_211_1,  s_210_1,  s_209_2,  s_208_2, 
 s_207_3,  s_206_3,  s_205_4,  s_204_4,  s_203_5,  s_202_5, 
 s_201_6,  s_200_6,  s_199_7,  s_198_7,  s_197_8,  s_196_8, 
 s_195_9,  s_194_9, s_193_10, s_192_10, s_191_11, s_190_11, 
s_189_12, s_188_12, s_187_13, s_186_13, s_185_14, s_184_14, 
s_183_15, s_182_15, s_181_16, s_180_16, s_179_17, s_178_17, 
s_177_18, s_176_18, s_175_19, s_174_19, s_173_20, s_172_20, 
s_171_21, s_170_21, s_169_22, s_168_22, s_167_23, s_166_23, 
s_165_24, s_164_24, s_163_25, s_162_25, s_161_26, s_160_26, 
s_159_27, s_158_27, s_157_28, s_156_28, s_155_29, s_154_29, 
s_153_30, s_152_30, s_151_31, s_150_31, s_149_32, s_148_32, 
s_147_33, s_146_33, s_145_34, s_144_34, s_143_35, s_142_35, 
s_141_36, s_140_36, s_139_37, s_138_37, s_137_38, s_136_38, 
s_135_39, s_134_39, s_133_40, s_132_40, s_131_41, s_130_41, 
s_129_42, s_128_42, s_127_42, s_126_42, s_125_42, s_124_42, 
s_123_42, s_122_42, s_121_42, s_120_42, s_119_42, s_118_42, 
s_117_42, s_116_42, s_115_42, s_114_42, s_113_42, s_112_42, 
s_111_42, s_110_42, s_109_42, s_108_42, s_107_42, s_106_42, 
s_105_42, s_104_42, s_103_42, s_102_42, s_101_42, s_100_42, 
 s_99_42,  s_98_42,  s_97_42,  s_96_42,  s_95_42,  s_94_42, 
 s_93_42,  s_92_42,  s_91_42,  s_90_42,  s_89_42,  s_88_42, 
 s_87_42,  s_86_42,  s_85_42,  s_84_42
} = partial_products[(width+2)*(42+1)-1:(width+2)*42];

assign {
 s_215_0,  s_214_0,  s_213_1,  s_212_1,  s_211_2,  s_210_2, 
 s_209_3,  s_208_3,  s_207_4,  s_206_4,  s_205_5,  s_204_5, 
 s_203_6,  s_202_6,  s_201_7,  s_200_7,  s_199_8,  s_198_8, 
 s_197_9,  s_196_9, s_195_10, s_194_10, s_193_11, s_192_11, 
s_191_12, s_190_12, s_189_13, s_188_13, s_187_14, s_186_14, 
s_185_15, s_184_15, s_183_16, s_182_16, s_181_17, s_180_17, 
s_179_18, s_178_18, s_177_19, s_176_19, s_175_20, s_174_20, 
s_173_21, s_172_21, s_171_22, s_170_22, s_169_23, s_168_23, 
s_167_24, s_166_24, s_165_25, s_164_25, s_163_26, s_162_26, 
s_161_27, s_160_27, s_159_28, s_158_28, s_157_29, s_156_29, 
s_155_30, s_154_30, s_153_31, s_152_31, s_151_32, s_150_32, 
s_149_33, s_148_33, s_147_34, s_146_34, s_145_35, s_144_35, 
s_143_36, s_142_36, s_141_37, s_140_37, s_139_38, s_138_38, 
s_137_39, s_136_39, s_135_40, s_134_40, s_133_41, s_132_41, 
s_131_42, s_130_42, s_129_43, s_128_43, s_127_43, s_126_43, 
s_125_43, s_124_43, s_123_43, s_122_43, s_121_43, s_120_43, 
s_119_43, s_118_43, s_117_43, s_116_43, s_115_43, s_114_43, 
s_113_43, s_112_43, s_111_43, s_110_43, s_109_43, s_108_43, 
s_107_43, s_106_43, s_105_43, s_104_43, s_103_43, s_102_43, 
s_101_43, s_100_43,  s_99_43,  s_98_43,  s_97_43,  s_96_43, 
 s_95_43,  s_94_43,  s_93_43,  s_92_43,  s_91_43,  s_90_43, 
 s_89_43,  s_88_43,  s_87_43,  s_86_43
} = partial_products[(width+2)*(43+1)-1:(width+2)*43];

assign {
 s_217_0,  s_216_0,  s_215_1,  s_214_1,  s_213_2,  s_212_2, 
 s_211_3,  s_210_3,  s_209_4,  s_208_4,  s_207_5,  s_206_5, 
 s_205_6,  s_204_6,  s_203_7,  s_202_7,  s_201_8,  s_200_8, 
 s_199_9,  s_198_9, s_197_10, s_196_10, s_195_11, s_194_11, 
s_193_12, s_192_12, s_191_13, s_190_13, s_189_14, s_188_14, 
s_187_15, s_186_15, s_185_16, s_184_16, s_183_17, s_182_17, 
s_181_18, s_180_18, s_179_19, s_178_19, s_177_20, s_176_20, 
s_175_21, s_174_21, s_173_22, s_172_22, s_171_23, s_170_23, 
s_169_24, s_168_24, s_167_25, s_166_25, s_165_26, s_164_26, 
s_163_27, s_162_27, s_161_28, s_160_28, s_159_29, s_158_29, 
s_157_30, s_156_30, s_155_31, s_154_31, s_153_32, s_152_32, 
s_151_33, s_150_33, s_149_34, s_148_34, s_147_35, s_146_35, 
s_145_36, s_144_36, s_143_37, s_142_37, s_141_38, s_140_38, 
s_139_39, s_138_39, s_137_40, s_136_40, s_135_41, s_134_41, 
s_133_42, s_132_42, s_131_43, s_130_43, s_129_44, s_128_44, 
s_127_44, s_126_44, s_125_44, s_124_44, s_123_44, s_122_44, 
s_121_44, s_120_44, s_119_44, s_118_44, s_117_44, s_116_44, 
s_115_44, s_114_44, s_113_44, s_112_44, s_111_44, s_110_44, 
s_109_44, s_108_44, s_107_44, s_106_44, s_105_44, s_104_44, 
s_103_44, s_102_44, s_101_44, s_100_44,  s_99_44,  s_98_44, 
 s_97_44,  s_96_44,  s_95_44,  s_94_44,  s_93_44,  s_92_44, 
 s_91_44,  s_90_44,  s_89_44,  s_88_44
} = partial_products[(width+2)*(44+1)-1:(width+2)*44];

assign {
 s_219_0,  s_218_0,  s_217_1,  s_216_1,  s_215_2,  s_214_2, 
 s_213_3,  s_212_3,  s_211_4,  s_210_4,  s_209_5,  s_208_5, 
 s_207_6,  s_206_6,  s_205_7,  s_204_7,  s_203_8,  s_202_8, 
 s_201_9,  s_200_9, s_199_10, s_198_10, s_197_11, s_196_11, 
s_195_12, s_194_12, s_193_13, s_192_13, s_191_14, s_190_14, 
s_189_15, s_188_15, s_187_16, s_186_16, s_185_17, s_184_17, 
s_183_18, s_182_18, s_181_19, s_180_19, s_179_20, s_178_20, 
s_177_21, s_176_21, s_175_22, s_174_22, s_173_23, s_172_23, 
s_171_24, s_170_24, s_169_25, s_168_25, s_167_26, s_166_26, 
s_165_27, s_164_27, s_163_28, s_162_28, s_161_29, s_160_29, 
s_159_30, s_158_30, s_157_31, s_156_31, s_155_32, s_154_32, 
s_153_33, s_152_33, s_151_34, s_150_34, s_149_35, s_148_35, 
s_147_36, s_146_36, s_145_37, s_144_37, s_143_38, s_142_38, 
s_141_39, s_140_39, s_139_40, s_138_40, s_137_41, s_136_41, 
s_135_42, s_134_42, s_133_43, s_132_43, s_131_44, s_130_44, 
s_129_45, s_128_45, s_127_45, s_126_45, s_125_45, s_124_45, 
s_123_45, s_122_45, s_121_45, s_120_45, s_119_45, s_118_45, 
s_117_45, s_116_45, s_115_45, s_114_45, s_113_45, s_112_45, 
s_111_45, s_110_45, s_109_45, s_108_45, s_107_45, s_106_45, 
s_105_45, s_104_45, s_103_45, s_102_45, s_101_45, s_100_45, 
 s_99_45,  s_98_45,  s_97_45,  s_96_45,  s_95_45,  s_94_45, 
 s_93_45,  s_92_45,  s_91_45,  s_90_45
} = partial_products[(width+2)*(45+1)-1:(width+2)*45];

assign {
 s_221_0,  s_220_0,  s_219_1,  s_218_1,  s_217_2,  s_216_2, 
 s_215_3,  s_214_3,  s_213_4,  s_212_4,  s_211_5,  s_210_5, 
 s_209_6,  s_208_6,  s_207_7,  s_206_7,  s_205_8,  s_204_8, 
 s_203_9,  s_202_9, s_201_10, s_200_10, s_199_11, s_198_11, 
s_197_12, s_196_12, s_195_13, s_194_13, s_193_14, s_192_14, 
s_191_15, s_190_15, s_189_16, s_188_16, s_187_17, s_186_17, 
s_185_18, s_184_18, s_183_19, s_182_19, s_181_20, s_180_20, 
s_179_21, s_178_21, s_177_22, s_176_22, s_175_23, s_174_23, 
s_173_24, s_172_24, s_171_25, s_170_25, s_169_26, s_168_26, 
s_167_27, s_166_27, s_165_28, s_164_28, s_163_29, s_162_29, 
s_161_30, s_160_30, s_159_31, s_158_31, s_157_32, s_156_32, 
s_155_33, s_154_33, s_153_34, s_152_34, s_151_35, s_150_35, 
s_149_36, s_148_36, s_147_37, s_146_37, s_145_38, s_144_38, 
s_143_39, s_142_39, s_141_40, s_140_40, s_139_41, s_138_41, 
s_137_42, s_136_42, s_135_43, s_134_43, s_133_44, s_132_44, 
s_131_45, s_130_45, s_129_46, s_128_46, s_127_46, s_126_46, 
s_125_46, s_124_46, s_123_46, s_122_46, s_121_46, s_120_46, 
s_119_46, s_118_46, s_117_46, s_116_46, s_115_46, s_114_46, 
s_113_46, s_112_46, s_111_46, s_110_46, s_109_46, s_108_46, 
s_107_46, s_106_46, s_105_46, s_104_46, s_103_46, s_102_46, 
s_101_46, s_100_46,  s_99_46,  s_98_46,  s_97_46,  s_96_46, 
 s_95_46,  s_94_46,  s_93_46,  s_92_46
} = partial_products[(width+2)*(46+1)-1:(width+2)*46];

assign {
 s_223_0,  s_222_0,  s_221_1,  s_220_1,  s_219_2,  s_218_2, 
 s_217_3,  s_216_3,  s_215_4,  s_214_4,  s_213_5,  s_212_5, 
 s_211_6,  s_210_6,  s_209_7,  s_208_7,  s_207_8,  s_206_8, 
 s_205_9,  s_204_9, s_203_10, s_202_10, s_201_11, s_200_11, 
s_199_12, s_198_12, s_197_13, s_196_13, s_195_14, s_194_14, 
s_193_15, s_192_15, s_191_16, s_190_16, s_189_17, s_188_17, 
s_187_18, s_186_18, s_185_19, s_184_19, s_183_20, s_182_20, 
s_181_21, s_180_21, s_179_22, s_178_22, s_177_23, s_176_23, 
s_175_24, s_174_24, s_173_25, s_172_25, s_171_26, s_170_26, 
s_169_27, s_168_27, s_167_28, s_166_28, s_165_29, s_164_29, 
s_163_30, s_162_30, s_161_31, s_160_31, s_159_32, s_158_32, 
s_157_33, s_156_33, s_155_34, s_154_34, s_153_35, s_152_35, 
s_151_36, s_150_36, s_149_37, s_148_37, s_147_38, s_146_38, 
s_145_39, s_144_39, s_143_40, s_142_40, s_141_41, s_140_41, 
s_139_42, s_138_42, s_137_43, s_136_43, s_135_44, s_134_44, 
s_133_45, s_132_45, s_131_46, s_130_46, s_129_47, s_128_47, 
s_127_47, s_126_47, s_125_47, s_124_47, s_123_47, s_122_47, 
s_121_47, s_120_47, s_119_47, s_118_47, s_117_47, s_116_47, 
s_115_47, s_114_47, s_113_47, s_112_47, s_111_47, s_110_47, 
s_109_47, s_108_47, s_107_47, s_106_47, s_105_47, s_104_47, 
s_103_47, s_102_47, s_101_47, s_100_47,  s_99_47,  s_98_47, 
 s_97_47,  s_96_47,  s_95_47,  s_94_47
} = partial_products[(width+2)*(47+1)-1:(width+2)*47];

assign {
 s_225_0,  s_224_0,  s_223_1,  s_222_1,  s_221_2,  s_220_2, 
 s_219_3,  s_218_3,  s_217_4,  s_216_4,  s_215_5,  s_214_5, 
 s_213_6,  s_212_6,  s_211_7,  s_210_7,  s_209_8,  s_208_8, 
 s_207_9,  s_206_9, s_205_10, s_204_10, s_203_11, s_202_11, 
s_201_12, s_200_12, s_199_13, s_198_13, s_197_14, s_196_14, 
s_195_15, s_194_15, s_193_16, s_192_16, s_191_17, s_190_17, 
s_189_18, s_188_18, s_187_19, s_186_19, s_185_20, s_184_20, 
s_183_21, s_182_21, s_181_22, s_180_22, s_179_23, s_178_23, 
s_177_24, s_176_24, s_175_25, s_174_25, s_173_26, s_172_26, 
s_171_27, s_170_27, s_169_28, s_168_28, s_167_29, s_166_29, 
s_165_30, s_164_30, s_163_31, s_162_31, s_161_32, s_160_32, 
s_159_33, s_158_33, s_157_34, s_156_34, s_155_35, s_154_35, 
s_153_36, s_152_36, s_151_37, s_150_37, s_149_38, s_148_38, 
s_147_39, s_146_39, s_145_40, s_144_40, s_143_41, s_142_41, 
s_141_42, s_140_42, s_139_43, s_138_43, s_137_44, s_136_44, 
s_135_45, s_134_45, s_133_46, s_132_46, s_131_47, s_130_47, 
s_129_48, s_128_48, s_127_48, s_126_48, s_125_48, s_124_48, 
s_123_48, s_122_48, s_121_48, s_120_48, s_119_48, s_118_48, 
s_117_48, s_116_48, s_115_48, s_114_48, s_113_48, s_112_48, 
s_111_48, s_110_48, s_109_48, s_108_48, s_107_48, s_106_48, 
s_105_48, s_104_48, s_103_48, s_102_48, s_101_48, s_100_48, 
 s_99_48,  s_98_48,  s_97_48,  s_96_48
} = partial_products[(width+2)*(48+1)-1:(width+2)*48];

assign {
 s_227_0,  s_226_0,  s_225_1,  s_224_1,  s_223_2,  s_222_2, 
 s_221_3,  s_220_3,  s_219_4,  s_218_4,  s_217_5,  s_216_5, 
 s_215_6,  s_214_6,  s_213_7,  s_212_7,  s_211_8,  s_210_8, 
 s_209_9,  s_208_9, s_207_10, s_206_10, s_205_11, s_204_11, 
s_203_12, s_202_12, s_201_13, s_200_13, s_199_14, s_198_14, 
s_197_15, s_196_15, s_195_16, s_194_16, s_193_17, s_192_17, 
s_191_18, s_190_18, s_189_19, s_188_19, s_187_20, s_186_20, 
s_185_21, s_184_21, s_183_22, s_182_22, s_181_23, s_180_23, 
s_179_24, s_178_24, s_177_25, s_176_25, s_175_26, s_174_26, 
s_173_27, s_172_27, s_171_28, s_170_28, s_169_29, s_168_29, 
s_167_30, s_166_30, s_165_31, s_164_31, s_163_32, s_162_32, 
s_161_33, s_160_33, s_159_34, s_158_34, s_157_35, s_156_35, 
s_155_36, s_154_36, s_153_37, s_152_37, s_151_38, s_150_38, 
s_149_39, s_148_39, s_147_40, s_146_40, s_145_41, s_144_41, 
s_143_42, s_142_42, s_141_43, s_140_43, s_139_44, s_138_44, 
s_137_45, s_136_45, s_135_46, s_134_46, s_133_47, s_132_47, 
s_131_48, s_130_48, s_129_49, s_128_49, s_127_49, s_126_49, 
s_125_49, s_124_49, s_123_49, s_122_49, s_121_49, s_120_49, 
s_119_49, s_118_49, s_117_49, s_116_49, s_115_49, s_114_49, 
s_113_49, s_112_49, s_111_49, s_110_49, s_109_49, s_108_49, 
s_107_49, s_106_49, s_105_49, s_104_49, s_103_49, s_102_49, 
s_101_49, s_100_49,  s_99_49,  s_98_49
} = partial_products[(width+2)*(49+1)-1:(width+2)*49];

assign {
 s_229_0,  s_228_0,  s_227_1,  s_226_1,  s_225_2,  s_224_2, 
 s_223_3,  s_222_3,  s_221_4,  s_220_4,  s_219_5,  s_218_5, 
 s_217_6,  s_216_6,  s_215_7,  s_214_7,  s_213_8,  s_212_8, 
 s_211_9,  s_210_9, s_209_10, s_208_10, s_207_11, s_206_11, 
s_205_12, s_204_12, s_203_13, s_202_13, s_201_14, s_200_14, 
s_199_15, s_198_15, s_197_16, s_196_16, s_195_17, s_194_17, 
s_193_18, s_192_18, s_191_19, s_190_19, s_189_20, s_188_20, 
s_187_21, s_186_21, s_185_22, s_184_22, s_183_23, s_182_23, 
s_181_24, s_180_24, s_179_25, s_178_25, s_177_26, s_176_26, 
s_175_27, s_174_27, s_173_28, s_172_28, s_171_29, s_170_29, 
s_169_30, s_168_30, s_167_31, s_166_31, s_165_32, s_164_32, 
s_163_33, s_162_33, s_161_34, s_160_34, s_159_35, s_158_35, 
s_157_36, s_156_36, s_155_37, s_154_37, s_153_38, s_152_38, 
s_151_39, s_150_39, s_149_40, s_148_40, s_147_41, s_146_41, 
s_145_42, s_144_42, s_143_43, s_142_43, s_141_44, s_140_44, 
s_139_45, s_138_45, s_137_46, s_136_46, s_135_47, s_134_47, 
s_133_48, s_132_48, s_131_49, s_130_49, s_129_50, s_128_50, 
s_127_50, s_126_50, s_125_50, s_124_50, s_123_50, s_122_50, 
s_121_50, s_120_50, s_119_50, s_118_50, s_117_50, s_116_50, 
s_115_50, s_114_50, s_113_50, s_112_50, s_111_50, s_110_50, 
s_109_50, s_108_50, s_107_50, s_106_50, s_105_50, s_104_50, 
s_103_50, s_102_50, s_101_50, s_100_50
} = partial_products[(width+2)*(50+1)-1:(width+2)*50];

assign {
 s_231_0,  s_230_0,  s_229_1,  s_228_1,  s_227_2,  s_226_2, 
 s_225_3,  s_224_3,  s_223_4,  s_222_4,  s_221_5,  s_220_5, 
 s_219_6,  s_218_6,  s_217_7,  s_216_7,  s_215_8,  s_214_8, 
 s_213_9,  s_212_9, s_211_10, s_210_10, s_209_11, s_208_11, 
s_207_12, s_206_12, s_205_13, s_204_13, s_203_14, s_202_14, 
s_201_15, s_200_15, s_199_16, s_198_16, s_197_17, s_196_17, 
s_195_18, s_194_18, s_193_19, s_192_19, s_191_20, s_190_20, 
s_189_21, s_188_21, s_187_22, s_186_22, s_185_23, s_184_23, 
s_183_24, s_182_24, s_181_25, s_180_25, s_179_26, s_178_26, 
s_177_27, s_176_27, s_175_28, s_174_28, s_173_29, s_172_29, 
s_171_30, s_170_30, s_169_31, s_168_31, s_167_32, s_166_32, 
s_165_33, s_164_33, s_163_34, s_162_34, s_161_35, s_160_35, 
s_159_36, s_158_36, s_157_37, s_156_37, s_155_38, s_154_38, 
s_153_39, s_152_39, s_151_40, s_150_40, s_149_41, s_148_41, 
s_147_42, s_146_42, s_145_43, s_144_43, s_143_44, s_142_44, 
s_141_45, s_140_45, s_139_46, s_138_46, s_137_47, s_136_47, 
s_135_48, s_134_48, s_133_49, s_132_49, s_131_50, s_130_50, 
s_129_51, s_128_51, s_127_51, s_126_51, s_125_51, s_124_51, 
s_123_51, s_122_51, s_121_51, s_120_51, s_119_51, s_118_51, 
s_117_51, s_116_51, s_115_51, s_114_51, s_113_51, s_112_51, 
s_111_51, s_110_51, s_109_51, s_108_51, s_107_51, s_106_51, 
s_105_51, s_104_51, s_103_51, s_102_51
} = partial_products[(width+2)*(51+1)-1:(width+2)*51];

assign {
 s_233_0,  s_232_0,  s_231_1,  s_230_1,  s_229_2,  s_228_2, 
 s_227_3,  s_226_3,  s_225_4,  s_224_4,  s_223_5,  s_222_5, 
 s_221_6,  s_220_6,  s_219_7,  s_218_7,  s_217_8,  s_216_8, 
 s_215_9,  s_214_9, s_213_10, s_212_10, s_211_11, s_210_11, 
s_209_12, s_208_12, s_207_13, s_206_13, s_205_14, s_204_14, 
s_203_15, s_202_15, s_201_16, s_200_16, s_199_17, s_198_17, 
s_197_18, s_196_18, s_195_19, s_194_19, s_193_20, s_192_20, 
s_191_21, s_190_21, s_189_22, s_188_22, s_187_23, s_186_23, 
s_185_24, s_184_24, s_183_25, s_182_25, s_181_26, s_180_26, 
s_179_27, s_178_27, s_177_28, s_176_28, s_175_29, s_174_29, 
s_173_30, s_172_30, s_171_31, s_170_31, s_169_32, s_168_32, 
s_167_33, s_166_33, s_165_34, s_164_34, s_163_35, s_162_35, 
s_161_36, s_160_36, s_159_37, s_158_37, s_157_38, s_156_38, 
s_155_39, s_154_39, s_153_40, s_152_40, s_151_41, s_150_41, 
s_149_42, s_148_42, s_147_43, s_146_43, s_145_44, s_144_44, 
s_143_45, s_142_45, s_141_46, s_140_46, s_139_47, s_138_47, 
s_137_48, s_136_48, s_135_49, s_134_49, s_133_50, s_132_50, 
s_131_51, s_130_51, s_129_52, s_128_52, s_127_52, s_126_52, 
s_125_52, s_124_52, s_123_52, s_122_52, s_121_52, s_120_52, 
s_119_52, s_118_52, s_117_52, s_116_52, s_115_52, s_114_52, 
s_113_52, s_112_52, s_111_52, s_110_52, s_109_52, s_108_52, 
s_107_52, s_106_52, s_105_52, s_104_52
} = partial_products[(width+2)*(52+1)-1:(width+2)*52];

assign {
 s_235_0,  s_234_0,  s_233_1,  s_232_1,  s_231_2,  s_230_2, 
 s_229_3,  s_228_3,  s_227_4,  s_226_4,  s_225_5,  s_224_5, 
 s_223_6,  s_222_6,  s_221_7,  s_220_7,  s_219_8,  s_218_8, 
 s_217_9,  s_216_9, s_215_10, s_214_10, s_213_11, s_212_11, 
s_211_12, s_210_12, s_209_13, s_208_13, s_207_14, s_206_14, 
s_205_15, s_204_15, s_203_16, s_202_16, s_201_17, s_200_17, 
s_199_18, s_198_18, s_197_19, s_196_19, s_195_20, s_194_20, 
s_193_21, s_192_21, s_191_22, s_190_22, s_189_23, s_188_23, 
s_187_24, s_186_24, s_185_25, s_184_25, s_183_26, s_182_26, 
s_181_27, s_180_27, s_179_28, s_178_28, s_177_29, s_176_29, 
s_175_30, s_174_30, s_173_31, s_172_31, s_171_32, s_170_32, 
s_169_33, s_168_33, s_167_34, s_166_34, s_165_35, s_164_35, 
s_163_36, s_162_36, s_161_37, s_160_37, s_159_38, s_158_38, 
s_157_39, s_156_39, s_155_40, s_154_40, s_153_41, s_152_41, 
s_151_42, s_150_42, s_149_43, s_148_43, s_147_44, s_146_44, 
s_145_45, s_144_45, s_143_46, s_142_46, s_141_47, s_140_47, 
s_139_48, s_138_48, s_137_49, s_136_49, s_135_50, s_134_50, 
s_133_51, s_132_51, s_131_52, s_130_52, s_129_53, s_128_53, 
s_127_53, s_126_53, s_125_53, s_124_53, s_123_53, s_122_53, 
s_121_53, s_120_53, s_119_53, s_118_53, s_117_53, s_116_53, 
s_115_53, s_114_53, s_113_53, s_112_53, s_111_53, s_110_53, 
s_109_53, s_108_53, s_107_53, s_106_53
} = partial_products[(width+2)*(53+1)-1:(width+2)*53];

assign {
 s_237_0,  s_236_0,  s_235_1,  s_234_1,  s_233_2,  s_232_2, 
 s_231_3,  s_230_3,  s_229_4,  s_228_4,  s_227_5,  s_226_5, 
 s_225_6,  s_224_6,  s_223_7,  s_222_7,  s_221_8,  s_220_8, 
 s_219_9,  s_218_9, s_217_10, s_216_10, s_215_11, s_214_11, 
s_213_12, s_212_12, s_211_13, s_210_13, s_209_14, s_208_14, 
s_207_15, s_206_15, s_205_16, s_204_16, s_203_17, s_202_17, 
s_201_18, s_200_18, s_199_19, s_198_19, s_197_20, s_196_20, 
s_195_21, s_194_21, s_193_22, s_192_22, s_191_23, s_190_23, 
s_189_24, s_188_24, s_187_25, s_186_25, s_185_26, s_184_26, 
s_183_27, s_182_27, s_181_28, s_180_28, s_179_29, s_178_29, 
s_177_30, s_176_30, s_175_31, s_174_31, s_173_32, s_172_32, 
s_171_33, s_170_33, s_169_34, s_168_34, s_167_35, s_166_35, 
s_165_36, s_164_36, s_163_37, s_162_37, s_161_38, s_160_38, 
s_159_39, s_158_39, s_157_40, s_156_40, s_155_41, s_154_41, 
s_153_42, s_152_42, s_151_43, s_150_43, s_149_44, s_148_44, 
s_147_45, s_146_45, s_145_46, s_144_46, s_143_47, s_142_47, 
s_141_48, s_140_48, s_139_49, s_138_49, s_137_50, s_136_50, 
s_135_51, s_134_51, s_133_52, s_132_52, s_131_53, s_130_53, 
s_129_54, s_128_54, s_127_54, s_126_54, s_125_54, s_124_54, 
s_123_54, s_122_54, s_121_54, s_120_54, s_119_54, s_118_54, 
s_117_54, s_116_54, s_115_54, s_114_54, s_113_54, s_112_54, 
s_111_54, s_110_54, s_109_54, s_108_54
} = partial_products[(width+2)*(54+1)-1:(width+2)*54];

assign {
 s_239_0,  s_238_0,  s_237_1,  s_236_1,  s_235_2,  s_234_2, 
 s_233_3,  s_232_3,  s_231_4,  s_230_4,  s_229_5,  s_228_5, 
 s_227_6,  s_226_6,  s_225_7,  s_224_7,  s_223_8,  s_222_8, 
 s_221_9,  s_220_9, s_219_10, s_218_10, s_217_11, s_216_11, 
s_215_12, s_214_12, s_213_13, s_212_13, s_211_14, s_210_14, 
s_209_15, s_208_15, s_207_16, s_206_16, s_205_17, s_204_17, 
s_203_18, s_202_18, s_201_19, s_200_19, s_199_20, s_198_20, 
s_197_21, s_196_21, s_195_22, s_194_22, s_193_23, s_192_23, 
s_191_24, s_190_24, s_189_25, s_188_25, s_187_26, s_186_26, 
s_185_27, s_184_27, s_183_28, s_182_28, s_181_29, s_180_29, 
s_179_30, s_178_30, s_177_31, s_176_31, s_175_32, s_174_32, 
s_173_33, s_172_33, s_171_34, s_170_34, s_169_35, s_168_35, 
s_167_36, s_166_36, s_165_37, s_164_37, s_163_38, s_162_38, 
s_161_39, s_160_39, s_159_40, s_158_40, s_157_41, s_156_41, 
s_155_42, s_154_42, s_153_43, s_152_43, s_151_44, s_150_44, 
s_149_45, s_148_45, s_147_46, s_146_46, s_145_47, s_144_47, 
s_143_48, s_142_48, s_141_49, s_140_49, s_139_50, s_138_50, 
s_137_51, s_136_51, s_135_52, s_134_52, s_133_53, s_132_53, 
s_131_54, s_130_54, s_129_55, s_128_55, s_127_55, s_126_55, 
s_125_55, s_124_55, s_123_55, s_122_55, s_121_55, s_120_55, 
s_119_55, s_118_55, s_117_55, s_116_55, s_115_55, s_114_55, 
s_113_55, s_112_55, s_111_55, s_110_55
} = partial_products[(width+2)*(55+1)-1:(width+2)*55];

assign {
 s_241_0,  s_240_0,  s_239_1,  s_238_1,  s_237_2,  s_236_2, 
 s_235_3,  s_234_3,  s_233_4,  s_232_4,  s_231_5,  s_230_5, 
 s_229_6,  s_228_6,  s_227_7,  s_226_7,  s_225_8,  s_224_8, 
 s_223_9,  s_222_9, s_221_10, s_220_10, s_219_11, s_218_11, 
s_217_12, s_216_12, s_215_13, s_214_13, s_213_14, s_212_14, 
s_211_15, s_210_15, s_209_16, s_208_16, s_207_17, s_206_17, 
s_205_18, s_204_18, s_203_19, s_202_19, s_201_20, s_200_20, 
s_199_21, s_198_21, s_197_22, s_196_22, s_195_23, s_194_23, 
s_193_24, s_192_24, s_191_25, s_190_25, s_189_26, s_188_26, 
s_187_27, s_186_27, s_185_28, s_184_28, s_183_29, s_182_29, 
s_181_30, s_180_30, s_179_31, s_178_31, s_177_32, s_176_32, 
s_175_33, s_174_33, s_173_34, s_172_34, s_171_35, s_170_35, 
s_169_36, s_168_36, s_167_37, s_166_37, s_165_38, s_164_38, 
s_163_39, s_162_39, s_161_40, s_160_40, s_159_41, s_158_41, 
s_157_42, s_156_42, s_155_43, s_154_43, s_153_44, s_152_44, 
s_151_45, s_150_45, s_149_46, s_148_46, s_147_47, s_146_47, 
s_145_48, s_144_48, s_143_49, s_142_49, s_141_50, s_140_50, 
s_139_51, s_138_51, s_137_52, s_136_52, s_135_53, s_134_53, 
s_133_54, s_132_54, s_131_55, s_130_55, s_129_56, s_128_56, 
s_127_56, s_126_56, s_125_56, s_124_56, s_123_56, s_122_56, 
s_121_56, s_120_56, s_119_56, s_118_56, s_117_56, s_116_56, 
s_115_56, s_114_56, s_113_56, s_112_56
} = partial_products[(width+2)*(56+1)-1:(width+2)*56];

assign {
 s_243_0,  s_242_0,  s_241_1,  s_240_1,  s_239_2,  s_238_2, 
 s_237_3,  s_236_3,  s_235_4,  s_234_4,  s_233_5,  s_232_5, 
 s_231_6,  s_230_6,  s_229_7,  s_228_7,  s_227_8,  s_226_8, 
 s_225_9,  s_224_9, s_223_10, s_222_10, s_221_11, s_220_11, 
s_219_12, s_218_12, s_217_13, s_216_13, s_215_14, s_214_14, 
s_213_15, s_212_15, s_211_16, s_210_16, s_209_17, s_208_17, 
s_207_18, s_206_18, s_205_19, s_204_19, s_203_20, s_202_20, 
s_201_21, s_200_21, s_199_22, s_198_22, s_197_23, s_196_23, 
s_195_24, s_194_24, s_193_25, s_192_25, s_191_26, s_190_26, 
s_189_27, s_188_27, s_187_28, s_186_28, s_185_29, s_184_29, 
s_183_30, s_182_30, s_181_31, s_180_31, s_179_32, s_178_32, 
s_177_33, s_176_33, s_175_34, s_174_34, s_173_35, s_172_35, 
s_171_36, s_170_36, s_169_37, s_168_37, s_167_38, s_166_38, 
s_165_39, s_164_39, s_163_40, s_162_40, s_161_41, s_160_41, 
s_159_42, s_158_42, s_157_43, s_156_43, s_155_44, s_154_44, 
s_153_45, s_152_45, s_151_46, s_150_46, s_149_47, s_148_47, 
s_147_48, s_146_48, s_145_49, s_144_49, s_143_50, s_142_50, 
s_141_51, s_140_51, s_139_52, s_138_52, s_137_53, s_136_53, 
s_135_54, s_134_54, s_133_55, s_132_55, s_131_56, s_130_56, 
s_129_57, s_128_57, s_127_57, s_126_57, s_125_57, s_124_57, 
s_123_57, s_122_57, s_121_57, s_120_57, s_119_57, s_118_57, 
s_117_57, s_116_57, s_115_57, s_114_57
} = partial_products[(width+2)*(57+1)-1:(width+2)*57];

assign {
 s_245_0,  s_244_0,  s_243_1,  s_242_1,  s_241_2,  s_240_2, 
 s_239_3,  s_238_3,  s_237_4,  s_236_4,  s_235_5,  s_234_5, 
 s_233_6,  s_232_6,  s_231_7,  s_230_7,  s_229_8,  s_228_8, 
 s_227_9,  s_226_9, s_225_10, s_224_10, s_223_11, s_222_11, 
s_221_12, s_220_12, s_219_13, s_218_13, s_217_14, s_216_14, 
s_215_15, s_214_15, s_213_16, s_212_16, s_211_17, s_210_17, 
s_209_18, s_208_18, s_207_19, s_206_19, s_205_20, s_204_20, 
s_203_21, s_202_21, s_201_22, s_200_22, s_199_23, s_198_23, 
s_197_24, s_196_24, s_195_25, s_194_25, s_193_26, s_192_26, 
s_191_27, s_190_27, s_189_28, s_188_28, s_187_29, s_186_29, 
s_185_30, s_184_30, s_183_31, s_182_31, s_181_32, s_180_32, 
s_179_33, s_178_33, s_177_34, s_176_34, s_175_35, s_174_35, 
s_173_36, s_172_36, s_171_37, s_170_37, s_169_38, s_168_38, 
s_167_39, s_166_39, s_165_40, s_164_40, s_163_41, s_162_41, 
s_161_42, s_160_42, s_159_43, s_158_43, s_157_44, s_156_44, 
s_155_45, s_154_45, s_153_46, s_152_46, s_151_47, s_150_47, 
s_149_48, s_148_48, s_147_49, s_146_49, s_145_50, s_144_50, 
s_143_51, s_142_51, s_141_52, s_140_52, s_139_53, s_138_53, 
s_137_54, s_136_54, s_135_55, s_134_55, s_133_56, s_132_56, 
s_131_57, s_130_57, s_129_58, s_128_58, s_127_58, s_126_58, 
s_125_58, s_124_58, s_123_58, s_122_58, s_121_58, s_120_58, 
s_119_58, s_118_58, s_117_58, s_116_58
} = partial_products[(width+2)*(58+1)-1:(width+2)*58];

assign {
 s_247_0,  s_246_0,  s_245_1,  s_244_1,  s_243_2,  s_242_2, 
 s_241_3,  s_240_3,  s_239_4,  s_238_4,  s_237_5,  s_236_5, 
 s_235_6,  s_234_6,  s_233_7,  s_232_7,  s_231_8,  s_230_8, 
 s_229_9,  s_228_9, s_227_10, s_226_10, s_225_11, s_224_11, 
s_223_12, s_222_12, s_221_13, s_220_13, s_219_14, s_218_14, 
s_217_15, s_216_15, s_215_16, s_214_16, s_213_17, s_212_17, 
s_211_18, s_210_18, s_209_19, s_208_19, s_207_20, s_206_20, 
s_205_21, s_204_21, s_203_22, s_202_22, s_201_23, s_200_23, 
s_199_24, s_198_24, s_197_25, s_196_25, s_195_26, s_194_26, 
s_193_27, s_192_27, s_191_28, s_190_28, s_189_29, s_188_29, 
s_187_30, s_186_30, s_185_31, s_184_31, s_183_32, s_182_32, 
s_181_33, s_180_33, s_179_34, s_178_34, s_177_35, s_176_35, 
s_175_36, s_174_36, s_173_37, s_172_37, s_171_38, s_170_38, 
s_169_39, s_168_39, s_167_40, s_166_40, s_165_41, s_164_41, 
s_163_42, s_162_42, s_161_43, s_160_43, s_159_44, s_158_44, 
s_157_45, s_156_45, s_155_46, s_154_46, s_153_47, s_152_47, 
s_151_48, s_150_48, s_149_49, s_148_49, s_147_50, s_146_50, 
s_145_51, s_144_51, s_143_52, s_142_52, s_141_53, s_140_53, 
s_139_54, s_138_54, s_137_55, s_136_55, s_135_56, s_134_56, 
s_133_57, s_132_57, s_131_58, s_130_58, s_129_59, s_128_59, 
s_127_59, s_126_59, s_125_59, s_124_59, s_123_59, s_122_59, 
s_121_59, s_120_59, s_119_59, s_118_59
} = partial_products[(width+2)*(59+1)-1:(width+2)*59];

assign {
 s_249_0,  s_248_0,  s_247_1,  s_246_1,  s_245_2,  s_244_2, 
 s_243_3,  s_242_3,  s_241_4,  s_240_4,  s_239_5,  s_238_5, 
 s_237_6,  s_236_6,  s_235_7,  s_234_7,  s_233_8,  s_232_8, 
 s_231_9,  s_230_9, s_229_10, s_228_10, s_227_11, s_226_11, 
s_225_12, s_224_12, s_223_13, s_222_13, s_221_14, s_220_14, 
s_219_15, s_218_15, s_217_16, s_216_16, s_215_17, s_214_17, 
s_213_18, s_212_18, s_211_19, s_210_19, s_209_20, s_208_20, 
s_207_21, s_206_21, s_205_22, s_204_22, s_203_23, s_202_23, 
s_201_24, s_200_24, s_199_25, s_198_25, s_197_26, s_196_26, 
s_195_27, s_194_27, s_193_28, s_192_28, s_191_29, s_190_29, 
s_189_30, s_188_30, s_187_31, s_186_31, s_185_32, s_184_32, 
s_183_33, s_182_33, s_181_34, s_180_34, s_179_35, s_178_35, 
s_177_36, s_176_36, s_175_37, s_174_37, s_173_38, s_172_38, 
s_171_39, s_170_39, s_169_40, s_168_40, s_167_41, s_166_41, 
s_165_42, s_164_42, s_163_43, s_162_43, s_161_44, s_160_44, 
s_159_45, s_158_45, s_157_46, s_156_46, s_155_47, s_154_47, 
s_153_48, s_152_48, s_151_49, s_150_49, s_149_50, s_148_50, 
s_147_51, s_146_51, s_145_52, s_144_52, s_143_53, s_142_53, 
s_141_54, s_140_54, s_139_55, s_138_55, s_137_56, s_136_56, 
s_135_57, s_134_57, s_133_58, s_132_58, s_131_59, s_130_59, 
s_129_60, s_128_60, s_127_60, s_126_60, s_125_60, s_124_60, 
s_123_60, s_122_60, s_121_60, s_120_60
} = partial_products[(width+2)*(60+1)-1:(width+2)*60];

assign {
 s_251_0,  s_250_0,  s_249_1,  s_248_1,  s_247_2,  s_246_2, 
 s_245_3,  s_244_3,  s_243_4,  s_242_4,  s_241_5,  s_240_5, 
 s_239_6,  s_238_6,  s_237_7,  s_236_7,  s_235_8,  s_234_8, 
 s_233_9,  s_232_9, s_231_10, s_230_10, s_229_11, s_228_11, 
s_227_12, s_226_12, s_225_13, s_224_13, s_223_14, s_222_14, 
s_221_15, s_220_15, s_219_16, s_218_16, s_217_17, s_216_17, 
s_215_18, s_214_18, s_213_19, s_212_19, s_211_20, s_210_20, 
s_209_21, s_208_21, s_207_22, s_206_22, s_205_23, s_204_23, 
s_203_24, s_202_24, s_201_25, s_200_25, s_199_26, s_198_26, 
s_197_27, s_196_27, s_195_28, s_194_28, s_193_29, s_192_29, 
s_191_30, s_190_30, s_189_31, s_188_31, s_187_32, s_186_32, 
s_185_33, s_184_33, s_183_34, s_182_34, s_181_35, s_180_35, 
s_179_36, s_178_36, s_177_37, s_176_37, s_175_38, s_174_38, 
s_173_39, s_172_39, s_171_40, s_170_40, s_169_41, s_168_41, 
s_167_42, s_166_42, s_165_43, s_164_43, s_163_44, s_162_44, 
s_161_45, s_160_45, s_159_46, s_158_46, s_157_47, s_156_47, 
s_155_48, s_154_48, s_153_49, s_152_49, s_151_50, s_150_50, 
s_149_51, s_148_51, s_147_52, s_146_52, s_145_53, s_144_53, 
s_143_54, s_142_54, s_141_55, s_140_55, s_139_56, s_138_56, 
s_137_57, s_136_57, s_135_58, s_134_58, s_133_59, s_132_59, 
s_131_60, s_130_60, s_129_61, s_128_61, s_127_61, s_126_61, 
s_125_61, s_124_61, s_123_61, s_122_61
} = partial_products[(width+2)*(61+1)-1:(width+2)*61];

assign {
 s_253_0,  s_252_0,  s_251_1,  s_250_1,  s_249_2,  s_248_2, 
 s_247_3,  s_246_3,  s_245_4,  s_244_4,  s_243_5,  s_242_5, 
 s_241_6,  s_240_6,  s_239_7,  s_238_7,  s_237_8,  s_236_8, 
 s_235_9,  s_234_9, s_233_10, s_232_10, s_231_11, s_230_11, 
s_229_12, s_228_12, s_227_13, s_226_13, s_225_14, s_224_14, 
s_223_15, s_222_15, s_221_16, s_220_16, s_219_17, s_218_17, 
s_217_18, s_216_18, s_215_19, s_214_19, s_213_20, s_212_20, 
s_211_21, s_210_21, s_209_22, s_208_22, s_207_23, s_206_23, 
s_205_24, s_204_24, s_203_25, s_202_25, s_201_26, s_200_26, 
s_199_27, s_198_27, s_197_28, s_196_28, s_195_29, s_194_29, 
s_193_30, s_192_30, s_191_31, s_190_31, s_189_32, s_188_32, 
s_187_33, s_186_33, s_185_34, s_184_34, s_183_35, s_182_35, 
s_181_36, s_180_36, s_179_37, s_178_37, s_177_38, s_176_38, 
s_175_39, s_174_39, s_173_40, s_172_40, s_171_41, s_170_41, 
s_169_42, s_168_42, s_167_43, s_166_43, s_165_44, s_164_44, 
s_163_45, s_162_45, s_161_46, s_160_46, s_159_47, s_158_47, 
s_157_48, s_156_48, s_155_49, s_154_49, s_153_50, s_152_50, 
s_151_51, s_150_51, s_149_52, s_148_52, s_147_53, s_146_53, 
s_145_54, s_144_54, s_143_55, s_142_55, s_141_56, s_140_56, 
s_139_57, s_138_57, s_137_58, s_136_58, s_135_59, s_134_59, 
s_133_60, s_132_60, s_131_61, s_130_61, s_129_62, s_128_62, 
s_127_62, s_126_62, s_125_62, s_124_62
} = partial_products[(width+2)*(62+1)-1:(width+2)*62];

assign {
 s_255_0,  s_254_0,  s_253_1,  s_252_1,  s_251_2,  s_250_2, 
 s_249_3,  s_248_3,  s_247_4,  s_246_4,  s_245_5,  s_244_5, 
 s_243_6,  s_242_6,  s_241_7,  s_240_7,  s_239_8,  s_238_8, 
 s_237_9,  s_236_9, s_235_10, s_234_10, s_233_11, s_232_11, 
s_231_12, s_230_12, s_229_13, s_228_13, s_227_14, s_226_14, 
s_225_15, s_224_15, s_223_16, s_222_16, s_221_17, s_220_17, 
s_219_18, s_218_18, s_217_19, s_216_19, s_215_20, s_214_20, 
s_213_21, s_212_21, s_211_22, s_210_22, s_209_23, s_208_23, 
s_207_24, s_206_24, s_205_25, s_204_25, s_203_26, s_202_26, 
s_201_27, s_200_27, s_199_28, s_198_28, s_197_29, s_196_29, 
s_195_30, s_194_30, s_193_31, s_192_31, s_191_32, s_190_32, 
s_189_33, s_188_33, s_187_34, s_186_34, s_185_35, s_184_35, 
s_183_36, s_182_36, s_181_37, s_180_37, s_179_38, s_178_38, 
s_177_39, s_176_39, s_175_40, s_174_40, s_173_41, s_172_41, 
s_171_42, s_170_42, s_169_43, s_168_43, s_167_44, s_166_44, 
s_165_45, s_164_45, s_163_46, s_162_46, s_161_47, s_160_47, 
s_159_48, s_158_48, s_157_49, s_156_49, s_155_50, s_154_50, 
s_153_51, s_152_51, s_151_52, s_150_52, s_149_53, s_148_53, 
s_147_54, s_146_54, s_145_55, s_144_55, s_143_56, s_142_56, 
s_141_57, s_140_57, s_139_58, s_138_58, s_137_59, s_136_59, 
s_135_60, s_134_60, s_133_61, s_132_61, s_131_62, s_130_62, 
s_129_63, s_128_63, s_127_63, s_126_63
} = partial_products[(width+2)*(63+1)-1:(width+2)*63];

assign {
 s_255_1,  s_254_1,  s_253_2,  s_252_2,  s_251_3,  s_250_3, 
 s_249_4,  s_248_4,  s_247_5,  s_246_5,  s_245_6,  s_244_6, 
 s_243_7,  s_242_7,  s_241_8,  s_240_8,  s_239_9,  s_238_9, 
s_237_10, s_236_10, s_235_11, s_234_11, s_233_12, s_232_12, 
s_231_13, s_230_13, s_229_14, s_228_14, s_227_15, s_226_15, 
s_225_16, s_224_16, s_223_17, s_222_17, s_221_18, s_220_18, 
s_219_19, s_218_19, s_217_20, s_216_20, s_215_21, s_214_21, 
s_213_22, s_212_22, s_211_23, s_210_23, s_209_24, s_208_24, 
s_207_25, s_206_25, s_205_26, s_204_26, s_203_27, s_202_27, 
s_201_28, s_200_28, s_199_29, s_198_29, s_197_30, s_196_30, 
s_195_31, s_194_31, s_193_32, s_192_32, s_191_33, s_190_33, 
s_189_34, s_188_34, s_187_35, s_186_35, s_185_36, s_184_36, 
s_183_37, s_182_37, s_181_38, s_180_38, s_179_39, s_178_39, 
s_177_40, s_176_40, s_175_41, s_174_41, s_173_42, s_172_42, 
s_171_43, s_170_43, s_169_44, s_168_44, s_167_45, s_166_45, 
s_165_46, s_164_46, s_163_47, s_162_47, s_161_48, s_160_48, 
s_159_49, s_158_49, s_157_50, s_156_50, s_155_51, s_154_51, 
s_153_52, s_152_52, s_151_53, s_150_53, s_149_54, s_148_54, 
s_147_55, s_146_55, s_145_56, s_144_56, s_143_57, s_142_57, 
s_141_58, s_140_58, s_139_59, s_138_59, s_137_60, s_136_60, 
s_135_61, s_134_61, s_133_62, s_132_62, s_131_63, s_130_63, 
s_129_64, s_128_64
} = partial_products[(width+2)*(width/2+1)-1:(width+2)*width/2+2];

/* u0_1 Output nets */
wire t_0,      t_1;
/* u1_2 Output nets */
wire t_2,      t_3;
/* u0_3 Output nets */
wire t_4,      t_5;
/* u1_4 Output nets */
wire t_6,      t_7;
/* u1_5 Output nets */
wire t_8,      t_9;
/* u2_6 Output nets */
wire t_10,     t_11,     t_12;
/* u2_7 Output nets */
wire t_13,     t_14,     t_15;
/* u2_8 Output nets */
wire t_16,     t_17,     t_18;
/* u0_9 Output nets */
wire t_19,     t_20;
/* u2_10 Output nets */
wire t_21,     t_22,     t_23;
/* u2_11 Output nets */
wire t_24,     t_25,     t_26;
/* u1_12 Output nets */
wire t_27,     t_28;
/* u2_13 Output nets */
wire t_29,     t_30,     t_31;
/* u0_14 Output nets */
wire t_32,     t_33;
/* u2_15 Output nets */
wire t_34,     t_35,     t_36;
/* u1_16 Output nets */
wire t_37,     t_38;
/* u2_17 Output nets */
wire t_39,     t_40,     t_41;
/* u1_18 Output nets */
wire t_42,     t_43;
/* u2_19 Output nets */
wire t_44,     t_45,     t_46;
/* u2_20 Output nets */
wire t_47,     t_48,     t_49;
/* u2_21 Output nets */
wire t_50,     t_51,     t_52;
/* u2_22 Output nets */
wire t_53,     t_54,     t_55;
/* u2_23 Output nets */
wire t_56,     t_57,     t_58;
/* u2_24 Output nets */
wire t_59,     t_60,     t_61;
/* u0_25 Output nets */
wire t_62,     t_63;
/* u2_26 Output nets */
wire t_64,     t_65,     t_66;
/* u2_27 Output nets */
wire t_67,     t_68,     t_69;
/* u2_28 Output nets */
wire t_70,     t_71,     t_72;
/* u2_29 Output nets */
wire t_73,     t_74,     t_75;
/* u1_30 Output nets */
wire t_76,     t_77;
/* u2_31 Output nets */
wire t_78,     t_79,     t_80;
/* u2_32 Output nets */
wire t_81,     t_82,     t_83;
/* u0_33 Output nets */
wire t_84,     t_85;
/* u2_34 Output nets */
wire t_86,     t_87,     t_88;
/* u2_35 Output nets */
wire t_89,     t_90,     t_91;
/* u1_36 Output nets */
wire t_92,     t_93;
/* u2_37 Output nets */
wire t_94,     t_95,     t_96;
/* u2_38 Output nets */
wire t_97,     t_98,     t_99;
/* u1_39 Output nets */
wire t_100,    t_101;
/* u2_40 Output nets */
wire t_102,    t_103,    t_104;
/* u2_41 Output nets */
wire t_105,    t_106,    t_107;
/* u2_42 Output nets */
wire t_108,    t_109,    t_110;
/* u2_43 Output nets */
wire t_111,    t_112,    t_113;
/* u2_44 Output nets */
wire t_114,    t_115,    t_116;
/* u2_45 Output nets */
wire t_117,    t_118,    t_119;
/* u2_46 Output nets */
wire t_120,    t_121,    t_122;
/* u2_47 Output nets */
wire t_123,    t_124,    t_125;
/* u2_48 Output nets */
wire t_126,    t_127,    t_128;
/* u0_49 Output nets */
wire t_129,    t_130;
/* u2_50 Output nets */
wire t_131,    t_132,    t_133;
/* u2_51 Output nets */
wire t_134,    t_135,    t_136;
/* u2_52 Output nets */
wire t_137,    t_138,    t_139;
/* u2_53 Output nets */
wire t_140,    t_141,    t_142;
/* u2_54 Output nets */
wire t_143,    t_144,    t_145;
/* u2_55 Output nets */
wire t_146,    t_147,    t_148;
/* u1_56 Output nets */
wire t_149,    t_150;
/* u2_57 Output nets */
wire t_151,    t_152,    t_153;
/* u2_58 Output nets */
wire t_154,    t_155,    t_156;
/* u2_59 Output nets */
wire t_157,    t_158,    t_159;
/* u0_60 Output nets */
wire t_160,    t_161;
/* u2_61 Output nets */
wire t_162,    t_163,    t_164;
/* u2_62 Output nets */
wire t_165,    t_166,    t_167;
/* u2_63 Output nets */
wire t_168,    t_169,    t_170;
/* u1_64 Output nets */
wire t_171,    t_172;
/* u2_65 Output nets */
wire t_173,    t_174,    t_175;
/* u2_66 Output nets */
wire t_176,    t_177,    t_178;
/* u2_67 Output nets */
wire t_179,    t_180,    t_181;
/* u1_68 Output nets */
wire t_182,    t_183;
/* u2_69 Output nets */
wire t_184,    t_185,    t_186;
/* u2_70 Output nets */
wire t_187,    t_188,    t_189;
/* u2_71 Output nets */
wire t_190,    t_191,    t_192;
/* u2_72 Output nets */
wire t_193,    t_194,    t_195;
/* u2_73 Output nets */
wire t_196,    t_197,    t_198;
/* u2_74 Output nets */
wire t_199,    t_200,    t_201;
/* u2_75 Output nets */
wire t_202,    t_203,    t_204;
/* u2_76 Output nets */
wire t_205,    t_206,    t_207;
/* u2_77 Output nets */
wire t_208,    t_209,    t_210;
/* u2_78 Output nets */
wire t_211,    t_212,    t_213;
/* u2_79 Output nets */
wire t_214,    t_215,    t_216;
/* u2_80 Output nets */
wire t_217,    t_218,    t_219;
/* u0_81 Output nets */
wire t_220,    t_221;
/* u2_82 Output nets */
wire t_222,    t_223,    t_224;
/* u2_83 Output nets */
wire t_225,    t_226,    t_227;
/* u2_84 Output nets */
wire t_228,    t_229,    t_230;
/* u2_85 Output nets */
wire t_231,    t_232,    t_233;
/* u2_86 Output nets */
wire t_234,    t_235,    t_236;
/* u2_87 Output nets */
wire t_237,    t_238,    t_239;
/* u2_88 Output nets */
wire t_240,    t_241,    t_242;
/* u2_89 Output nets */
wire t_243,    t_244,    t_245;
/* u1_90 Output nets */
wire t_246,    t_247;
/* u2_91 Output nets */
wire t_248,    t_249,    t_250;
/* u2_92 Output nets */
wire t_251,    t_252,    t_253;
/* u2_93 Output nets */
wire t_254,    t_255,    t_256;
/* u2_94 Output nets */
wire t_257,    t_258,    t_259;
/* u0_95 Output nets */
wire t_260,    t_261;
/* u2_96 Output nets */
wire t_262,    t_263,    t_264;
/* u2_97 Output nets */
wire t_265,    t_266,    t_267;
/* u2_98 Output nets */
wire t_268,    t_269,    t_270;
/* u2_99 Output nets */
wire t_271,    t_272,    t_273;
/* u1_100 Output nets */
wire t_274,    t_275;
/* u2_101 Output nets */
wire t_276,    t_277,    t_278;
/* u2_102 Output nets */
wire t_279,    t_280,    t_281;
/* u2_103 Output nets */
wire t_282,    t_283,    t_284;
/* u2_104 Output nets */
wire t_285,    t_286,    t_287;
/* u1_105 Output nets */
wire t_288,    t_289;
/* u2_106 Output nets */
wire t_290,    t_291,    t_292;
/* u2_107 Output nets */
wire t_293,    t_294,    t_295;
/* u2_108 Output nets */
wire t_296,    t_297,    t_298;
/* u2_109 Output nets */
wire t_299,    t_300,    t_301;
/* u2_110 Output nets */
wire t_302,    t_303,    t_304;
/* u2_111 Output nets */
wire t_305,    t_306,    t_307;
/* u2_112 Output nets */
wire t_308,    t_309,    t_310;
/* u2_113 Output nets */
wire t_311,    t_312,    t_313;
/* u2_114 Output nets */
wire t_314,    t_315,    t_316;
/* u2_115 Output nets */
wire t_317,    t_318,    t_319;
/* u2_116 Output nets */
wire t_320,    t_321,    t_322;
/* u2_117 Output nets */
wire t_323,    t_324,    t_325;
/* u2_118 Output nets */
wire t_326,    t_327,    t_328;
/* u2_119 Output nets */
wire t_329,    t_330,    t_331;
/* u2_120 Output nets */
wire t_332,    t_333,    t_334;
/* u0_121 Output nets */
wire t_335,    t_336;
/* u2_122 Output nets */
wire t_337,    t_338,    t_339;
/* u2_123 Output nets */
wire t_340,    t_341,    t_342;
/* u2_124 Output nets */
wire t_343,    t_344,    t_345;
/* u2_125 Output nets */
wire t_346,    t_347,    t_348;
/* u2_126 Output nets */
wire t_349,    t_350,    t_351;
/* u2_127 Output nets */
wire t_352,    t_353,    t_354;
/* u2_128 Output nets */
wire t_355,    t_356,    t_357;
/* u2_129 Output nets */
wire t_358,    t_359,    t_360;
/* u2_130 Output nets */
wire t_361,    t_362,    t_363;
/* u2_131 Output nets */
wire t_364,    t_365,    t_366;
/* u1_132 Output nets */
wire t_367,    t_368;
/* u2_133 Output nets */
wire t_369,    t_370,    t_371;
/* u2_134 Output nets */
wire t_372,    t_373,    t_374;
/* u2_135 Output nets */
wire t_375,    t_376,    t_377;
/* u2_136 Output nets */
wire t_378,    t_379,    t_380;
/* u2_137 Output nets */
wire t_381,    t_382,    t_383;
/* u0_138 Output nets */
wire t_384,    t_385;
/* u2_139 Output nets */
wire t_386,    t_387,    t_388;
/* u2_140 Output nets */
wire t_389,    t_390,    t_391;
/* u2_141 Output nets */
wire t_392,    t_393,    t_394;
/* u2_142 Output nets */
wire t_395,    t_396,    t_397;
/* u2_143 Output nets */
wire t_398,    t_399,    t_400;
/* u1_144 Output nets */
wire t_401,    t_402;
/* u2_145 Output nets */
wire t_403,    t_404,    t_405;
/* u2_146 Output nets */
wire t_406,    t_407,    t_408;
/* u2_147 Output nets */
wire t_409,    t_410,    t_411;
/* u2_148 Output nets */
wire t_412,    t_413,    t_414;
/* u2_149 Output nets */
wire t_415,    t_416,    t_417;
/* u1_150 Output nets */
wire t_418,    t_419;
/* u2_151 Output nets */
wire t_420,    t_421,    t_422;
/* u2_152 Output nets */
wire t_423,    t_424,    t_425;
/* u2_153 Output nets */
wire t_426,    t_427,    t_428;
/* u2_154 Output nets */
wire t_429,    t_430,    t_431;
/* u2_155 Output nets */
wire t_432,    t_433,    t_434;
/* u2_156 Output nets */
wire t_435,    t_436,    t_437;
/* u2_157 Output nets */
wire t_438,    t_439,    t_440;
/* u2_158 Output nets */
wire t_441,    t_442,    t_443;
/* u2_159 Output nets */
wire t_444,    t_445,    t_446;
/* u2_160 Output nets */
wire t_447,    t_448,    t_449;
/* u2_161 Output nets */
wire t_450,    t_451,    t_452;
/* u2_162 Output nets */
wire t_453,    t_454,    t_455;
/* u2_163 Output nets */
wire t_456,    t_457,    t_458;
/* u2_164 Output nets */
wire t_459,    t_460,    t_461;
/* u2_165 Output nets */
wire t_462,    t_463,    t_464;
/* u2_166 Output nets */
wire t_465,    t_466,    t_467;
/* u2_167 Output nets */
wire t_468,    t_469,    t_470;
/* u2_168 Output nets */
wire t_471,    t_472,    t_473;
/* u0_169 Output nets */
wire t_474,    t_475;
/* u2_170 Output nets */
wire t_476,    t_477,    t_478;
/* u2_171 Output nets */
wire t_479,    t_480,    t_481;
/* u2_172 Output nets */
wire t_482,    t_483,    t_484;
/* u2_173 Output nets */
wire t_485,    t_486,    t_487;
/* u2_174 Output nets */
wire t_488,    t_489,    t_490;
/* u2_175 Output nets */
wire t_491,    t_492,    t_493;
/* u2_176 Output nets */
wire t_494,    t_495,    t_496;
/* u2_177 Output nets */
wire t_497,    t_498,    t_499;
/* u2_178 Output nets */
wire t_500,    t_501,    t_502;
/* u2_179 Output nets */
wire t_503,    t_504,    t_505;
/* u2_180 Output nets */
wire t_506,    t_507,    t_508;
/* u2_181 Output nets */
wire t_509,    t_510,    t_511;
/* u1_182 Output nets */
wire t_512,    t_513;
/* u2_183 Output nets */
wire t_514,    t_515,    t_516;
/* u2_184 Output nets */
wire t_517,    t_518,    t_519;
/* u2_185 Output nets */
wire t_520,    t_521,    t_522;
/* u2_186 Output nets */
wire t_523,    t_524,    t_525;
/* u2_187 Output nets */
wire t_526,    t_527,    t_528;
/* u2_188 Output nets */
wire t_529,    t_530,    t_531;
/* u0_189 Output nets */
wire t_532,    t_533;
/* u2_190 Output nets */
wire t_534,    t_535,    t_536;
/* u2_191 Output nets */
wire t_537,    t_538,    t_539;
/* u2_192 Output nets */
wire t_540,    t_541,    t_542;
/* u2_193 Output nets */
wire t_543,    t_544,    t_545;
/* u2_194 Output nets */
wire t_546,    t_547,    t_548;
/* u2_195 Output nets */
wire t_549,    t_550,    t_551;
/* u1_196 Output nets */
wire t_552,    t_553;
/* u2_197 Output nets */
wire t_554,    t_555,    t_556;
/* u2_198 Output nets */
wire t_557,    t_558,    t_559;
/* u2_199 Output nets */
wire t_560,    t_561,    t_562;
/* u2_200 Output nets */
wire t_563,    t_564,    t_565;
/* u2_201 Output nets */
wire t_566,    t_567,    t_568;
/* u2_202 Output nets */
wire t_569,    t_570,    t_571;
/* u1_203 Output nets */
wire t_572,    t_573;
/* u2_204 Output nets */
wire t_574,    t_575,    t_576;
/* u2_205 Output nets */
wire t_577,    t_578,    t_579;
/* u2_206 Output nets */
wire t_580,    t_581,    t_582;
/* u2_207 Output nets */
wire t_583,    t_584,    t_585;
/* u2_208 Output nets */
wire t_586,    t_587,    t_588;
/* u2_209 Output nets */
wire t_589,    t_590,    t_591;
/* u2_210 Output nets */
wire t_592,    t_593,    t_594;
/* u2_211 Output nets */
wire t_595,    t_596,    t_597;
/* u2_212 Output nets */
wire t_598,    t_599,    t_600;
/* u2_213 Output nets */
wire t_601,    t_602,    t_603;
/* u2_214 Output nets */
wire t_604,    t_605,    t_606;
/* u2_215 Output nets */
wire t_607,    t_608,    t_609;
/* u2_216 Output nets */
wire t_610,    t_611,    t_612;
/* u2_217 Output nets */
wire t_613,    t_614,    t_615;
/* u2_218 Output nets */
wire t_616,    t_617,    t_618;
/* u2_219 Output nets */
wire t_619,    t_620,    t_621;
/* u2_220 Output nets */
wire t_622,    t_623,    t_624;
/* u2_221 Output nets */
wire t_625,    t_626,    t_627;
/* u2_222 Output nets */
wire t_628,    t_629,    t_630;
/* u2_223 Output nets */
wire t_631,    t_632,    t_633;
/* u2_224 Output nets */
wire t_634,    t_635,    t_636;
/* u0_225 Output nets */
wire t_637,    t_638;
/* u2_226 Output nets */
wire t_639,    t_640,    t_641;
/* u2_227 Output nets */
wire t_642,    t_643,    t_644;
/* u2_228 Output nets */
wire t_645,    t_646,    t_647;
/* u2_229 Output nets */
wire t_648,    t_649,    t_650;
/* u2_230 Output nets */
wire t_651,    t_652,    t_653;
/* u2_231 Output nets */
wire t_654,    t_655,    t_656;
/* u2_232 Output nets */
wire t_657,    t_658,    t_659;
/* u2_233 Output nets */
wire t_660,    t_661,    t_662;
/* u2_234 Output nets */
wire t_663,    t_664,    t_665;
/* u2_235 Output nets */
wire t_666,    t_667,    t_668;
/* u2_236 Output nets */
wire t_669,    t_670,    t_671;
/* u2_237 Output nets */
wire t_672,    t_673,    t_674;
/* u2_238 Output nets */
wire t_675,    t_676,    t_677;
/* u2_239 Output nets */
wire t_678,    t_679,    t_680;
/* u1_240 Output nets */
wire t_681,    t_682;
/* u2_241 Output nets */
wire t_683,    t_684,    t_685;
/* u2_242 Output nets */
wire t_686,    t_687,    t_688;
/* u2_243 Output nets */
wire t_689,    t_690,    t_691;
/* u2_244 Output nets */
wire t_692,    t_693,    t_694;
/* u2_245 Output nets */
wire t_695,    t_696,    t_697;
/* u2_246 Output nets */
wire t_698,    t_699,    t_700;
/* u2_247 Output nets */
wire t_701,    t_702,    t_703;
/* u0_248 Output nets */
wire t_704,    t_705;
/* u2_249 Output nets */
wire t_706,    t_707,    t_708;
/* u2_250 Output nets */
wire t_709,    t_710,    t_711;
/* u2_251 Output nets */
wire t_712,    t_713,    t_714;
/* u2_252 Output nets */
wire t_715,    t_716,    t_717;
/* u2_253 Output nets */
wire t_718,    t_719,    t_720;
/* u2_254 Output nets */
wire t_721,    t_722,    t_723;
/* u2_255 Output nets */
wire t_724,    t_725,    t_726;
/* u1_256 Output nets */
wire t_727,    t_728;
/* u2_257 Output nets */
wire t_729,    t_730,    t_731;
/* u2_258 Output nets */
wire t_732,    t_733,    t_734;
/* u2_259 Output nets */
wire t_735,    t_736,    t_737;
/* u2_260 Output nets */
wire t_738,    t_739,    t_740;
/* u2_261 Output nets */
wire t_741,    t_742,    t_743;
/* u2_262 Output nets */
wire t_744,    t_745,    t_746;
/* u2_263 Output nets */
wire t_747,    t_748,    t_749;
/* u1_264 Output nets */
wire t_750,    t_751;
/* u2_265 Output nets */
wire t_752,    t_753,    t_754;
/* u2_266 Output nets */
wire t_755,    t_756,    t_757;
/* u2_267 Output nets */
wire t_758,    t_759,    t_760;
/* u2_268 Output nets */
wire t_761,    t_762,    t_763;
/* u2_269 Output nets */
wire t_764,    t_765,    t_766;
/* u2_270 Output nets */
wire t_767,    t_768,    t_769;
/* u2_271 Output nets */
wire t_770,    t_771,    t_772;
/* u2_272 Output nets */
wire t_773,    t_774,    t_775;
/* u2_273 Output nets */
wire t_776,    t_777,    t_778;
/* u2_274 Output nets */
wire t_779,    t_780,    t_781;
/* u2_275 Output nets */
wire t_782,    t_783,    t_784;
/* u2_276 Output nets */
wire t_785,    t_786,    t_787;
/* u2_277 Output nets */
wire t_788,    t_789,    t_790;
/* u2_278 Output nets */
wire t_791,    t_792,    t_793;
/* u2_279 Output nets */
wire t_794,    t_795,    t_796;
/* u2_280 Output nets */
wire t_797,    t_798,    t_799;
/* u2_281 Output nets */
wire t_800,    t_801,    t_802;
/* u2_282 Output nets */
wire t_803,    t_804,    t_805;
/* u2_283 Output nets */
wire t_806,    t_807,    t_808;
/* u2_284 Output nets */
wire t_809,    t_810,    t_811;
/* u2_285 Output nets */
wire t_812,    t_813,    t_814;
/* u2_286 Output nets */
wire t_815,    t_816,    t_817;
/* u2_287 Output nets */
wire t_818,    t_819,    t_820;
/* u2_288 Output nets */
wire t_821,    t_822,    t_823;
/* u0_289 Output nets */
wire t_824,    t_825;
/* u2_290 Output nets */
wire t_826,    t_827,    t_828;
/* u2_291 Output nets */
wire t_829,    t_830,    t_831;
/* u2_292 Output nets */
wire t_832,    t_833,    t_834;
/* u2_293 Output nets */
wire t_835,    t_836,    t_837;
/* u2_294 Output nets */
wire t_838,    t_839,    t_840;
/* u2_295 Output nets */
wire t_841,    t_842,    t_843;
/* u2_296 Output nets */
wire t_844,    t_845,    t_846;
/* u2_297 Output nets */
wire t_847,    t_848,    t_849;
/* u2_298 Output nets */
wire t_850,    t_851,    t_852;
/* u2_299 Output nets */
wire t_853,    t_854,    t_855;
/* u2_300 Output nets */
wire t_856,    t_857,    t_858;
/* u2_301 Output nets */
wire t_859,    t_860,    t_861;
/* u2_302 Output nets */
wire t_862,    t_863,    t_864;
/* u2_303 Output nets */
wire t_865,    t_866,    t_867;
/* u2_304 Output nets */
wire t_868,    t_869,    t_870;
/* u2_305 Output nets */
wire t_871,    t_872,    t_873;
/* u1_306 Output nets */
wire t_874,    t_875;
/* u2_307 Output nets */
wire t_876,    t_877,    t_878;
/* u2_308 Output nets */
wire t_879,    t_880,    t_881;
/* u2_309 Output nets */
wire t_882,    t_883,    t_884;
/* u2_310 Output nets */
wire t_885,    t_886,    t_887;
/* u2_311 Output nets */
wire t_888,    t_889,    t_890;
/* u2_312 Output nets */
wire t_891,    t_892,    t_893;
/* u2_313 Output nets */
wire t_894,    t_895,    t_896;
/* u2_314 Output nets */
wire t_897,    t_898,    t_899;
/* u0_315 Output nets */
wire t_900,    t_901;
/* u2_316 Output nets */
wire t_902,    t_903,    t_904;
/* u2_317 Output nets */
wire t_905,    t_906,    t_907;
/* u2_318 Output nets */
wire t_908,    t_909,    t_910;
/* u2_319 Output nets */
wire t_911,    t_912,    t_913;
/* u2_320 Output nets */
wire t_914,    t_915,    t_916;
/* u2_321 Output nets */
wire t_917,    t_918,    t_919;
/* u2_322 Output nets */
wire t_920,    t_921,    t_922;
/* u2_323 Output nets */
wire t_923,    t_924,    t_925;
/* u1_324 Output nets */
wire t_926,    t_927;
/* u2_325 Output nets */
wire t_928,    t_929,    t_930;
/* u2_326 Output nets */
wire t_931,    t_932,    t_933;
/* u2_327 Output nets */
wire t_934,    t_935,    t_936;
/* u2_328 Output nets */
wire t_937,    t_938,    t_939;
/* u2_329 Output nets */
wire t_940,    t_941,    t_942;
/* u2_330 Output nets */
wire t_943,    t_944,    t_945;
/* u2_331 Output nets */
wire t_946,    t_947,    t_948;
/* u2_332 Output nets */
wire t_949,    t_950,    t_951;
/* u1_333 Output nets */
wire t_952,    t_953;
/* u2_334 Output nets */
wire t_954,    t_955,    t_956;
/* u2_335 Output nets */
wire t_957,    t_958,    t_959;
/* u2_336 Output nets */
wire t_960,    t_961,    t_962;
/* u2_337 Output nets */
wire t_963,    t_964,    t_965;
/* u2_338 Output nets */
wire t_966,    t_967,    t_968;
/* u2_339 Output nets */
wire t_969,    t_970,    t_971;
/* u2_340 Output nets */
wire t_972,    t_973,    t_974;
/* u2_341 Output nets */
wire t_975,    t_976,    t_977;
/* u2_342 Output nets */
wire t_978,    t_979,    t_980;
/* u2_343 Output nets */
wire t_981,    t_982,    t_983;
/* u2_344 Output nets */
wire t_984,    t_985,    t_986;
/* u2_345 Output nets */
wire t_987,    t_988,    t_989;
/* u2_346 Output nets */
wire t_990,    t_991,    t_992;
/* u2_347 Output nets */
wire t_993,    t_994,    t_995;
/* u2_348 Output nets */
wire t_996,    t_997,    t_998;
/* u2_349 Output nets */
wire t_999,   t_1000,   t_1001;
/* u2_350 Output nets */
wire t_1002,   t_1003,   t_1004;
/* u2_351 Output nets */
wire t_1005,   t_1006,   t_1007;
/* u2_352 Output nets */
wire t_1008,   t_1009,   t_1010;
/* u2_353 Output nets */
wire t_1011,   t_1012,   t_1013;
/* u2_354 Output nets */
wire t_1014,   t_1015,   t_1016;
/* u2_355 Output nets */
wire t_1017,   t_1018,   t_1019;
/* u2_356 Output nets */
wire t_1020,   t_1021,   t_1022;
/* u2_357 Output nets */
wire t_1023,   t_1024,   t_1025;
/* u2_358 Output nets */
wire t_1026,   t_1027,   t_1028;
/* u2_359 Output nets */
wire t_1029,   t_1030,   t_1031;
/* u2_360 Output nets */
wire t_1032,   t_1033,   t_1034;
/* u0_361 Output nets */
wire t_1035,   t_1036;
/* u2_362 Output nets */
wire t_1037,   t_1038,   t_1039;
/* u2_363 Output nets */
wire t_1040,   t_1041,   t_1042;
/* u2_364 Output nets */
wire t_1043,   t_1044,   t_1045;
/* u2_365 Output nets */
wire t_1046,   t_1047,   t_1048;
/* u2_366 Output nets */
wire t_1049,   t_1050,   t_1051;
/* u2_367 Output nets */
wire t_1052,   t_1053,   t_1054;
/* u2_368 Output nets */
wire t_1055,   t_1056,   t_1057;
/* u2_369 Output nets */
wire t_1058,   t_1059,   t_1060;
/* u2_370 Output nets */
wire t_1061,   t_1062,   t_1063;
/* u2_371 Output nets */
wire t_1064,   t_1065,   t_1066;
/* u2_372 Output nets */
wire t_1067,   t_1068,   t_1069;
/* u2_373 Output nets */
wire t_1070,   t_1071,   t_1072;
/* u2_374 Output nets */
wire t_1073,   t_1074,   t_1075;
/* u2_375 Output nets */
wire t_1076,   t_1077,   t_1078;
/* u2_376 Output nets */
wire t_1079,   t_1080,   t_1081;
/* u2_377 Output nets */
wire t_1082,   t_1083,   t_1084;
/* u2_378 Output nets */
wire t_1085,   t_1086,   t_1087;
/* u2_379 Output nets */
wire t_1088,   t_1089,   t_1090;
/* u1_380 Output nets */
wire t_1091,   t_1092;
/* u2_381 Output nets */
wire t_1093,   t_1094,   t_1095;
/* u2_382 Output nets */
wire t_1096,   t_1097,   t_1098;
/* u2_383 Output nets */
wire t_1099,   t_1100,   t_1101;
/* u2_384 Output nets */
wire t_1102,   t_1103,   t_1104;
/* u2_385 Output nets */
wire t_1105,   t_1106,   t_1107;
/* u2_386 Output nets */
wire t_1108,   t_1109,   t_1110;
/* u2_387 Output nets */
wire t_1111,   t_1112,   t_1113;
/* u2_388 Output nets */
wire t_1114,   t_1115,   t_1116;
/* u2_389 Output nets */
wire t_1117,   t_1118,   t_1119;
/* u0_390 Output nets */
wire t_1120,   t_1121;
/* u2_391 Output nets */
wire t_1122,   t_1123,   t_1124;
/* u2_392 Output nets */
wire t_1125,   t_1126,   t_1127;
/* u2_393 Output nets */
wire t_1128,   t_1129,   t_1130;
/* u2_394 Output nets */
wire t_1131,   t_1132,   t_1133;
/* u2_395 Output nets */
wire t_1134,   t_1135,   t_1136;
/* u2_396 Output nets */
wire t_1137,   t_1138,   t_1139;
/* u2_397 Output nets */
wire t_1140,   t_1141,   t_1142;
/* u2_398 Output nets */
wire t_1143,   t_1144,   t_1145;
/* u2_399 Output nets */
wire t_1146,   t_1147,   t_1148;
/* u1_400 Output nets */
wire t_1149,   t_1150;
/* u2_401 Output nets */
wire t_1151,   t_1152,   t_1153;
/* u2_402 Output nets */
wire t_1154,   t_1155,   t_1156;
/* u2_403 Output nets */
wire t_1157,   t_1158,   t_1159;
/* u2_404 Output nets */
wire t_1160,   t_1161,   t_1162;
/* u2_405 Output nets */
wire t_1163,   t_1164,   t_1165;
/* u2_406 Output nets */
wire t_1166,   t_1167,   t_1168;
/* u2_407 Output nets */
wire t_1169,   t_1170,   t_1171;
/* u2_408 Output nets */
wire t_1172,   t_1173,   t_1174;
/* u2_409 Output nets */
wire t_1175,   t_1176,   t_1177;
/* u1_410 Output nets */
wire t_1178,   t_1179;
/* u2_411 Output nets */
wire t_1180,   t_1181,   t_1182;
/* u2_412 Output nets */
wire t_1183,   t_1184,   t_1185;
/* u2_413 Output nets */
wire t_1186,   t_1187,   t_1188;
/* u2_414 Output nets */
wire t_1189,   t_1190,   t_1191;
/* u2_415 Output nets */
wire t_1192,   t_1193,   t_1194;
/* u2_416 Output nets */
wire t_1195,   t_1196,   t_1197;
/* u2_417 Output nets */
wire t_1198,   t_1199,   t_1200;
/* u2_418 Output nets */
wire t_1201,   t_1202,   t_1203;
/* u2_419 Output nets */
wire t_1204,   t_1205,   t_1206;
/* u2_420 Output nets */
wire t_1207,   t_1208,   t_1209;
/* u2_421 Output nets */
wire t_1210,   t_1211,   t_1212;
/* u2_422 Output nets */
wire t_1213,   t_1214,   t_1215;
/* u2_423 Output nets */
wire t_1216,   t_1217,   t_1218;
/* u2_424 Output nets */
wire t_1219,   t_1220,   t_1221;
/* u2_425 Output nets */
wire t_1222,   t_1223,   t_1224;
/* u2_426 Output nets */
wire t_1225,   t_1226,   t_1227;
/* u2_427 Output nets */
wire t_1228,   t_1229,   t_1230;
/* u2_428 Output nets */
wire t_1231,   t_1232,   t_1233;
/* u2_429 Output nets */
wire t_1234,   t_1235,   t_1236;
/* u2_430 Output nets */
wire t_1237,   t_1238,   t_1239;
/* u2_431 Output nets */
wire t_1240,   t_1241,   t_1242;
/* u2_432 Output nets */
wire t_1243,   t_1244,   t_1245;
/* u2_433 Output nets */
wire t_1246,   t_1247,   t_1248;
/* u2_434 Output nets */
wire t_1249,   t_1250,   t_1251;
/* u2_435 Output nets */
wire t_1252,   t_1253,   t_1254;
/* u2_436 Output nets */
wire t_1255,   t_1256,   t_1257;
/* u2_437 Output nets */
wire t_1258,   t_1259,   t_1260;
/* u2_438 Output nets */
wire t_1261,   t_1262,   t_1263;
/* u2_439 Output nets */
wire t_1264,   t_1265,   t_1266;
/* u2_440 Output nets */
wire t_1267,   t_1268,   t_1269;
/* u0_441 Output nets */
wire t_1270,   t_1271;
/* u2_442 Output nets */
wire t_1272,   t_1273,   t_1274;
/* u2_443 Output nets */
wire t_1275,   t_1276,   t_1277;
/* u2_444 Output nets */
wire t_1278,   t_1279,   t_1280;
/* u2_445 Output nets */
wire t_1281,   t_1282,   t_1283;
/* u2_446 Output nets */
wire t_1284,   t_1285,   t_1286;
/* u2_447 Output nets */
wire t_1287,   t_1288,   t_1289;
/* u2_448 Output nets */
wire t_1290,   t_1291,   t_1292;
/* u2_449 Output nets */
wire t_1293,   t_1294,   t_1295;
/* u2_450 Output nets */
wire t_1296,   t_1297,   t_1298;
/* u2_451 Output nets */
wire t_1299,   t_1300,   t_1301;
/* u2_452 Output nets */
wire t_1302,   t_1303,   t_1304;
/* u2_453 Output nets */
wire t_1305,   t_1306,   t_1307;
/* u2_454 Output nets */
wire t_1308,   t_1309,   t_1310;
/* u2_455 Output nets */
wire t_1311,   t_1312,   t_1313;
/* u2_456 Output nets */
wire t_1314,   t_1315,   t_1316;
/* u2_457 Output nets */
wire t_1317,   t_1318,   t_1319;
/* u2_458 Output nets */
wire t_1320,   t_1321,   t_1322;
/* u2_459 Output nets */
wire t_1323,   t_1324,   t_1325;
/* u2_460 Output nets */
wire t_1326,   t_1327,   t_1328;
/* u2_461 Output nets */
wire t_1329,   t_1330,   t_1331;
/* u1_462 Output nets */
wire t_1332,   t_1333;
/* u2_463 Output nets */
wire t_1334,   t_1335,   t_1336;
/* u2_464 Output nets */
wire t_1337,   t_1338,   t_1339;
/* u2_465 Output nets */
wire t_1340,   t_1341,   t_1342;
/* u2_466 Output nets */
wire t_1343,   t_1344,   t_1345;
/* u2_467 Output nets */
wire t_1346,   t_1347,   t_1348;
/* u2_468 Output nets */
wire t_1349,   t_1350,   t_1351;
/* u2_469 Output nets */
wire t_1352,   t_1353,   t_1354;
/* u2_470 Output nets */
wire t_1355,   t_1356,   t_1357;
/* u2_471 Output nets */
wire t_1358,   t_1359,   t_1360;
/* u2_472 Output nets */
wire t_1361,   t_1362,   t_1363;
/* u0_473 Output nets */
wire t_1364,   t_1365;
/* u2_474 Output nets */
wire t_1366,   t_1367,   t_1368;
/* u2_475 Output nets */
wire t_1369,   t_1370,   t_1371;
/* u2_476 Output nets */
wire t_1372,   t_1373,   t_1374;
/* u2_477 Output nets */
wire t_1375,   t_1376,   t_1377;
/* u2_478 Output nets */
wire t_1378,   t_1379,   t_1380;
/* u2_479 Output nets */
wire t_1381,   t_1382,   t_1383;
/* u2_480 Output nets */
wire t_1384,   t_1385,   t_1386;
/* u2_481 Output nets */
wire t_1387,   t_1388,   t_1389;
/* u2_482 Output nets */
wire t_1390,   t_1391,   t_1392;
/* u2_483 Output nets */
wire t_1393,   t_1394,   t_1395;
/* u1_484 Output nets */
wire t_1396,   t_1397;
/* u2_485 Output nets */
wire t_1398,   t_1399,   t_1400;
/* u2_486 Output nets */
wire t_1401,   t_1402,   t_1403;
/* u2_487 Output nets */
wire t_1404,   t_1405,   t_1406;
/* u2_488 Output nets */
wire t_1407,   t_1408,   t_1409;
/* u2_489 Output nets */
wire t_1410,   t_1411,   t_1412;
/* u2_490 Output nets */
wire t_1413,   t_1414,   t_1415;
/* u2_491 Output nets */
wire t_1416,   t_1417,   t_1418;
/* u2_492 Output nets */
wire t_1419,   t_1420,   t_1421;
/* u2_493 Output nets */
wire t_1422,   t_1423,   t_1424;
/* u2_494 Output nets */
wire t_1425,   t_1426,   t_1427;
/* u1_495 Output nets */
wire t_1428,   t_1429;
/* u2_496 Output nets */
wire t_1430,   t_1431,   t_1432;
/* u2_497 Output nets */
wire t_1433,   t_1434,   t_1435;
/* u2_498 Output nets */
wire t_1436,   t_1437,   t_1438;
/* u2_499 Output nets */
wire t_1439,   t_1440,   t_1441;
/* u2_500 Output nets */
wire t_1442,   t_1443,   t_1444;
/* u2_501 Output nets */
wire t_1445,   t_1446,   t_1447;
/* u2_502 Output nets */
wire t_1448,   t_1449,   t_1450;
/* u2_503 Output nets */
wire t_1451,   t_1452,   t_1453;
/* u2_504 Output nets */
wire t_1454,   t_1455,   t_1456;
/* u2_505 Output nets */
wire t_1457,   t_1458,   t_1459;
/* u2_506 Output nets */
wire t_1460,   t_1461,   t_1462;
/* u2_507 Output nets */
wire t_1463,   t_1464,   t_1465;
/* u2_508 Output nets */
wire t_1466,   t_1467,   t_1468;
/* u2_509 Output nets */
wire t_1469,   t_1470,   t_1471;
/* u2_510 Output nets */
wire t_1472,   t_1473,   t_1474;
/* u2_511 Output nets */
wire t_1475,   t_1476,   t_1477;
/* u2_512 Output nets */
wire t_1478,   t_1479,   t_1480;
/* u2_513 Output nets */
wire t_1481,   t_1482,   t_1483;
/* u2_514 Output nets */
wire t_1484,   t_1485,   t_1486;
/* u2_515 Output nets */
wire t_1487,   t_1488,   t_1489;
/* u2_516 Output nets */
wire t_1490,   t_1491,   t_1492;
/* u2_517 Output nets */
wire t_1493,   t_1494,   t_1495;
/* u2_518 Output nets */
wire t_1496,   t_1497,   t_1498;
/* u2_519 Output nets */
wire t_1499,   t_1500,   t_1501;
/* u2_520 Output nets */
wire t_1502,   t_1503,   t_1504;
/* u2_521 Output nets */
wire t_1505,   t_1506,   t_1507;
/* u2_522 Output nets */
wire t_1508,   t_1509,   t_1510;
/* u2_523 Output nets */
wire t_1511,   t_1512,   t_1513;
/* u2_524 Output nets */
wire t_1514,   t_1515,   t_1516;
/* u2_525 Output nets */
wire t_1517,   t_1518,   t_1519;
/* u2_526 Output nets */
wire t_1520,   t_1521,   t_1522;
/* u2_527 Output nets */
wire t_1523,   t_1524,   t_1525;
/* u2_528 Output nets */
wire t_1526,   t_1527,   t_1528;
/* u0_529 Output nets */
wire t_1529,   t_1530;
/* u2_530 Output nets */
wire t_1531,   t_1532,   t_1533;
/* u2_531 Output nets */
wire t_1534,   t_1535,   t_1536;
/* u2_532 Output nets */
wire t_1537,   t_1538,   t_1539;
/* u2_533 Output nets */
wire t_1540,   t_1541,   t_1542;
/* u2_534 Output nets */
wire t_1543,   t_1544,   t_1545;
/* u2_535 Output nets */
wire t_1546,   t_1547,   t_1548;
/* u2_536 Output nets */
wire t_1549,   t_1550,   t_1551;
/* u2_537 Output nets */
wire t_1552,   t_1553,   t_1554;
/* u2_538 Output nets */
wire t_1555,   t_1556,   t_1557;
/* u2_539 Output nets */
wire t_1558,   t_1559,   t_1560;
/* u2_540 Output nets */
wire t_1561,   t_1562,   t_1563;
/* u2_541 Output nets */
wire t_1564,   t_1565,   t_1566;
/* u2_542 Output nets */
wire t_1567,   t_1568,   t_1569;
/* u2_543 Output nets */
wire t_1570,   t_1571,   t_1572;
/* u2_544 Output nets */
wire t_1573,   t_1574,   t_1575;
/* u2_545 Output nets */
wire t_1576,   t_1577,   t_1578;
/* u2_546 Output nets */
wire t_1579,   t_1580,   t_1581;
/* u2_547 Output nets */
wire t_1582,   t_1583,   t_1584;
/* u2_548 Output nets */
wire t_1585,   t_1586,   t_1587;
/* u2_549 Output nets */
wire t_1588,   t_1589,   t_1590;
/* u2_550 Output nets */
wire t_1591,   t_1592,   t_1593;
/* u2_551 Output nets */
wire t_1594,   t_1595,   t_1596;
/* u1_552 Output nets */
wire t_1597,   t_1598;
/* u2_553 Output nets */
wire t_1599,   t_1600,   t_1601;
/* u2_554 Output nets */
wire t_1602,   t_1603,   t_1604;
/* u2_555 Output nets */
wire t_1605,   t_1606,   t_1607;
/* u2_556 Output nets */
wire t_1608,   t_1609,   t_1610;
/* u2_557 Output nets */
wire t_1611,   t_1612,   t_1613;
/* u2_558 Output nets */
wire t_1614,   t_1615,   t_1616;
/* u2_559 Output nets */
wire t_1617,   t_1618,   t_1619;
/* u2_560 Output nets */
wire t_1620,   t_1621,   t_1622;
/* u2_561 Output nets */
wire t_1623,   t_1624,   t_1625;
/* u2_562 Output nets */
wire t_1626,   t_1627,   t_1628;
/* u2_563 Output nets */
wire t_1629,   t_1630,   t_1631;
/* u0_564 Output nets */
wire t_1632,   t_1633;
/* u2_565 Output nets */
wire t_1634,   t_1635,   t_1636;
/* u2_566 Output nets */
wire t_1637,   t_1638,   t_1639;
/* u2_567 Output nets */
wire t_1640,   t_1641,   t_1642;
/* u2_568 Output nets */
wire t_1643,   t_1644,   t_1645;
/* u2_569 Output nets */
wire t_1646,   t_1647,   t_1648;
/* u2_570 Output nets */
wire t_1649,   t_1650,   t_1651;
/* u2_571 Output nets */
wire t_1652,   t_1653,   t_1654;
/* u2_572 Output nets */
wire t_1655,   t_1656,   t_1657;
/* u2_573 Output nets */
wire t_1658,   t_1659,   t_1660;
/* u2_574 Output nets */
wire t_1661,   t_1662,   t_1663;
/* u2_575 Output nets */
wire t_1664,   t_1665,   t_1666;
/* u1_576 Output nets */
wire t_1667,   t_1668;
/* u2_577 Output nets */
wire t_1669,   t_1670,   t_1671;
/* u2_578 Output nets */
wire t_1672,   t_1673,   t_1674;
/* u2_579 Output nets */
wire t_1675,   t_1676,   t_1677;
/* u2_580 Output nets */
wire t_1678,   t_1679,   t_1680;
/* u2_581 Output nets */
wire t_1681,   t_1682,   t_1683;
/* u2_582 Output nets */
wire t_1684,   t_1685,   t_1686;
/* u2_583 Output nets */
wire t_1687,   t_1688,   t_1689;
/* u2_584 Output nets */
wire t_1690,   t_1691,   t_1692;
/* u2_585 Output nets */
wire t_1693,   t_1694,   t_1695;
/* u2_586 Output nets */
wire t_1696,   t_1697,   t_1698;
/* u2_587 Output nets */
wire t_1699,   t_1700,   t_1701;
/* u1_588 Output nets */
wire t_1702,   t_1703;
/* u2_589 Output nets */
wire t_1704,   t_1705,   t_1706;
/* u2_590 Output nets */
wire t_1707,   t_1708,   t_1709;
/* u2_591 Output nets */
wire t_1710,   t_1711,   t_1712;
/* u2_592 Output nets */
wire t_1713,   t_1714,   t_1715;
/* u2_593 Output nets */
wire t_1716,   t_1717,   t_1718;
/* u2_594 Output nets */
wire t_1719,   t_1720,   t_1721;
/* u2_595 Output nets */
wire t_1722,   t_1723,   t_1724;
/* u2_596 Output nets */
wire t_1725,   t_1726,   t_1727;
/* u2_597 Output nets */
wire t_1728,   t_1729,   t_1730;
/* u2_598 Output nets */
wire t_1731,   t_1732,   t_1733;
/* u2_599 Output nets */
wire t_1734,   t_1735,   t_1736;
/* u2_600 Output nets */
wire t_1737,   t_1738,   t_1739;
/* u2_601 Output nets */
wire t_1740,   t_1741,   t_1742;
/* u2_602 Output nets */
wire t_1743,   t_1744,   t_1745;
/* u2_603 Output nets */
wire t_1746,   t_1747,   t_1748;
/* u2_604 Output nets */
wire t_1749,   t_1750,   t_1751;
/* u2_605 Output nets */
wire t_1752,   t_1753,   t_1754;
/* u2_606 Output nets */
wire t_1755,   t_1756,   t_1757;
/* u2_607 Output nets */
wire t_1758,   t_1759,   t_1760;
/* u2_608 Output nets */
wire t_1761,   t_1762,   t_1763;
/* u2_609 Output nets */
wire t_1764,   t_1765,   t_1766;
/* u2_610 Output nets */
wire t_1767,   t_1768,   t_1769;
/* u2_611 Output nets */
wire t_1770,   t_1771,   t_1772;
/* u2_612 Output nets */
wire t_1773,   t_1774,   t_1775;
/* u2_613 Output nets */
wire t_1776,   t_1777,   t_1778;
/* u2_614 Output nets */
wire t_1779,   t_1780,   t_1781;
/* u2_615 Output nets */
wire t_1782,   t_1783,   t_1784;
/* u2_616 Output nets */
wire t_1785,   t_1786,   t_1787;
/* u2_617 Output nets */
wire t_1788,   t_1789,   t_1790;
/* u2_618 Output nets */
wire t_1791,   t_1792,   t_1793;
/* u2_619 Output nets */
wire t_1794,   t_1795,   t_1796;
/* u2_620 Output nets */
wire t_1797,   t_1798,   t_1799;
/* u2_621 Output nets */
wire t_1800,   t_1801,   t_1802;
/* u2_622 Output nets */
wire t_1803,   t_1804,   t_1805;
/* u2_623 Output nets */
wire t_1806,   t_1807,   t_1808;
/* u2_624 Output nets */
wire t_1809,   t_1810,   t_1811;
/* u0_625 Output nets */
wire t_1812,   t_1813;
/* u2_626 Output nets */
wire t_1814,   t_1815,   t_1816;
/* u2_627 Output nets */
wire t_1817,   t_1818,   t_1819;
/* u2_628 Output nets */
wire t_1820,   t_1821,   t_1822;
/* u2_629 Output nets */
wire t_1823,   t_1824,   t_1825;
/* u2_630 Output nets */
wire t_1826,   t_1827,   t_1828;
/* u2_631 Output nets */
wire t_1829,   t_1830,   t_1831;
/* u2_632 Output nets */
wire t_1832,   t_1833,   t_1834;
/* u2_633 Output nets */
wire t_1835,   t_1836,   t_1837;
/* u2_634 Output nets */
wire t_1838,   t_1839,   t_1840;
/* u2_635 Output nets */
wire t_1841,   t_1842,   t_1843;
/* u2_636 Output nets */
wire t_1844,   t_1845,   t_1846;
/* u2_637 Output nets */
wire t_1847,   t_1848,   t_1849;
/* u2_638 Output nets */
wire t_1850,   t_1851,   t_1852;
/* u2_639 Output nets */
wire t_1853,   t_1854,   t_1855;
/* u2_640 Output nets */
wire t_1856,   t_1857,   t_1858;
/* u2_641 Output nets */
wire t_1859,   t_1860,   t_1861;
/* u2_642 Output nets */
wire t_1862,   t_1863,   t_1864;
/* u2_643 Output nets */
wire t_1865,   t_1866,   t_1867;
/* u2_644 Output nets */
wire t_1868,   t_1869,   t_1870;
/* u2_645 Output nets */
wire t_1871,   t_1872,   t_1873;
/* u2_646 Output nets */
wire t_1874,   t_1875,   t_1876;
/* u2_647 Output nets */
wire t_1877,   t_1878,   t_1879;
/* u2_648 Output nets */
wire t_1880,   t_1881,   t_1882;
/* u2_649 Output nets */
wire t_1883,   t_1884,   t_1885;
/* u1_650 Output nets */
wire t_1886,   t_1887;
/* u2_651 Output nets */
wire t_1888,   t_1889,   t_1890;
/* u2_652 Output nets */
wire t_1891,   t_1892,   t_1893;
/* u2_653 Output nets */
wire t_1894,   t_1895,   t_1896;
/* u2_654 Output nets */
wire t_1897,   t_1898,   t_1899;
/* u2_655 Output nets */
wire t_1900,   t_1901,   t_1902;
/* u2_656 Output nets */
wire t_1903,   t_1904,   t_1905;
/* u2_657 Output nets */
wire t_1906,   t_1907,   t_1908;
/* u2_658 Output nets */
wire t_1909,   t_1910,   t_1911;
/* u2_659 Output nets */
wire t_1912,   t_1913,   t_1914;
/* u2_660 Output nets */
wire t_1915,   t_1916,   t_1917;
/* u2_661 Output nets */
wire t_1918,   t_1919,   t_1920;
/* u2_662 Output nets */
wire t_1921,   t_1922,   t_1923;
/* u0_663 Output nets */
wire t_1924,   t_1925;
/* u2_664 Output nets */
wire t_1926,   t_1927,   t_1928;
/* u2_665 Output nets */
wire t_1929,   t_1930,   t_1931;
/* u2_666 Output nets */
wire t_1932,   t_1933,   t_1934;
/* u2_667 Output nets */
wire t_1935,   t_1936,   t_1937;
/* u2_668 Output nets */
wire t_1938,   t_1939,   t_1940;
/* u2_669 Output nets */
wire t_1941,   t_1942,   t_1943;
/* u2_670 Output nets */
wire t_1944,   t_1945,   t_1946;
/* u2_671 Output nets */
wire t_1947,   t_1948,   t_1949;
/* u2_672 Output nets */
wire t_1950,   t_1951,   t_1952;
/* u2_673 Output nets */
wire t_1953,   t_1954,   t_1955;
/* u2_674 Output nets */
wire t_1956,   t_1957,   t_1958;
/* u2_675 Output nets */
wire t_1959,   t_1960,   t_1961;
/* u1_676 Output nets */
wire t_1962,   t_1963;
/* u2_677 Output nets */
wire t_1964,   t_1965,   t_1966;
/* u2_678 Output nets */
wire t_1967,   t_1968,   t_1969;
/* u2_679 Output nets */
wire t_1970,   t_1971,   t_1972;
/* u2_680 Output nets */
wire t_1973,   t_1974,   t_1975;
/* u2_681 Output nets */
wire t_1976,   t_1977,   t_1978;
/* u2_682 Output nets */
wire t_1979,   t_1980,   t_1981;
/* u2_683 Output nets */
wire t_1982,   t_1983,   t_1984;
/* u2_684 Output nets */
wire t_1985,   t_1986,   t_1987;
/* u2_685 Output nets */
wire t_1988,   t_1989,   t_1990;
/* u2_686 Output nets */
wire t_1991,   t_1992,   t_1993;
/* u2_687 Output nets */
wire t_1994,   t_1995,   t_1996;
/* u2_688 Output nets */
wire t_1997,   t_1998,   t_1999;
/* u1_689 Output nets */
wire t_2000,   t_2001;
/* u2_690 Output nets */
wire t_2002,   t_2003,   t_2004;
/* u2_691 Output nets */
wire t_2005,   t_2006,   t_2007;
/* u2_692 Output nets */
wire t_2008,   t_2009,   t_2010;
/* u2_693 Output nets */
wire t_2011,   t_2012,   t_2013;
/* u2_694 Output nets */
wire t_2014,   t_2015,   t_2016;
/* u2_695 Output nets */
wire t_2017,   t_2018,   t_2019;
/* u2_696 Output nets */
wire t_2020,   t_2021,   t_2022;
/* u2_697 Output nets */
wire t_2023,   t_2024,   t_2025;
/* u2_698 Output nets */
wire t_2026,   t_2027,   t_2028;
/* u2_699 Output nets */
wire t_2029,   t_2030,   t_2031;
/* u2_700 Output nets */
wire t_2032,   t_2033,   t_2034;
/* u2_701 Output nets */
wire t_2035,   t_2036,   t_2037;
/* u2_702 Output nets */
wire t_2038,   t_2039,   t_2040;
/* u2_703 Output nets */
wire t_2041,   t_2042,   t_2043;
/* u2_704 Output nets */
wire t_2044,   t_2045,   t_2046;
/* u2_705 Output nets */
wire t_2047,   t_2048,   t_2049;
/* u2_706 Output nets */
wire t_2050,   t_2051,   t_2052;
/* u2_707 Output nets */
wire t_2053,   t_2054,   t_2055;
/* u2_708 Output nets */
wire t_2056,   t_2057,   t_2058;
/* u2_709 Output nets */
wire t_2059,   t_2060,   t_2061;
/* u2_710 Output nets */
wire t_2062,   t_2063,   t_2064;
/* u2_711 Output nets */
wire t_2065,   t_2066,   t_2067;
/* u2_712 Output nets */
wire t_2068,   t_2069,   t_2070;
/* u2_713 Output nets */
wire t_2071,   t_2072,   t_2073;
/* u2_714 Output nets */
wire t_2074,   t_2075,   t_2076;
/* u2_715 Output nets */
wire t_2077,   t_2078,   t_2079;
/* u2_716 Output nets */
wire t_2080,   t_2081,   t_2082;
/* u2_717 Output nets */
wire t_2083,   t_2084,   t_2085;
/* u2_718 Output nets */
wire t_2086,   t_2087,   t_2088;
/* u2_719 Output nets */
wire t_2089,   t_2090,   t_2091;
/* u2_720 Output nets */
wire t_2092,   t_2093,   t_2094;
/* u2_721 Output nets */
wire t_2095,   t_2096,   t_2097;
/* u2_722 Output nets */
wire t_2098,   t_2099,   t_2100;
/* u2_723 Output nets */
wire t_2101,   t_2102,   t_2103;
/* u2_724 Output nets */
wire t_2104,   t_2105,   t_2106;
/* u2_725 Output nets */
wire t_2107,   t_2108,   t_2109;
/* u2_726 Output nets */
wire t_2110,   t_2111,   t_2112;
/* u2_727 Output nets */
wire t_2113,   t_2114,   t_2115;
/* u2_728 Output nets */
wire t_2116,   t_2117,   t_2118;
/* u0_729 Output nets */
wire t_2119,   t_2120;
/* u2_730 Output nets */
wire t_2121,   t_2122,   t_2123;
/* u2_731 Output nets */
wire t_2124,   t_2125,   t_2126;
/* u2_732 Output nets */
wire t_2127,   t_2128,   t_2129;
/* u2_733 Output nets */
wire t_2130,   t_2131,   t_2132;
/* u2_734 Output nets */
wire t_2133,   t_2134,   t_2135;
/* u2_735 Output nets */
wire t_2136,   t_2137,   t_2138;
/* u2_736 Output nets */
wire t_2139,   t_2140,   t_2141;
/* u2_737 Output nets */
wire t_2142,   t_2143,   t_2144;
/* u2_738 Output nets */
wire t_2145,   t_2146,   t_2147;
/* u2_739 Output nets */
wire t_2148,   t_2149,   t_2150;
/* u2_740 Output nets */
wire t_2151,   t_2152,   t_2153;
/* u2_741 Output nets */
wire t_2154,   t_2155,   t_2156;
/* u2_742 Output nets */
wire t_2157,   t_2158,   t_2159;
/* u2_743 Output nets */
wire t_2160,   t_2161,   t_2162;
/* u2_744 Output nets */
wire t_2163,   t_2164,   t_2165;
/* u2_745 Output nets */
wire t_2166,   t_2167,   t_2168;
/* u2_746 Output nets */
wire t_2169,   t_2170,   t_2171;
/* u2_747 Output nets */
wire t_2172,   t_2173,   t_2174;
/* u2_748 Output nets */
wire t_2175,   t_2176,   t_2177;
/* u2_749 Output nets */
wire t_2178,   t_2179,   t_2180;
/* u2_750 Output nets */
wire t_2181,   t_2182,   t_2183;
/* u2_751 Output nets */
wire t_2184,   t_2185,   t_2186;
/* u2_752 Output nets */
wire t_2187,   t_2188,   t_2189;
/* u2_753 Output nets */
wire t_2190,   t_2191,   t_2192;
/* u2_754 Output nets */
wire t_2193,   t_2194,   t_2195;
/* u2_755 Output nets */
wire t_2196,   t_2197,   t_2198;
/* u1_756 Output nets */
wire t_2199,   t_2200;
/* u2_757 Output nets */
wire t_2201,   t_2202,   t_2203;
/* u2_758 Output nets */
wire t_2204,   t_2205,   t_2206;
/* u2_759 Output nets */
wire t_2207,   t_2208,   t_2209;
/* u2_760 Output nets */
wire t_2210,   t_2211,   t_2212;
/* u2_761 Output nets */
wire t_2213,   t_2214,   t_2215;
/* u2_762 Output nets */
wire t_2216,   t_2217,   t_2218;
/* u2_763 Output nets */
wire t_2219,   t_2220,   t_2221;
/* u2_764 Output nets */
wire t_2222,   t_2223,   t_2224;
/* u2_765 Output nets */
wire t_2225,   t_2226,   t_2227;
/* u2_766 Output nets */
wire t_2228,   t_2229,   t_2230;
/* u2_767 Output nets */
wire t_2231,   t_2232,   t_2233;
/* u2_768 Output nets */
wire t_2234,   t_2235,   t_2236;
/* u2_769 Output nets */
wire t_2237,   t_2238,   t_2239;
/* u0_770 Output nets */
wire t_2240,   t_2241;
/* u2_771 Output nets */
wire t_2242,   t_2243,   t_2244;
/* u2_772 Output nets */
wire t_2245,   t_2246,   t_2247;
/* u2_773 Output nets */
wire t_2248,   t_2249,   t_2250;
/* u2_774 Output nets */
wire t_2251,   t_2252,   t_2253;
/* u2_775 Output nets */
wire t_2254,   t_2255,   t_2256;
/* u2_776 Output nets */
wire t_2257,   t_2258,   t_2259;
/* u2_777 Output nets */
wire t_2260,   t_2261,   t_2262;
/* u2_778 Output nets */
wire t_2263,   t_2264,   t_2265;
/* u2_779 Output nets */
wire t_2266,   t_2267,   t_2268;
/* u2_780 Output nets */
wire t_2269,   t_2270,   t_2271;
/* u2_781 Output nets */
wire t_2272,   t_2273,   t_2274;
/* u2_782 Output nets */
wire t_2275,   t_2276,   t_2277;
/* u2_783 Output nets */
wire t_2278,   t_2279,   t_2280;
/* u1_784 Output nets */
wire t_2281,   t_2282;
/* u2_785 Output nets */
wire t_2283,   t_2284,   t_2285;
/* u2_786 Output nets */
wire t_2286,   t_2287,   t_2288;
/* u2_787 Output nets */
wire t_2289,   t_2290,   t_2291;
/* u2_788 Output nets */
wire t_2292,   t_2293,   t_2294;
/* u2_789 Output nets */
wire t_2295,   t_2296,   t_2297;
/* u2_790 Output nets */
wire t_2298,   t_2299,   t_2300;
/* u2_791 Output nets */
wire t_2301,   t_2302,   t_2303;
/* u2_792 Output nets */
wire t_2304,   t_2305,   t_2306;
/* u2_793 Output nets */
wire t_2307,   t_2308,   t_2309;
/* u2_794 Output nets */
wire t_2310,   t_2311,   t_2312;
/* u2_795 Output nets */
wire t_2313,   t_2314,   t_2315;
/* u2_796 Output nets */
wire t_2316,   t_2317,   t_2318;
/* u2_797 Output nets */
wire t_2319,   t_2320,   t_2321;
/* u1_798 Output nets */
wire t_2322,   t_2323;
/* u2_799 Output nets */
wire t_2324,   t_2325,   t_2326;
/* u2_800 Output nets */
wire t_2327,   t_2328,   t_2329;
/* u2_801 Output nets */
wire t_2330,   t_2331,   t_2332;
/* u2_802 Output nets */
wire t_2333,   t_2334,   t_2335;
/* u2_803 Output nets */
wire t_2336,   t_2337,   t_2338;
/* u2_804 Output nets */
wire t_2339,   t_2340,   t_2341;
/* u2_805 Output nets */
wire t_2342,   t_2343,   t_2344;
/* u2_806 Output nets */
wire t_2345,   t_2346,   t_2347;
/* u2_807 Output nets */
wire t_2348,   t_2349,   t_2350;
/* u2_808 Output nets */
wire t_2351,   t_2352,   t_2353;
/* u2_809 Output nets */
wire t_2354,   t_2355,   t_2356;
/* u2_810 Output nets */
wire t_2357,   t_2358,   t_2359;
/* u2_811 Output nets */
wire t_2360,   t_2361,   t_2362;
/* u2_812 Output nets */
wire t_2363,   t_2364,   t_2365;
/* u2_813 Output nets */
wire t_2366,   t_2367,   t_2368;
/* u2_814 Output nets */
wire t_2369,   t_2370,   t_2371;
/* u2_815 Output nets */
wire t_2372,   t_2373,   t_2374;
/* u2_816 Output nets */
wire t_2375,   t_2376,   t_2377;
/* u2_817 Output nets */
wire t_2378,   t_2379,   t_2380;
/* u2_818 Output nets */
wire t_2381,   t_2382,   t_2383;
/* u2_819 Output nets */
wire t_2384,   t_2385,   t_2386;
/* u2_820 Output nets */
wire t_2387,   t_2388,   t_2389;
/* u2_821 Output nets */
wire t_2390,   t_2391,   t_2392;
/* u2_822 Output nets */
wire t_2393,   t_2394,   t_2395;
/* u2_823 Output nets */
wire t_2396,   t_2397,   t_2398;
/* u2_824 Output nets */
wire t_2399,   t_2400,   t_2401;
/* u2_825 Output nets */
wire t_2402,   t_2403,   t_2404;
/* u2_826 Output nets */
wire t_2405,   t_2406,   t_2407;
/* u2_827 Output nets */
wire t_2408,   t_2409,   t_2410;
/* u2_828 Output nets */
wire t_2411,   t_2412,   t_2413;
/* u2_829 Output nets */
wire t_2414,   t_2415,   t_2416;
/* u2_830 Output nets */
wire t_2417,   t_2418,   t_2419;
/* u2_831 Output nets */
wire t_2420,   t_2421,   t_2422;
/* u2_832 Output nets */
wire t_2423,   t_2424,   t_2425;
/* u2_833 Output nets */
wire t_2426,   t_2427,   t_2428;
/* u2_834 Output nets */
wire t_2429,   t_2430,   t_2431;
/* u2_835 Output nets */
wire t_2432,   t_2433,   t_2434;
/* u2_836 Output nets */
wire t_2435,   t_2436,   t_2437;
/* u2_837 Output nets */
wire t_2438,   t_2439,   t_2440;
/* u2_838 Output nets */
wire t_2441,   t_2442,   t_2443;
/* u2_839 Output nets */
wire t_2444,   t_2445,   t_2446;
/* u2_840 Output nets */
wire t_2447,   t_2448,   t_2449;
/* u0_841 Output nets */
wire t_2450,   t_2451;
/* u2_842 Output nets */
wire t_2452,   t_2453,   t_2454;
/* u2_843 Output nets */
wire t_2455,   t_2456,   t_2457;
/* u2_844 Output nets */
wire t_2458,   t_2459,   t_2460;
/* u2_845 Output nets */
wire t_2461,   t_2462,   t_2463;
/* u2_846 Output nets */
wire t_2464,   t_2465,   t_2466;
/* u2_847 Output nets */
wire t_2467,   t_2468,   t_2469;
/* u2_848 Output nets */
wire t_2470,   t_2471,   t_2472;
/* u2_849 Output nets */
wire t_2473,   t_2474,   t_2475;
/* u2_850 Output nets */
wire t_2476,   t_2477,   t_2478;
/* u2_851 Output nets */
wire t_2479,   t_2480,   t_2481;
/* u2_852 Output nets */
wire t_2482,   t_2483,   t_2484;
/* u2_853 Output nets */
wire t_2485,   t_2486,   t_2487;
/* u2_854 Output nets */
wire t_2488,   t_2489,   t_2490;
/* u2_855 Output nets */
wire t_2491,   t_2492,   t_2493;
/* u2_856 Output nets */
wire t_2494,   t_2495,   t_2496;
/* u2_857 Output nets */
wire t_2497,   t_2498,   t_2499;
/* u2_858 Output nets */
wire t_2500,   t_2501,   t_2502;
/* u2_859 Output nets */
wire t_2503,   t_2504,   t_2505;
/* u2_860 Output nets */
wire t_2506,   t_2507,   t_2508;
/* u2_861 Output nets */
wire t_2509,   t_2510,   t_2511;
/* u2_862 Output nets */
wire t_2512,   t_2513,   t_2514;
/* u2_863 Output nets */
wire t_2515,   t_2516,   t_2517;
/* u2_864 Output nets */
wire t_2518,   t_2519,   t_2520;
/* u2_865 Output nets */
wire t_2521,   t_2522,   t_2523;
/* u2_866 Output nets */
wire t_2524,   t_2525,   t_2526;
/* u2_867 Output nets */
wire t_2527,   t_2528,   t_2529;
/* u2_868 Output nets */
wire t_2530,   t_2531,   t_2532;
/* u2_869 Output nets */
wire t_2533,   t_2534,   t_2535;
/* u1_870 Output nets */
wire t_2536,   t_2537;
/* u2_871 Output nets */
wire t_2538,   t_2539,   t_2540;
/* u2_872 Output nets */
wire t_2541,   t_2542,   t_2543;
/* u2_873 Output nets */
wire t_2544,   t_2545,   t_2546;
/* u2_874 Output nets */
wire t_2547,   t_2548,   t_2549;
/* u2_875 Output nets */
wire t_2550,   t_2551,   t_2552;
/* u2_876 Output nets */
wire t_2553,   t_2554,   t_2555;
/* u2_877 Output nets */
wire t_2556,   t_2557,   t_2558;
/* u2_878 Output nets */
wire t_2559,   t_2560,   t_2561;
/* u2_879 Output nets */
wire t_2562,   t_2563,   t_2564;
/* u2_880 Output nets */
wire t_2565,   t_2566,   t_2567;
/* u2_881 Output nets */
wire t_2568,   t_2569,   t_2570;
/* u2_882 Output nets */
wire t_2571,   t_2572,   t_2573;
/* u2_883 Output nets */
wire t_2574,   t_2575,   t_2576;
/* u2_884 Output nets */
wire t_2577,   t_2578,   t_2579;
/* u0_885 Output nets */
wire t_2580,   t_2581;
/* u2_886 Output nets */
wire t_2582,   t_2583,   t_2584;
/* u2_887 Output nets */
wire t_2585,   t_2586,   t_2587;
/* u2_888 Output nets */
wire t_2588,   t_2589,   t_2590;
/* u2_889 Output nets */
wire t_2591,   t_2592,   t_2593;
/* u2_890 Output nets */
wire t_2594,   t_2595,   t_2596;
/* u2_891 Output nets */
wire t_2597,   t_2598,   t_2599;
/* u2_892 Output nets */
wire t_2600,   t_2601,   t_2602;
/* u2_893 Output nets */
wire t_2603,   t_2604,   t_2605;
/* u2_894 Output nets */
wire t_2606,   t_2607,   t_2608;
/* u2_895 Output nets */
wire t_2609,   t_2610,   t_2611;
/* u2_896 Output nets */
wire t_2612,   t_2613,   t_2614;
/* u2_897 Output nets */
wire t_2615,   t_2616,   t_2617;
/* u2_898 Output nets */
wire t_2618,   t_2619,   t_2620;
/* u2_899 Output nets */
wire t_2621,   t_2622,   t_2623;
/* u1_900 Output nets */
wire t_2624,   t_2625;
/* u2_901 Output nets */
wire t_2626,   t_2627,   t_2628;
/* u2_902 Output nets */
wire t_2629,   t_2630,   t_2631;
/* u2_903 Output nets */
wire t_2632,   t_2633,   t_2634;
/* u2_904 Output nets */
wire t_2635,   t_2636,   t_2637;
/* u2_905 Output nets */
wire t_2638,   t_2639,   t_2640;
/* u2_906 Output nets */
wire t_2641,   t_2642,   t_2643;
/* u2_907 Output nets */
wire t_2644,   t_2645,   t_2646;
/* u2_908 Output nets */
wire t_2647,   t_2648,   t_2649;
/* u2_909 Output nets */
wire t_2650,   t_2651,   t_2652;
/* u2_910 Output nets */
wire t_2653,   t_2654,   t_2655;
/* u2_911 Output nets */
wire t_2656,   t_2657,   t_2658;
/* u2_912 Output nets */
wire t_2659,   t_2660,   t_2661;
/* u2_913 Output nets */
wire t_2662,   t_2663,   t_2664;
/* u2_914 Output nets */
wire t_2665,   t_2666,   t_2667;
/* u1_915 Output nets */
wire t_2668,   t_2669;
/* u2_916 Output nets */
wire t_2670,   t_2671,   t_2672;
/* u2_917 Output nets */
wire t_2673,   t_2674,   t_2675;
/* u2_918 Output nets */
wire t_2676,   t_2677,   t_2678;
/* u2_919 Output nets */
wire t_2679,   t_2680,   t_2681;
/* u2_920 Output nets */
wire t_2682,   t_2683,   t_2684;
/* u2_921 Output nets */
wire t_2685,   t_2686,   t_2687;
/* u2_922 Output nets */
wire t_2688,   t_2689,   t_2690;
/* u2_923 Output nets */
wire t_2691,   t_2692,   t_2693;
/* u2_924 Output nets */
wire t_2694,   t_2695,   t_2696;
/* u2_925 Output nets */
wire t_2697,   t_2698,   t_2699;
/* u2_926 Output nets */
wire t_2700,   t_2701,   t_2702;
/* u2_927 Output nets */
wire t_2703,   t_2704,   t_2705;
/* u2_928 Output nets */
wire t_2706,   t_2707,   t_2708;
/* u2_929 Output nets */
wire t_2709,   t_2710,   t_2711;
/* u2_930 Output nets */
wire t_2712,   t_2713,   t_2714;
/* u2_931 Output nets */
wire t_2715,   t_2716,   t_2717;
/* u2_932 Output nets */
wire t_2718,   t_2719,   t_2720;
/* u2_933 Output nets */
wire t_2721,   t_2722,   t_2723;
/* u2_934 Output nets */
wire t_2724,   t_2725,   t_2726;
/* u2_935 Output nets */
wire t_2727,   t_2728,   t_2729;
/* u2_936 Output nets */
wire t_2730,   t_2731,   t_2732;
/* u2_937 Output nets */
wire t_2733,   t_2734,   t_2735;
/* u2_938 Output nets */
wire t_2736,   t_2737,   t_2738;
/* u2_939 Output nets */
wire t_2739,   t_2740,   t_2741;
/* u2_940 Output nets */
wire t_2742,   t_2743,   t_2744;
/* u2_941 Output nets */
wire t_2745,   t_2746,   t_2747;
/* u2_942 Output nets */
wire t_2748,   t_2749,   t_2750;
/* u2_943 Output nets */
wire t_2751,   t_2752,   t_2753;
/* u2_944 Output nets */
wire t_2754,   t_2755,   t_2756;
/* u2_945 Output nets */
wire t_2757,   t_2758,   t_2759;
/* u2_946 Output nets */
wire t_2760,   t_2761,   t_2762;
/* u2_947 Output nets */
wire t_2763,   t_2764,   t_2765;
/* u2_948 Output nets */
wire t_2766,   t_2767,   t_2768;
/* u2_949 Output nets */
wire t_2769,   t_2770,   t_2771;
/* u2_950 Output nets */
wire t_2772,   t_2773,   t_2774;
/* u2_951 Output nets */
wire t_2775,   t_2776,   t_2777;
/* u2_952 Output nets */
wire t_2778,   t_2779,   t_2780;
/* u2_953 Output nets */
wire t_2781,   t_2782,   t_2783;
/* u2_954 Output nets */
wire t_2784,   t_2785,   t_2786;
/* u2_955 Output nets */
wire t_2787,   t_2788,   t_2789;
/* u2_956 Output nets */
wire t_2790,   t_2791,   t_2792;
/* u2_957 Output nets */
wire t_2793,   t_2794,   t_2795;
/* u2_958 Output nets */
wire t_2796,   t_2797,   t_2798;
/* u2_959 Output nets */
wire t_2799,   t_2800,   t_2801;
/* u2_960 Output nets */
wire t_2802,   t_2803,   t_2804;
/* u0_961 Output nets */
wire t_2805,   t_2806;
/* u2_962 Output nets */
wire t_2807,   t_2808,   t_2809;
/* u2_963 Output nets */
wire t_2810,   t_2811,   t_2812;
/* u2_964 Output nets */
wire t_2813,   t_2814,   t_2815;
/* u2_965 Output nets */
wire t_2816,   t_2817,   t_2818;
/* u2_966 Output nets */
wire t_2819,   t_2820,   t_2821;
/* u2_967 Output nets */
wire t_2822,   t_2823,   t_2824;
/* u2_968 Output nets */
wire t_2825,   t_2826,   t_2827;
/* u2_969 Output nets */
wire t_2828,   t_2829,   t_2830;
/* u2_970 Output nets */
wire t_2831,   t_2832,   t_2833;
/* u2_971 Output nets */
wire t_2834,   t_2835,   t_2836;
/* u2_972 Output nets */
wire t_2837,   t_2838,   t_2839;
/* u2_973 Output nets */
wire t_2840,   t_2841,   t_2842;
/* u2_974 Output nets */
wire t_2843,   t_2844,   t_2845;
/* u2_975 Output nets */
wire t_2846,   t_2847,   t_2848;
/* u2_976 Output nets */
wire t_2849,   t_2850,   t_2851;
/* u2_977 Output nets */
wire t_2852,   t_2853,   t_2854;
/* u2_978 Output nets */
wire t_2855,   t_2856,   t_2857;
/* u2_979 Output nets */
wire t_2858,   t_2859,   t_2860;
/* u2_980 Output nets */
wire t_2861,   t_2862,   t_2863;
/* u2_981 Output nets */
wire t_2864,   t_2865,   t_2866;
/* u2_982 Output nets */
wire t_2867,   t_2868,   t_2869;
/* u2_983 Output nets */
wire t_2870,   t_2871,   t_2872;
/* u2_984 Output nets */
wire t_2873,   t_2874,   t_2875;
/* u2_985 Output nets */
wire t_2876,   t_2877,   t_2878;
/* u2_986 Output nets */
wire t_2879,   t_2880,   t_2881;
/* u2_987 Output nets */
wire t_2882,   t_2883,   t_2884;
/* u2_988 Output nets */
wire t_2885,   t_2886,   t_2887;
/* u2_989 Output nets */
wire t_2888,   t_2889,   t_2890;
/* u2_990 Output nets */
wire t_2891,   t_2892,   t_2893;
/* u2_991 Output nets */
wire t_2894,   t_2895,   t_2896;
/* u1_992 Output nets */
wire t_2897,   t_2898;
/* u2_993 Output nets */
wire t_2899,   t_2900,   t_2901;
/* u2_994 Output nets */
wire t_2902,   t_2903,   t_2904;
/* u2_995 Output nets */
wire t_2905,   t_2906,   t_2907;
/* u2_996 Output nets */
wire t_2908,   t_2909,   t_2910;
/* u2_997 Output nets */
wire t_2911,   t_2912,   t_2913;
/* u2_998 Output nets */
wire t_2914,   t_2915,   t_2916;
/* u2_999 Output nets */
wire t_2917,   t_2918,   t_2919;
/* u2_1000 Output nets */
wire t_2920,   t_2921,   t_2922;
/* u2_1001 Output nets */
wire t_2923,   t_2924,   t_2925;
/* u2_1002 Output nets */
wire t_2926,   t_2927,   t_2928;
/* u2_1003 Output nets */
wire t_2929,   t_2930,   t_2931;
/* u2_1004 Output nets */
wire t_2932,   t_2933,   t_2934;
/* u2_1005 Output nets */
wire t_2935,   t_2936,   t_2937;
/* u2_1006 Output nets */
wire t_2938,   t_2939,   t_2940;
/* u2_1007 Output nets */
wire t_2941,   t_2942,   t_2943;
/* u0_1008 Output nets */
wire t_2944,   t_2945;
/* u2_1009 Output nets */
wire t_2946,   t_2947,   t_2948;
/* u2_1010 Output nets */
wire t_2949,   t_2950,   t_2951;
/* u2_1011 Output nets */
wire t_2952,   t_2953,   t_2954;
/* u2_1012 Output nets */
wire t_2955,   t_2956,   t_2957;
/* u2_1013 Output nets */
wire t_2958,   t_2959,   t_2960;
/* u2_1014 Output nets */
wire t_2961,   t_2962,   t_2963;
/* u2_1015 Output nets */
wire t_2964,   t_2965,   t_2966;
/* u2_1016 Output nets */
wire t_2967,   t_2968,   t_2969;
/* u2_1017 Output nets */
wire t_2970,   t_2971,   t_2972;
/* u2_1018 Output nets */
wire t_2973,   t_2974,   t_2975;
/* u2_1019 Output nets */
wire t_2976,   t_2977,   t_2978;
/* u2_1020 Output nets */
wire t_2979,   t_2980,   t_2981;
/* u2_1021 Output nets */
wire t_2982,   t_2983,   t_2984;
/* u2_1022 Output nets */
wire t_2985,   t_2986,   t_2987;
/* u2_1023 Output nets */
wire t_2988,   t_2989,   t_2990;
/* u1_1024 Output nets */
wire t_2991,   t_2992;
/* u2_1025 Output nets */
wire t_2993,   t_2994,   t_2995;
/* u2_1026 Output nets */
wire t_2996,   t_2997,   t_2998;
/* u2_1027 Output nets */
wire t_2999,   t_3000,   t_3001;
/* u2_1028 Output nets */
wire t_3002,   t_3003,   t_3004;
/* u2_1029 Output nets */
wire t_3005,   t_3006,   t_3007;
/* u2_1030 Output nets */
wire t_3008,   t_3009,   t_3010;
/* u2_1031 Output nets */
wire t_3011,   t_3012,   t_3013;
/* u2_1032 Output nets */
wire t_3014,   t_3015,   t_3016;
/* u2_1033 Output nets */
wire t_3017,   t_3018,   t_3019;
/* u2_1034 Output nets */
wire t_3020,   t_3021,   t_3022;
/* u2_1035 Output nets */
wire t_3023,   t_3024,   t_3025;
/* u2_1036 Output nets */
wire t_3026,   t_3027,   t_3028;
/* u2_1037 Output nets */
wire t_3029,   t_3030,   t_3031;
/* u2_1038 Output nets */
wire t_3032,   t_3033,   t_3034;
/* u2_1039 Output nets */
wire t_3035,   t_3036,   t_3037;
/* u1_1040 Output nets */
wire t_3038,   t_3039;
/* u2_1041 Output nets */
wire t_3040,   t_3041,   t_3042;
/* u2_1042 Output nets */
wire t_3043,   t_3044,   t_3045;
/* u2_1043 Output nets */
wire t_3046,   t_3047,   t_3048;
/* u2_1044 Output nets */
wire t_3049,   t_3050,   t_3051;
/* u2_1045 Output nets */
wire t_3052,   t_3053,   t_3054;
/* u2_1046 Output nets */
wire t_3055,   t_3056,   t_3057;
/* u2_1047 Output nets */
wire t_3058,   t_3059,   t_3060;
/* u2_1048 Output nets */
wire t_3061,   t_3062,   t_3063;
/* u2_1049 Output nets */
wire t_3064,   t_3065,   t_3066;
/* u2_1050 Output nets */
wire t_3067,   t_3068,   t_3069;
/* u2_1051 Output nets */
wire t_3070,   t_3071,   t_3072;
/* u2_1052 Output nets */
wire t_3073,   t_3074,   t_3075;
/* u2_1053 Output nets */
wire t_3076,   t_3077,   t_3078;
/* u2_1054 Output nets */
wire t_3079,   t_3080,   t_3081;
/* u2_1055 Output nets */
wire t_3082,   t_3083,   t_3084;
/* u2_1056 Output nets */
wire t_3085,   t_3086,   t_3087;
/* u2_1057 Output nets */
wire t_3088,   t_3089,   t_3090;
/* u2_1058 Output nets */
wire t_3091,   t_3092,   t_3093;
/* u2_1059 Output nets */
wire t_3094,   t_3095,   t_3096;
/* u2_1060 Output nets */
wire t_3097,   t_3098,   t_3099;
/* u2_1061 Output nets */
wire t_3100,   t_3101,   t_3102;
/* u2_1062 Output nets */
wire t_3103,   t_3104,   t_3105;
/* u2_1063 Output nets */
wire t_3106,   t_3107,   t_3108;
/* u2_1064 Output nets */
wire t_3109,   t_3110,   t_3111;
/* u2_1065 Output nets */
wire t_3112,   t_3113,   t_3114;
/* u2_1066 Output nets */
wire t_3115,   t_3116,   t_3117;
/* u2_1067 Output nets */
wire t_3118,   t_3119,   t_3120;
/* u2_1068 Output nets */
wire t_3121,   t_3122,   t_3123;
/* u2_1069 Output nets */
wire t_3124,   t_3125,   t_3126;
/* u2_1070 Output nets */
wire t_3127,   t_3128,   t_3129;
/* u2_1071 Output nets */
wire t_3130,   t_3131,   t_3132;
/* u2_1072 Output nets */
wire t_3133,   t_3134,   t_3135;
/* u2_1073 Output nets */
wire t_3136,   t_3137,   t_3138;
/* u2_1074 Output nets */
wire t_3139,   t_3140,   t_3141;
/* u2_1075 Output nets */
wire t_3142,   t_3143,   t_3144;
/* u2_1076 Output nets */
wire t_3145,   t_3146,   t_3147;
/* u2_1077 Output nets */
wire t_3148,   t_3149,   t_3150;
/* u2_1078 Output nets */
wire t_3151,   t_3152,   t_3153;
/* u2_1079 Output nets */
wire t_3154,   t_3155,   t_3156;
/* u2_1080 Output nets */
wire t_3157,   t_3158,   t_3159;
/* u2_1081 Output nets */
wire t_3160,   t_3161,   t_3162;
/* u2_1082 Output nets */
wire t_3163,   t_3164,   t_3165;
/* u2_1083 Output nets */
wire t_3166,   t_3167,   t_3168;
/* u2_1084 Output nets */
wire t_3169,   t_3170,   t_3171;
/* u2_1085 Output nets */
wire t_3172,   t_3173,   t_3174;
/* u2_1086 Output nets */
wire t_3175,   t_3176,   t_3177;
/* u2_1087 Output nets */
wire t_3178,   t_3179,   t_3180;
/* u2_1088 Output nets */
wire t_3181,   t_3182,   t_3183;
/* u2_1089 Output nets */
wire t_3184,   t_3185,   t_3186;
/* u2_1090 Output nets */
wire t_3187,   t_3188,   t_3189;
/* u2_1091 Output nets */
wire t_3190,   t_3191,   t_3192;
/* u2_1092 Output nets */
wire t_3193,   t_3194,   t_3195;
/* u2_1093 Output nets */
wire t_3196,   t_3197,   t_3198;
/* u2_1094 Output nets */
wire t_3199,   t_3200,   t_3201;
/* u2_1095 Output nets */
wire t_3202,   t_3203,   t_3204;
/* u2_1096 Output nets */
wire t_3205,   t_3206,   t_3207;
/* u2_1097 Output nets */
wire t_3208,   t_3209,   t_3210;
/* u2_1098 Output nets */
wire t_3211,   t_3212,   t_3213;
/* u2_1099 Output nets */
wire t_3214,   t_3215,   t_3216;
/* u2_1100 Output nets */
wire t_3217,   t_3218,   t_3219;
/* u2_1101 Output nets */
wire t_3220,   t_3221,   t_3222;
/* u2_1102 Output nets */
wire t_3223,   t_3224,   t_3225;
/* u2_1103 Output nets */
wire t_3226,   t_3227,   t_3228;
/* u2_1104 Output nets */
wire t_3229,   t_3230,   t_3231;
/* u2_1105 Output nets */
wire t_3232,   t_3233,   t_3234;
/* u2_1106 Output nets */
wire t_3235,   t_3236,   t_3237;
/* u2_1107 Output nets */
wire t_3238,   t_3239,   t_3240;
/* u2_1108 Output nets */
wire t_3241,   t_3242,   t_3243;
/* u2_1109 Output nets */
wire t_3244,   t_3245,   t_3246;
/* u2_1110 Output nets */
wire t_3247,   t_3248,   t_3249;
/* u2_1111 Output nets */
wire t_3250,   t_3251,   t_3252;
/* u2_1112 Output nets */
wire t_3253,   t_3254,   t_3255;
/* u2_1113 Output nets */
wire t_3256,   t_3257,   t_3258;
/* u2_1114 Output nets */
wire t_3259,   t_3260,   t_3261;
/* u2_1115 Output nets */
wire t_3262,   t_3263,   t_3264;
/* u2_1116 Output nets */
wire t_3265,   t_3266,   t_3267;
/* u2_1117 Output nets */
wire t_3268,   t_3269,   t_3270;
/* u2_1118 Output nets */
wire t_3271,   t_3272,   t_3273;
/* u2_1119 Output nets */
wire t_3274,   t_3275,   t_3276;
/* u2_1120 Output nets */
wire t_3277,   t_3278,   t_3279;
/* u2_1121 Output nets */
wire t_3280,   t_3281,   t_3282;
/* u2_1122 Output nets */
wire t_3283,   t_3284,   t_3285;
/* u2_1123 Output nets */
wire t_3286,   t_3287,   t_3288;
/* u2_1124 Output nets */
wire t_3289,   t_3290,   t_3291;
/* u2_1125 Output nets */
wire t_3292,   t_3293,   t_3294;
/* u2_1126 Output nets */
wire t_3295,   t_3296,   t_3297;
/* u2_1127 Output nets */
wire t_3298,   t_3299,   t_3300;
/* u2_1128 Output nets */
wire t_3301,   t_3302,   t_3303;
/* u2_1129 Output nets */
wire t_3304,   t_3305,   t_3306;
/* u2_1130 Output nets */
wire t_3307,   t_3308,   t_3309;
/* u2_1131 Output nets */
wire t_3310,   t_3311,   t_3312;
/* u2_1132 Output nets */
wire t_3313,   t_3314,   t_3315;
/* u2_1133 Output nets */
wire t_3316,   t_3317,   t_3318;
/* u2_1134 Output nets */
wire t_3319,   t_3320,   t_3321;
/* u2_1135 Output nets */
wire t_3322,   t_3323,   t_3324;
/* u2_1136 Output nets */
wire t_3325,   t_3326,   t_3327;
/* u2_1137 Output nets */
wire t_3328,   t_3329,   t_3330;
/* u2_1138 Output nets */
wire t_3331,   t_3332,   t_3333;
/* u2_1139 Output nets */
wire t_3334,   t_3335,   t_3336;
/* u2_1140 Output nets */
wire t_3337,   t_3338,   t_3339;
/* u2_1141 Output nets */
wire t_3340,   t_3341,   t_3342;
/* u2_1142 Output nets */
wire t_3343,   t_3344,   t_3345;
/* u2_1143 Output nets */
wire t_3346,   t_3347,   t_3348;
/* u2_1144 Output nets */
wire t_3349,   t_3350,   t_3351;
/* u2_1145 Output nets */
wire t_3352,   t_3353,   t_3354;
/* u2_1146 Output nets */
wire t_3355,   t_3356,   t_3357;
/* u2_1147 Output nets */
wire t_3358,   t_3359,   t_3360;
/* u2_1148 Output nets */
wire t_3361,   t_3362,   t_3363;
/* u2_1149 Output nets */
wire t_3364,   t_3365,   t_3366;
/* u2_1150 Output nets */
wire t_3367,   t_3368,   t_3369;
/* u2_1151 Output nets */
wire t_3370,   t_3371,   t_3372;
/* u1_1152 Output nets */
wire t_3373,   t_3374;
/* u2_1153 Output nets */
wire t_3375,   t_3376,   t_3377;
/* u2_1154 Output nets */
wire t_3378,   t_3379,   t_3380;
/* u2_1155 Output nets */
wire t_3381,   t_3382,   t_3383;
/* u2_1156 Output nets */
wire t_3384,   t_3385,   t_3386;
/* u2_1157 Output nets */
wire t_3387,   t_3388,   t_3389;
/* u2_1158 Output nets */
wire t_3390,   t_3391,   t_3392;
/* u2_1159 Output nets */
wire t_3393,   t_3394,   t_3395;
/* u2_1160 Output nets */
wire t_3396,   t_3397,   t_3398;
/* u2_1161 Output nets */
wire t_3399,   t_3400,   t_3401;
/* u2_1162 Output nets */
wire t_3402,   t_3403,   t_3404;
/* u2_1163 Output nets */
wire t_3405,   t_3406,   t_3407;
/* u2_1164 Output nets */
wire t_3408,   t_3409,   t_3410;
/* u2_1165 Output nets */
wire t_3411,   t_3412,   t_3413;
/* u2_1166 Output nets */
wire t_3414,   t_3415,   t_3416;
/* u2_1167 Output nets */
wire t_3417,   t_3418,   t_3419;
/* u1_1168 Output nets */
wire t_3420,   t_3421;
/* u2_1169 Output nets */
wire t_3422,   t_3423,   t_3424;
/* u2_1170 Output nets */
wire t_3425,   t_3426,   t_3427;
/* u2_1171 Output nets */
wire t_3428,   t_3429,   t_3430;
/* u2_1172 Output nets */
wire t_3431,   t_3432,   t_3433;
/* u2_1173 Output nets */
wire t_3434,   t_3435,   t_3436;
/* u2_1174 Output nets */
wire t_3437,   t_3438,   t_3439;
/* u2_1175 Output nets */
wire t_3440,   t_3441,   t_3442;
/* u2_1176 Output nets */
wire t_3443,   t_3444,   t_3445;
/* u2_1177 Output nets */
wire t_3446,   t_3447,   t_3448;
/* u2_1178 Output nets */
wire t_3449,   t_3450,   t_3451;
/* u2_1179 Output nets */
wire t_3452,   t_3453,   t_3454;
/* u2_1180 Output nets */
wire t_3455,   t_3456,   t_3457;
/* u2_1181 Output nets */
wire t_3458,   t_3459,   t_3460;
/* u2_1182 Output nets */
wire t_3461,   t_3462,   t_3463;
/* u2_1183 Output nets */
wire t_3464,   t_3465,   t_3466;
/* u0_1184 Output nets */
wire t_3467,   t_3468;
/* u2_1185 Output nets */
wire t_3469,   t_3470,   t_3471;
/* u2_1186 Output nets */
wire t_3472,   t_3473,   t_3474;
/* u2_1187 Output nets */
wire t_3475,   t_3476,   t_3477;
/* u2_1188 Output nets */
wire t_3478,   t_3479,   t_3480;
/* u2_1189 Output nets */
wire t_3481,   t_3482,   t_3483;
/* u2_1190 Output nets */
wire t_3484,   t_3485,   t_3486;
/* u2_1191 Output nets */
wire t_3487,   t_3488,   t_3489;
/* u2_1192 Output nets */
wire t_3490,   t_3491,   t_3492;
/* u2_1193 Output nets */
wire t_3493,   t_3494,   t_3495;
/* u2_1194 Output nets */
wire t_3496,   t_3497,   t_3498;
/* u2_1195 Output nets */
wire t_3499,   t_3500,   t_3501;
/* u2_1196 Output nets */
wire t_3502,   t_3503,   t_3504;
/* u2_1197 Output nets */
wire t_3505,   t_3506,   t_3507;
/* u2_1198 Output nets */
wire t_3508,   t_3509,   t_3510;
/* u2_1199 Output nets */
wire t_3511,   t_3512,   t_3513;
/* u0_1200 Output nets */
wire t_3514,   t_3515;
/* u2_1201 Output nets */
wire t_3516,   t_3517,   t_3518;
/* u2_1202 Output nets */
wire t_3519,   t_3520,   t_3521;
/* u2_1203 Output nets */
wire t_3522,   t_3523,   t_3524;
/* u2_1204 Output nets */
wire t_3525,   t_3526,   t_3527;
/* u2_1205 Output nets */
wire t_3528,   t_3529,   t_3530;
/* u2_1206 Output nets */
wire t_3531,   t_3532,   t_3533;
/* u2_1207 Output nets */
wire t_3534,   t_3535,   t_3536;
/* u2_1208 Output nets */
wire t_3537,   t_3538,   t_3539;
/* u2_1209 Output nets */
wire t_3540,   t_3541,   t_3542;
/* u2_1210 Output nets */
wire t_3543,   t_3544,   t_3545;
/* u2_1211 Output nets */
wire t_3546,   t_3547,   t_3548;
/* u2_1212 Output nets */
wire t_3549,   t_3550,   t_3551;
/* u2_1213 Output nets */
wire t_3552,   t_3553,   t_3554;
/* u2_1214 Output nets */
wire t_3555,   t_3556,   t_3557;
/* u2_1215 Output nets */
wire t_3558,   t_3559,   t_3560;
/* u2_1216 Output nets */
wire t_3561,   t_3562,   t_3563;
/* u2_1217 Output nets */
wire t_3564,   t_3565,   t_3566;
/* u2_1218 Output nets */
wire t_3567,   t_3568,   t_3569;
/* u2_1219 Output nets */
wire t_3570,   t_3571,   t_3572;
/* u2_1220 Output nets */
wire t_3573,   t_3574,   t_3575;
/* u2_1221 Output nets */
wire t_3576,   t_3577,   t_3578;
/* u2_1222 Output nets */
wire t_3579,   t_3580,   t_3581;
/* u2_1223 Output nets */
wire t_3582,   t_3583,   t_3584;
/* u2_1224 Output nets */
wire t_3585,   t_3586,   t_3587;
/* u2_1225 Output nets */
wire t_3588,   t_3589,   t_3590;
/* u2_1226 Output nets */
wire t_3591,   t_3592,   t_3593;
/* u2_1227 Output nets */
wire t_3594,   t_3595,   t_3596;
/* u2_1228 Output nets */
wire t_3597,   t_3598,   t_3599;
/* u2_1229 Output nets */
wire t_3600,   t_3601,   t_3602;
/* u2_1230 Output nets */
wire t_3603,   t_3604,   t_3605;
/* u2_1231 Output nets */
wire t_3606,   t_3607,   t_3608;
/* u2_1232 Output nets */
wire t_3609,   t_3610,   t_3611;
/* u2_1233 Output nets */
wire t_3612,   t_3613,   t_3614;
/* u2_1234 Output nets */
wire t_3615,   t_3616,   t_3617;
/* u2_1235 Output nets */
wire t_3618,   t_3619,   t_3620;
/* u2_1236 Output nets */
wire t_3621,   t_3622,   t_3623;
/* u2_1237 Output nets */
wire t_3624,   t_3625,   t_3626;
/* u2_1238 Output nets */
wire t_3627,   t_3628,   t_3629;
/* u2_1239 Output nets */
wire t_3630,   t_3631,   t_3632;
/* u2_1240 Output nets */
wire t_3633,   t_3634,   t_3635;
/* u2_1241 Output nets */
wire t_3636,   t_3637,   t_3638;
/* u2_1242 Output nets */
wire t_3639,   t_3640,   t_3641;
/* u2_1243 Output nets */
wire t_3642,   t_3643,   t_3644;
/* u2_1244 Output nets */
wire t_3645,   t_3646,   t_3647;
/* u2_1245 Output nets */
wire t_3648,   t_3649,   t_3650;
/* u2_1246 Output nets */
wire t_3651,   t_3652,   t_3653;
/* u2_1247 Output nets */
wire t_3654,   t_3655,   t_3656;
/* u2_1248 Output nets */
wire t_3657,   t_3658,   t_3659;
/* u2_1249 Output nets */
wire t_3660,   t_3661,   t_3662;
/* u2_1250 Output nets */
wire t_3663,   t_3664,   t_3665;
/* u2_1251 Output nets */
wire t_3666,   t_3667,   t_3668;
/* u2_1252 Output nets */
wire t_3669,   t_3670,   t_3671;
/* u2_1253 Output nets */
wire t_3672,   t_3673,   t_3674;
/* u2_1254 Output nets */
wire t_3675,   t_3676,   t_3677;
/* u2_1255 Output nets */
wire t_3678,   t_3679,   t_3680;
/* u2_1256 Output nets */
wire t_3681,   t_3682,   t_3683;
/* u2_1257 Output nets */
wire t_3684,   t_3685,   t_3686;
/* u2_1258 Output nets */
wire t_3687,   t_3688,   t_3689;
/* u2_1259 Output nets */
wire t_3690,   t_3691,   t_3692;
/* u2_1260 Output nets */
wire t_3693,   t_3694,   t_3695;
/* u2_1261 Output nets */
wire t_3696,   t_3697,   t_3698;
/* u2_1262 Output nets */
wire t_3699,   t_3700,   t_3701;
/* u2_1263 Output nets */
wire t_3702,   t_3703,   t_3704;
/* u2_1264 Output nets */
wire t_3705,   t_3706,   t_3707;
/* u2_1265 Output nets */
wire t_3708,   t_3709,   t_3710;
/* u2_1266 Output nets */
wire t_3711,   t_3712,   t_3713;
/* u2_1267 Output nets */
wire t_3714,   t_3715,   t_3716;
/* u2_1268 Output nets */
wire t_3717,   t_3718,   t_3719;
/* u2_1269 Output nets */
wire t_3720,   t_3721,   t_3722;
/* u2_1270 Output nets */
wire t_3723,   t_3724,   t_3725;
/* u2_1271 Output nets */
wire t_3726,   t_3727,   t_3728;
/* u2_1272 Output nets */
wire t_3729,   t_3730,   t_3731;
/* u2_1273 Output nets */
wire t_3732,   t_3733,   t_3734;
/* u2_1274 Output nets */
wire t_3735,   t_3736,   t_3737;
/* u1_1275 Output nets */
wire t_3738,   t_3739;
/* u2_1276 Output nets */
wire t_3740,   t_3741,   t_3742;
/* u2_1277 Output nets */
wire t_3743,   t_3744,   t_3745;
/* u2_1278 Output nets */
wire t_3746,   t_3747,   t_3748;
/* u2_1279 Output nets */
wire t_3749,   t_3750,   t_3751;
/* u2_1280 Output nets */
wire t_3752,   t_3753,   t_3754;
/* u2_1281 Output nets */
wire t_3755,   t_3756,   t_3757;
/* u2_1282 Output nets */
wire t_3758,   t_3759,   t_3760;
/* u2_1283 Output nets */
wire t_3761,   t_3762,   t_3763;
/* u2_1284 Output nets */
wire t_3764,   t_3765,   t_3766;
/* u2_1285 Output nets */
wire t_3767,   t_3768,   t_3769;
/* u2_1286 Output nets */
wire t_3770,   t_3771,   t_3772;
/* u2_1287 Output nets */
wire t_3773,   t_3774,   t_3775;
/* u2_1288 Output nets */
wire t_3776,   t_3777,   t_3778;
/* u2_1289 Output nets */
wire t_3779,   t_3780,   t_3781;
/* u1_1290 Output nets */
wire t_3782,   t_3783;
/* u2_1291 Output nets */
wire t_3784,   t_3785,   t_3786;
/* u2_1292 Output nets */
wire t_3787,   t_3788,   t_3789;
/* u2_1293 Output nets */
wire t_3790,   t_3791,   t_3792;
/* u2_1294 Output nets */
wire t_3793,   t_3794,   t_3795;
/* u2_1295 Output nets */
wire t_3796,   t_3797,   t_3798;
/* u2_1296 Output nets */
wire t_3799,   t_3800,   t_3801;
/* u2_1297 Output nets */
wire t_3802,   t_3803,   t_3804;
/* u2_1298 Output nets */
wire t_3805,   t_3806,   t_3807;
/* u2_1299 Output nets */
wire t_3808,   t_3809,   t_3810;
/* u2_1300 Output nets */
wire t_3811,   t_3812,   t_3813;
/* u2_1301 Output nets */
wire t_3814,   t_3815,   t_3816;
/* u2_1302 Output nets */
wire t_3817,   t_3818,   t_3819;
/* u2_1303 Output nets */
wire t_3820,   t_3821,   t_3822;
/* u2_1304 Output nets */
wire t_3823,   t_3824,   t_3825;
/* u0_1305 Output nets */
wire t_3826,   t_3827;
/* u2_1306 Output nets */
wire t_3828,   t_3829,   t_3830;
/* u2_1307 Output nets */
wire t_3831,   t_3832,   t_3833;
/* u2_1308 Output nets */
wire t_3834,   t_3835,   t_3836;
/* u2_1309 Output nets */
wire t_3837,   t_3838,   t_3839;
/* u2_1310 Output nets */
wire t_3840,   t_3841,   t_3842;
/* u2_1311 Output nets */
wire t_3843,   t_3844,   t_3845;
/* u2_1312 Output nets */
wire t_3846,   t_3847,   t_3848;
/* u2_1313 Output nets */
wire t_3849,   t_3850,   t_3851;
/* u2_1314 Output nets */
wire t_3852,   t_3853,   t_3854;
/* u2_1315 Output nets */
wire t_3855,   t_3856,   t_3857;
/* u2_1316 Output nets */
wire t_3858,   t_3859,   t_3860;
/* u2_1317 Output nets */
wire t_3861,   t_3862,   t_3863;
/* u2_1318 Output nets */
wire t_3864,   t_3865,   t_3866;
/* u2_1319 Output nets */
wire t_3867,   t_3868,   t_3869;
/* u0_1320 Output nets */
wire t_3870,   t_3871;
/* u2_1321 Output nets */
wire t_3872,   t_3873,   t_3874;
/* u2_1322 Output nets */
wire t_3875,   t_3876,   t_3877;
/* u2_1323 Output nets */
wire t_3878,   t_3879,   t_3880;
/* u2_1324 Output nets */
wire t_3881,   t_3882,   t_3883;
/* u2_1325 Output nets */
wire t_3884,   t_3885,   t_3886;
/* u2_1326 Output nets */
wire t_3887,   t_3888,   t_3889;
/* u2_1327 Output nets */
wire t_3890,   t_3891,   t_3892;
/* u2_1328 Output nets */
wire t_3893,   t_3894,   t_3895;
/* u2_1329 Output nets */
wire t_3896,   t_3897,   t_3898;
/* u2_1330 Output nets */
wire t_3899,   t_3900,   t_3901;
/* u2_1331 Output nets */
wire t_3902,   t_3903,   t_3904;
/* u2_1332 Output nets */
wire t_3905,   t_3906,   t_3907;
/* u2_1333 Output nets */
wire t_3908,   t_3909,   t_3910;
/* u2_1334 Output nets */
wire t_3911,   t_3912,   t_3913;
/* u2_1335 Output nets */
wire t_3914,   t_3915,   t_3916;
/* u2_1336 Output nets */
wire t_3917,   t_3918,   t_3919;
/* u2_1337 Output nets */
wire t_3920,   t_3921,   t_3922;
/* u2_1338 Output nets */
wire t_3923,   t_3924,   t_3925;
/* u2_1339 Output nets */
wire t_3926,   t_3927,   t_3928;
/* u2_1340 Output nets */
wire t_3929,   t_3930,   t_3931;
/* u2_1341 Output nets */
wire t_3932,   t_3933,   t_3934;
/* u2_1342 Output nets */
wire t_3935,   t_3936,   t_3937;
/* u2_1343 Output nets */
wire t_3938,   t_3939,   t_3940;
/* u2_1344 Output nets */
wire t_3941,   t_3942,   t_3943;
/* u2_1345 Output nets */
wire t_3944,   t_3945,   t_3946;
/* u2_1346 Output nets */
wire t_3947,   t_3948,   t_3949;
/* u2_1347 Output nets */
wire t_3950,   t_3951,   t_3952;
/* u2_1348 Output nets */
wire t_3953,   t_3954,   t_3955;
/* u2_1349 Output nets */
wire t_3956,   t_3957,   t_3958;
/* u2_1350 Output nets */
wire t_3959,   t_3960,   t_3961;
/* u2_1351 Output nets */
wire t_3962,   t_3963,   t_3964;
/* u2_1352 Output nets */
wire t_3965,   t_3966,   t_3967;
/* u2_1353 Output nets */
wire t_3968,   t_3969,   t_3970;
/* u2_1354 Output nets */
wire t_3971,   t_3972,   t_3973;
/* u2_1355 Output nets */
wire t_3974,   t_3975,   t_3976;
/* u2_1356 Output nets */
wire t_3977,   t_3978,   t_3979;
/* u2_1357 Output nets */
wire t_3980,   t_3981,   t_3982;
/* u2_1358 Output nets */
wire t_3983,   t_3984,   t_3985;
/* u2_1359 Output nets */
wire t_3986,   t_3987,   t_3988;
/* u2_1360 Output nets */
wire t_3989,   t_3990,   t_3991;
/* u2_1361 Output nets */
wire t_3992,   t_3993,   t_3994;
/* u2_1362 Output nets */
wire t_3995,   t_3996,   t_3997;
/* u2_1363 Output nets */
wire t_3998,   t_3999,   t_4000;
/* u2_1364 Output nets */
wire t_4001,   t_4002,   t_4003;
/* u2_1365 Output nets */
wire t_4004,   t_4005,   t_4006;
/* u2_1366 Output nets */
wire t_4007,   t_4008,   t_4009;
/* u2_1367 Output nets */
wire t_4010,   t_4011,   t_4012;
/* u2_1368 Output nets */
wire t_4013,   t_4014,   t_4015;
/* u2_1369 Output nets */
wire t_4016,   t_4017,   t_4018;
/* u2_1370 Output nets */
wire t_4019,   t_4020,   t_4021;
/* u2_1371 Output nets */
wire t_4022,   t_4023,   t_4024;
/* u2_1372 Output nets */
wire t_4025,   t_4026,   t_4027;
/* u2_1373 Output nets */
wire t_4028,   t_4029,   t_4030;
/* u2_1374 Output nets */
wire t_4031,   t_4032,   t_4033;
/* u2_1375 Output nets */
wire t_4034,   t_4035,   t_4036;
/* u2_1376 Output nets */
wire t_4037,   t_4038,   t_4039;
/* u2_1377 Output nets */
wire t_4040,   t_4041,   t_4042;
/* u2_1378 Output nets */
wire t_4043,   t_4044,   t_4045;
/* u2_1379 Output nets */
wire t_4046,   t_4047,   t_4048;
/* u2_1380 Output nets */
wire t_4049,   t_4050,   t_4051;
/* u2_1381 Output nets */
wire t_4052,   t_4053,   t_4054;
/* u2_1382 Output nets */
wire t_4055,   t_4056,   t_4057;
/* u2_1383 Output nets */
wire t_4058,   t_4059,   t_4060;
/* u2_1384 Output nets */
wire t_4061,   t_4062,   t_4063;
/* u2_1385 Output nets */
wire t_4064,   t_4065,   t_4066;
/* u2_1386 Output nets */
wire t_4067,   t_4068,   t_4069;
/* u2_1387 Output nets */
wire t_4070,   t_4071,   t_4072;
/* u2_1388 Output nets */
wire t_4073,   t_4074,   t_4075;
/* u2_1389 Output nets */
wire t_4076,   t_4077,   t_4078;
/* u1_1390 Output nets */
wire t_4079,   t_4080;
/* u2_1391 Output nets */
wire t_4081,   t_4082,   t_4083;
/* u2_1392 Output nets */
wire t_4084,   t_4085,   t_4086;
/* u2_1393 Output nets */
wire t_4087,   t_4088,   t_4089;
/* u2_1394 Output nets */
wire t_4090,   t_4091,   t_4092;
/* u2_1395 Output nets */
wire t_4093,   t_4094,   t_4095;
/* u2_1396 Output nets */
wire t_4096,   t_4097,   t_4098;
/* u2_1397 Output nets */
wire t_4099,   t_4100,   t_4101;
/* u2_1398 Output nets */
wire t_4102,   t_4103,   t_4104;
/* u2_1399 Output nets */
wire t_4105,   t_4106,   t_4107;
/* u2_1400 Output nets */
wire t_4108,   t_4109,   t_4110;
/* u2_1401 Output nets */
wire t_4111,   t_4112,   t_4113;
/* u2_1402 Output nets */
wire t_4114,   t_4115,   t_4116;
/* u2_1403 Output nets */
wire t_4117,   t_4118,   t_4119;
/* u1_1404 Output nets */
wire t_4120,   t_4121;
/* u2_1405 Output nets */
wire t_4122,   t_4123,   t_4124;
/* u2_1406 Output nets */
wire t_4125,   t_4126,   t_4127;
/* u2_1407 Output nets */
wire t_4128,   t_4129,   t_4130;
/* u2_1408 Output nets */
wire t_4131,   t_4132,   t_4133;
/* u2_1409 Output nets */
wire t_4134,   t_4135,   t_4136;
/* u2_1410 Output nets */
wire t_4137,   t_4138,   t_4139;
/* u2_1411 Output nets */
wire t_4140,   t_4141,   t_4142;
/* u2_1412 Output nets */
wire t_4143,   t_4144,   t_4145;
/* u2_1413 Output nets */
wire t_4146,   t_4147,   t_4148;
/* u2_1414 Output nets */
wire t_4149,   t_4150,   t_4151;
/* u2_1415 Output nets */
wire t_4152,   t_4153,   t_4154;
/* u2_1416 Output nets */
wire t_4155,   t_4156,   t_4157;
/* u2_1417 Output nets */
wire t_4158,   t_4159,   t_4160;
/* u0_1418 Output nets */
wire t_4161,   t_4162;
/* u2_1419 Output nets */
wire t_4163,   t_4164,   t_4165;
/* u2_1420 Output nets */
wire t_4166,   t_4167,   t_4168;
/* u2_1421 Output nets */
wire t_4169,   t_4170,   t_4171;
/* u2_1422 Output nets */
wire t_4172,   t_4173,   t_4174;
/* u2_1423 Output nets */
wire t_4175,   t_4176,   t_4177;
/* u2_1424 Output nets */
wire t_4178,   t_4179,   t_4180;
/* u2_1425 Output nets */
wire t_4181,   t_4182,   t_4183;
/* u2_1426 Output nets */
wire t_4184,   t_4185,   t_4186;
/* u2_1427 Output nets */
wire t_4187,   t_4188,   t_4189;
/* u2_1428 Output nets */
wire t_4190,   t_4191,   t_4192;
/* u2_1429 Output nets */
wire t_4193,   t_4194,   t_4195;
/* u2_1430 Output nets */
wire t_4196,   t_4197,   t_4198;
/* u2_1431 Output nets */
wire t_4199,   t_4200,   t_4201;
/* u0_1432 Output nets */
wire t_4202,   t_4203;
/* u2_1433 Output nets */
wire t_4204,   t_4205,   t_4206;
/* u2_1434 Output nets */
wire t_4207,   t_4208,   t_4209;
/* u2_1435 Output nets */
wire t_4210,   t_4211,   t_4212;
/* u2_1436 Output nets */
wire t_4213,   t_4214,   t_4215;
/* u2_1437 Output nets */
wire t_4216,   t_4217,   t_4218;
/* u2_1438 Output nets */
wire t_4219,   t_4220,   t_4221;
/* u2_1439 Output nets */
wire t_4222,   t_4223,   t_4224;
/* u2_1440 Output nets */
wire t_4225,   t_4226,   t_4227;
/* u2_1441 Output nets */
wire t_4228,   t_4229,   t_4230;
/* u2_1442 Output nets */
wire t_4231,   t_4232,   t_4233;
/* u2_1443 Output nets */
wire t_4234,   t_4235,   t_4236;
/* u2_1444 Output nets */
wire t_4237,   t_4238,   t_4239;
/* u2_1445 Output nets */
wire t_4240,   t_4241,   t_4242;
/* u2_1446 Output nets */
wire t_4243,   t_4244,   t_4245;
/* u2_1447 Output nets */
wire t_4246,   t_4247,   t_4248;
/* u2_1448 Output nets */
wire t_4249,   t_4250,   t_4251;
/* u2_1449 Output nets */
wire t_4252,   t_4253,   t_4254;
/* u2_1450 Output nets */
wire t_4255,   t_4256,   t_4257;
/* u2_1451 Output nets */
wire t_4258,   t_4259,   t_4260;
/* u2_1452 Output nets */
wire t_4261,   t_4262,   t_4263;
/* u2_1453 Output nets */
wire t_4264,   t_4265,   t_4266;
/* u2_1454 Output nets */
wire t_4267,   t_4268,   t_4269;
/* u2_1455 Output nets */
wire t_4270,   t_4271,   t_4272;
/* u2_1456 Output nets */
wire t_4273,   t_4274,   t_4275;
/* u2_1457 Output nets */
wire t_4276,   t_4277,   t_4278;
/* u2_1458 Output nets */
wire t_4279,   t_4280,   t_4281;
/* u2_1459 Output nets */
wire t_4282,   t_4283,   t_4284;
/* u2_1460 Output nets */
wire t_4285,   t_4286,   t_4287;
/* u2_1461 Output nets */
wire t_4288,   t_4289,   t_4290;
/* u2_1462 Output nets */
wire t_4291,   t_4292,   t_4293;
/* u2_1463 Output nets */
wire t_4294,   t_4295,   t_4296;
/* u2_1464 Output nets */
wire t_4297,   t_4298,   t_4299;
/* u2_1465 Output nets */
wire t_4300,   t_4301,   t_4302;
/* u2_1466 Output nets */
wire t_4303,   t_4304,   t_4305;
/* u2_1467 Output nets */
wire t_4306,   t_4307,   t_4308;
/* u2_1468 Output nets */
wire t_4309,   t_4310,   t_4311;
/* u2_1469 Output nets */
wire t_4312,   t_4313,   t_4314;
/* u2_1470 Output nets */
wire t_4315,   t_4316,   t_4317;
/* u2_1471 Output nets */
wire t_4318,   t_4319,   t_4320;
/* u2_1472 Output nets */
wire t_4321,   t_4322,   t_4323;
/* u2_1473 Output nets */
wire t_4324,   t_4325,   t_4326;
/* u2_1474 Output nets */
wire t_4327,   t_4328,   t_4329;
/* u2_1475 Output nets */
wire t_4330,   t_4331,   t_4332;
/* u2_1476 Output nets */
wire t_4333,   t_4334,   t_4335;
/* u2_1477 Output nets */
wire t_4336,   t_4337,   t_4338;
/* u2_1478 Output nets */
wire t_4339,   t_4340,   t_4341;
/* u2_1479 Output nets */
wire t_4342,   t_4343,   t_4344;
/* u2_1480 Output nets */
wire t_4345,   t_4346,   t_4347;
/* u2_1481 Output nets */
wire t_4348,   t_4349,   t_4350;
/* u2_1482 Output nets */
wire t_4351,   t_4352,   t_4353;
/* u2_1483 Output nets */
wire t_4354,   t_4355,   t_4356;
/* u2_1484 Output nets */
wire t_4357,   t_4358,   t_4359;
/* u2_1485 Output nets */
wire t_4360,   t_4361,   t_4362;
/* u2_1486 Output nets */
wire t_4363,   t_4364,   t_4365;
/* u2_1487 Output nets */
wire t_4366,   t_4367,   t_4368;
/* u2_1488 Output nets */
wire t_4369,   t_4370,   t_4371;
/* u2_1489 Output nets */
wire t_4372,   t_4373,   t_4374;
/* u2_1490 Output nets */
wire t_4375,   t_4376,   t_4377;
/* u2_1491 Output nets */
wire t_4378,   t_4379,   t_4380;
/* u2_1492 Output nets */
wire t_4381,   t_4382,   t_4383;
/* u2_1493 Output nets */
wire t_4384,   t_4385,   t_4386;
/* u2_1494 Output nets */
wire t_4387,   t_4388,   t_4389;
/* u2_1495 Output nets */
wire t_4390,   t_4391,   t_4392;
/* u2_1496 Output nets */
wire t_4393,   t_4394,   t_4395;
/* u1_1497 Output nets */
wire t_4396,   t_4397;
/* u2_1498 Output nets */
wire t_4398,   t_4399,   t_4400;
/* u2_1499 Output nets */
wire t_4401,   t_4402,   t_4403;
/* u2_1500 Output nets */
wire t_4404,   t_4405,   t_4406;
/* u2_1501 Output nets */
wire t_4407,   t_4408,   t_4409;
/* u2_1502 Output nets */
wire t_4410,   t_4411,   t_4412;
/* u2_1503 Output nets */
wire t_4413,   t_4414,   t_4415;
/* u2_1504 Output nets */
wire t_4416,   t_4417,   t_4418;
/* u2_1505 Output nets */
wire t_4419,   t_4420,   t_4421;
/* u2_1506 Output nets */
wire t_4422,   t_4423,   t_4424;
/* u2_1507 Output nets */
wire t_4425,   t_4426,   t_4427;
/* u2_1508 Output nets */
wire t_4428,   t_4429,   t_4430;
/* u2_1509 Output nets */
wire t_4431,   t_4432,   t_4433;
/* u1_1510 Output nets */
wire t_4434,   t_4435;
/* u2_1511 Output nets */
wire t_4436,   t_4437,   t_4438;
/* u2_1512 Output nets */
wire t_4439,   t_4440,   t_4441;
/* u2_1513 Output nets */
wire t_4442,   t_4443,   t_4444;
/* u2_1514 Output nets */
wire t_4445,   t_4446,   t_4447;
/* u2_1515 Output nets */
wire t_4448,   t_4449,   t_4450;
/* u2_1516 Output nets */
wire t_4451,   t_4452,   t_4453;
/* u2_1517 Output nets */
wire t_4454,   t_4455,   t_4456;
/* u2_1518 Output nets */
wire t_4457,   t_4458,   t_4459;
/* u2_1519 Output nets */
wire t_4460,   t_4461,   t_4462;
/* u2_1520 Output nets */
wire t_4463,   t_4464,   t_4465;
/* u2_1521 Output nets */
wire t_4466,   t_4467,   t_4468;
/* u2_1522 Output nets */
wire t_4469,   t_4470,   t_4471;
/* u0_1523 Output nets */
wire t_4472,   t_4473;
/* u2_1524 Output nets */
wire t_4474,   t_4475,   t_4476;
/* u2_1525 Output nets */
wire t_4477,   t_4478,   t_4479;
/* u2_1526 Output nets */
wire t_4480,   t_4481,   t_4482;
/* u2_1527 Output nets */
wire t_4483,   t_4484,   t_4485;
/* u2_1528 Output nets */
wire t_4486,   t_4487,   t_4488;
/* u2_1529 Output nets */
wire t_4489,   t_4490,   t_4491;
/* u2_1530 Output nets */
wire t_4492,   t_4493,   t_4494;
/* u2_1531 Output nets */
wire t_4495,   t_4496,   t_4497;
/* u2_1532 Output nets */
wire t_4498,   t_4499,   t_4500;
/* u2_1533 Output nets */
wire t_4501,   t_4502,   t_4503;
/* u2_1534 Output nets */
wire t_4504,   t_4505,   t_4506;
/* u2_1535 Output nets */
wire t_4507,   t_4508,   t_4509;
/* u0_1536 Output nets */
wire t_4510,   t_4511;
/* u2_1537 Output nets */
wire t_4512,   t_4513,   t_4514;
/* u2_1538 Output nets */
wire t_4515,   t_4516,   t_4517;
/* u2_1539 Output nets */
wire t_4518,   t_4519,   t_4520;
/* u2_1540 Output nets */
wire t_4521,   t_4522,   t_4523;
/* u2_1541 Output nets */
wire t_4524,   t_4525,   t_4526;
/* u2_1542 Output nets */
wire t_4527,   t_4528,   t_4529;
/* u2_1543 Output nets */
wire t_4530,   t_4531,   t_4532;
/* u2_1544 Output nets */
wire t_4533,   t_4534,   t_4535;
/* u2_1545 Output nets */
wire t_4536,   t_4537,   t_4538;
/* u2_1546 Output nets */
wire t_4539,   t_4540,   t_4541;
/* u2_1547 Output nets */
wire t_4542,   t_4543,   t_4544;
/* u2_1548 Output nets */
wire t_4545,   t_4546,   t_4547;
/* u2_1549 Output nets */
wire t_4548,   t_4549,   t_4550;
/* u2_1550 Output nets */
wire t_4551,   t_4552,   t_4553;
/* u2_1551 Output nets */
wire t_4554,   t_4555,   t_4556;
/* u2_1552 Output nets */
wire t_4557,   t_4558,   t_4559;
/* u2_1553 Output nets */
wire t_4560,   t_4561,   t_4562;
/* u2_1554 Output nets */
wire t_4563,   t_4564,   t_4565;
/* u2_1555 Output nets */
wire t_4566,   t_4567,   t_4568;
/* u2_1556 Output nets */
wire t_4569,   t_4570,   t_4571;
/* u2_1557 Output nets */
wire t_4572,   t_4573,   t_4574;
/* u2_1558 Output nets */
wire t_4575,   t_4576,   t_4577;
/* u2_1559 Output nets */
wire t_4578,   t_4579,   t_4580;
/* u2_1560 Output nets */
wire t_4581,   t_4582,   t_4583;
/* u2_1561 Output nets */
wire t_4584,   t_4585,   t_4586;
/* u2_1562 Output nets */
wire t_4587,   t_4588,   t_4589;
/* u2_1563 Output nets */
wire t_4590,   t_4591,   t_4592;
/* u2_1564 Output nets */
wire t_4593,   t_4594,   t_4595;
/* u2_1565 Output nets */
wire t_4596,   t_4597,   t_4598;
/* u2_1566 Output nets */
wire t_4599,   t_4600,   t_4601;
/* u2_1567 Output nets */
wire t_4602,   t_4603,   t_4604;
/* u2_1568 Output nets */
wire t_4605,   t_4606,   t_4607;
/* u2_1569 Output nets */
wire t_4608,   t_4609,   t_4610;
/* u2_1570 Output nets */
wire t_4611,   t_4612,   t_4613;
/* u2_1571 Output nets */
wire t_4614,   t_4615,   t_4616;
/* u2_1572 Output nets */
wire t_4617,   t_4618,   t_4619;
/* u2_1573 Output nets */
wire t_4620,   t_4621,   t_4622;
/* u2_1574 Output nets */
wire t_4623,   t_4624,   t_4625;
/* u2_1575 Output nets */
wire t_4626,   t_4627,   t_4628;
/* u2_1576 Output nets */
wire t_4629,   t_4630,   t_4631;
/* u2_1577 Output nets */
wire t_4632,   t_4633,   t_4634;
/* u2_1578 Output nets */
wire t_4635,   t_4636,   t_4637;
/* u2_1579 Output nets */
wire t_4638,   t_4639,   t_4640;
/* u2_1580 Output nets */
wire t_4641,   t_4642,   t_4643;
/* u2_1581 Output nets */
wire t_4644,   t_4645,   t_4646;
/* u2_1582 Output nets */
wire t_4647,   t_4648,   t_4649;
/* u2_1583 Output nets */
wire t_4650,   t_4651,   t_4652;
/* u2_1584 Output nets */
wire t_4653,   t_4654,   t_4655;
/* u2_1585 Output nets */
wire t_4656,   t_4657,   t_4658;
/* u2_1586 Output nets */
wire t_4659,   t_4660,   t_4661;
/* u2_1587 Output nets */
wire t_4662,   t_4663,   t_4664;
/* u2_1588 Output nets */
wire t_4665,   t_4666,   t_4667;
/* u2_1589 Output nets */
wire t_4668,   t_4669,   t_4670;
/* u2_1590 Output nets */
wire t_4671,   t_4672,   t_4673;
/* u2_1591 Output nets */
wire t_4674,   t_4675,   t_4676;
/* u2_1592 Output nets */
wire t_4677,   t_4678,   t_4679;
/* u2_1593 Output nets */
wire t_4680,   t_4681,   t_4682;
/* u2_1594 Output nets */
wire t_4683,   t_4684,   t_4685;
/* u2_1595 Output nets */
wire t_4686,   t_4687,   t_4688;
/* u1_1596 Output nets */
wire t_4689,   t_4690;
/* u2_1597 Output nets */
wire t_4691,   t_4692,   t_4693;
/* u2_1598 Output nets */
wire t_4694,   t_4695,   t_4696;
/* u2_1599 Output nets */
wire t_4697,   t_4698,   t_4699;
/* u2_1600 Output nets */
wire t_4700,   t_4701,   t_4702;
/* u2_1601 Output nets */
wire t_4703,   t_4704,   t_4705;
/* u2_1602 Output nets */
wire t_4706,   t_4707,   t_4708;
/* u2_1603 Output nets */
wire t_4709,   t_4710,   t_4711;
/* u2_1604 Output nets */
wire t_4712,   t_4713,   t_4714;
/* u2_1605 Output nets */
wire t_4715,   t_4716,   t_4717;
/* u2_1606 Output nets */
wire t_4718,   t_4719,   t_4720;
/* u2_1607 Output nets */
wire t_4721,   t_4722,   t_4723;
/* u1_1608 Output nets */
wire t_4724,   t_4725;
/* u2_1609 Output nets */
wire t_4726,   t_4727,   t_4728;
/* u2_1610 Output nets */
wire t_4729,   t_4730,   t_4731;
/* u2_1611 Output nets */
wire t_4732,   t_4733,   t_4734;
/* u2_1612 Output nets */
wire t_4735,   t_4736,   t_4737;
/* u2_1613 Output nets */
wire t_4738,   t_4739,   t_4740;
/* u2_1614 Output nets */
wire t_4741,   t_4742,   t_4743;
/* u2_1615 Output nets */
wire t_4744,   t_4745,   t_4746;
/* u2_1616 Output nets */
wire t_4747,   t_4748,   t_4749;
/* u2_1617 Output nets */
wire t_4750,   t_4751,   t_4752;
/* u2_1618 Output nets */
wire t_4753,   t_4754,   t_4755;
/* u2_1619 Output nets */
wire t_4756,   t_4757,   t_4758;
/* u0_1620 Output nets */
wire t_4759,   t_4760;
/* u2_1621 Output nets */
wire t_4761,   t_4762,   t_4763;
/* u2_1622 Output nets */
wire t_4764,   t_4765,   t_4766;
/* u2_1623 Output nets */
wire t_4767,   t_4768,   t_4769;
/* u2_1624 Output nets */
wire t_4770,   t_4771,   t_4772;
/* u2_1625 Output nets */
wire t_4773,   t_4774,   t_4775;
/* u2_1626 Output nets */
wire t_4776,   t_4777,   t_4778;
/* u2_1627 Output nets */
wire t_4779,   t_4780,   t_4781;
/* u2_1628 Output nets */
wire t_4782,   t_4783,   t_4784;
/* u2_1629 Output nets */
wire t_4785,   t_4786,   t_4787;
/* u2_1630 Output nets */
wire t_4788,   t_4789,   t_4790;
/* u2_1631 Output nets */
wire t_4791,   t_4792,   t_4793;
/* u0_1632 Output nets */
wire t_4794,   t_4795;
/* u2_1633 Output nets */
wire t_4796,   t_4797,   t_4798;
/* u2_1634 Output nets */
wire t_4799,   t_4800,   t_4801;
/* u2_1635 Output nets */
wire t_4802,   t_4803,   t_4804;
/* u2_1636 Output nets */
wire t_4805,   t_4806,   t_4807;
/* u2_1637 Output nets */
wire t_4808,   t_4809,   t_4810;
/* u2_1638 Output nets */
wire t_4811,   t_4812,   t_4813;
/* u2_1639 Output nets */
wire t_4814,   t_4815,   t_4816;
/* u2_1640 Output nets */
wire t_4817,   t_4818,   t_4819;
/* u2_1641 Output nets */
wire t_4820,   t_4821,   t_4822;
/* u2_1642 Output nets */
wire t_4823,   t_4824,   t_4825;
/* u2_1643 Output nets */
wire t_4826,   t_4827,   t_4828;
/* u2_1644 Output nets */
wire t_4829,   t_4830,   t_4831;
/* u2_1645 Output nets */
wire t_4832,   t_4833,   t_4834;
/* u2_1646 Output nets */
wire t_4835,   t_4836,   t_4837;
/* u2_1647 Output nets */
wire t_4838,   t_4839,   t_4840;
/* u2_1648 Output nets */
wire t_4841,   t_4842,   t_4843;
/* u2_1649 Output nets */
wire t_4844,   t_4845,   t_4846;
/* u2_1650 Output nets */
wire t_4847,   t_4848,   t_4849;
/* u2_1651 Output nets */
wire t_4850,   t_4851,   t_4852;
/* u2_1652 Output nets */
wire t_4853,   t_4854,   t_4855;
/* u2_1653 Output nets */
wire t_4856,   t_4857,   t_4858;
/* u2_1654 Output nets */
wire t_4859,   t_4860,   t_4861;
/* u2_1655 Output nets */
wire t_4862,   t_4863,   t_4864;
/* u2_1656 Output nets */
wire t_4865,   t_4866,   t_4867;
/* u2_1657 Output nets */
wire t_4868,   t_4869,   t_4870;
/* u2_1658 Output nets */
wire t_4871,   t_4872,   t_4873;
/* u2_1659 Output nets */
wire t_4874,   t_4875,   t_4876;
/* u2_1660 Output nets */
wire t_4877,   t_4878,   t_4879;
/* u2_1661 Output nets */
wire t_4880,   t_4881,   t_4882;
/* u2_1662 Output nets */
wire t_4883,   t_4884,   t_4885;
/* u2_1663 Output nets */
wire t_4886,   t_4887,   t_4888;
/* u2_1664 Output nets */
wire t_4889,   t_4890,   t_4891;
/* u2_1665 Output nets */
wire t_4892,   t_4893,   t_4894;
/* u2_1666 Output nets */
wire t_4895,   t_4896,   t_4897;
/* u2_1667 Output nets */
wire t_4898,   t_4899,   t_4900;
/* u2_1668 Output nets */
wire t_4901,   t_4902,   t_4903;
/* u2_1669 Output nets */
wire t_4904,   t_4905,   t_4906;
/* u2_1670 Output nets */
wire t_4907,   t_4908,   t_4909;
/* u2_1671 Output nets */
wire t_4910,   t_4911,   t_4912;
/* u2_1672 Output nets */
wire t_4913,   t_4914,   t_4915;
/* u2_1673 Output nets */
wire t_4916,   t_4917,   t_4918;
/* u2_1674 Output nets */
wire t_4919,   t_4920,   t_4921;
/* u2_1675 Output nets */
wire t_4922,   t_4923,   t_4924;
/* u2_1676 Output nets */
wire t_4925,   t_4926,   t_4927;
/* u2_1677 Output nets */
wire t_4928,   t_4929,   t_4930;
/* u2_1678 Output nets */
wire t_4931,   t_4932,   t_4933;
/* u2_1679 Output nets */
wire t_4934,   t_4935,   t_4936;
/* u2_1680 Output nets */
wire t_4937,   t_4938,   t_4939;
/* u2_1681 Output nets */
wire t_4940,   t_4941,   t_4942;
/* u2_1682 Output nets */
wire t_4943,   t_4944,   t_4945;
/* u2_1683 Output nets */
wire t_4946,   t_4947,   t_4948;
/* u2_1684 Output nets */
wire t_4949,   t_4950,   t_4951;
/* u2_1685 Output nets */
wire t_4952,   t_4953,   t_4954;
/* u2_1686 Output nets */
wire t_4955,   t_4956,   t_4957;
/* u1_1687 Output nets */
wire t_4958,   t_4959;
/* u2_1688 Output nets */
wire t_4960,   t_4961,   t_4962;
/* u2_1689 Output nets */
wire t_4963,   t_4964,   t_4965;
/* u2_1690 Output nets */
wire t_4966,   t_4967,   t_4968;
/* u2_1691 Output nets */
wire t_4969,   t_4970,   t_4971;
/* u2_1692 Output nets */
wire t_4972,   t_4973,   t_4974;
/* u2_1693 Output nets */
wire t_4975,   t_4976,   t_4977;
/* u2_1694 Output nets */
wire t_4978,   t_4979,   t_4980;
/* u2_1695 Output nets */
wire t_4981,   t_4982,   t_4983;
/* u2_1696 Output nets */
wire t_4984,   t_4985,   t_4986;
/* u2_1697 Output nets */
wire t_4987,   t_4988,   t_4989;
/* u1_1698 Output nets */
wire t_4990,   t_4991;
/* u2_1699 Output nets */
wire t_4992,   t_4993,   t_4994;
/* u2_1700 Output nets */
wire t_4995,   t_4996,   t_4997;
/* u2_1701 Output nets */
wire t_4998,   t_4999,   t_5000;
/* u2_1702 Output nets */
wire t_5001,   t_5002,   t_5003;
/* u2_1703 Output nets */
wire t_5004,   t_5005,   t_5006;
/* u2_1704 Output nets */
wire t_5007,   t_5008,   t_5009;
/* u2_1705 Output nets */
wire t_5010,   t_5011,   t_5012;
/* u2_1706 Output nets */
wire t_5013,   t_5014,   t_5015;
/* u2_1707 Output nets */
wire t_5016,   t_5017,   t_5018;
/* u2_1708 Output nets */
wire t_5019,   t_5020,   t_5021;
/* u0_1709 Output nets */
wire t_5022,   t_5023;
/* u2_1710 Output nets */
wire t_5024,   t_5025,   t_5026;
/* u2_1711 Output nets */
wire t_5027,   t_5028,   t_5029;
/* u2_1712 Output nets */
wire t_5030,   t_5031,   t_5032;
/* u2_1713 Output nets */
wire t_5033,   t_5034,   t_5035;
/* u2_1714 Output nets */
wire t_5036,   t_5037,   t_5038;
/* u2_1715 Output nets */
wire t_5039,   t_5040,   t_5041;
/* u2_1716 Output nets */
wire t_5042,   t_5043,   t_5044;
/* u2_1717 Output nets */
wire t_5045,   t_5046,   t_5047;
/* u2_1718 Output nets */
wire t_5048,   t_5049,   t_5050;
/* u2_1719 Output nets */
wire t_5051,   t_5052,   t_5053;
/* u0_1720 Output nets */
wire t_5054,   t_5055;
/* u2_1721 Output nets */
wire t_5056,   t_5057,   t_5058;
/* u2_1722 Output nets */
wire t_5059,   t_5060,   t_5061;
/* u2_1723 Output nets */
wire t_5062,   t_5063,   t_5064;
/* u2_1724 Output nets */
wire t_5065,   t_5066,   t_5067;
/* u2_1725 Output nets */
wire t_5068,   t_5069,   t_5070;
/* u2_1726 Output nets */
wire t_5071,   t_5072,   t_5073;
/* u2_1727 Output nets */
wire t_5074,   t_5075,   t_5076;
/* u2_1728 Output nets */
wire t_5077,   t_5078,   t_5079;
/* u2_1729 Output nets */
wire t_5080,   t_5081,   t_5082;
/* u2_1730 Output nets */
wire t_5083,   t_5084,   t_5085;
/* u2_1731 Output nets */
wire t_5086,   t_5087,   t_5088;
/* u2_1732 Output nets */
wire t_5089,   t_5090,   t_5091;
/* u2_1733 Output nets */
wire t_5092,   t_5093,   t_5094;
/* u2_1734 Output nets */
wire t_5095,   t_5096,   t_5097;
/* u2_1735 Output nets */
wire t_5098,   t_5099,   t_5100;
/* u2_1736 Output nets */
wire t_5101,   t_5102,   t_5103;
/* u2_1737 Output nets */
wire t_5104,   t_5105,   t_5106;
/* u2_1738 Output nets */
wire t_5107,   t_5108,   t_5109;
/* u2_1739 Output nets */
wire t_5110,   t_5111,   t_5112;
/* u2_1740 Output nets */
wire t_5113,   t_5114,   t_5115;
/* u2_1741 Output nets */
wire t_5116,   t_5117,   t_5118;
/* u2_1742 Output nets */
wire t_5119,   t_5120,   t_5121;
/* u2_1743 Output nets */
wire t_5122,   t_5123,   t_5124;
/* u2_1744 Output nets */
wire t_5125,   t_5126,   t_5127;
/* u2_1745 Output nets */
wire t_5128,   t_5129,   t_5130;
/* u2_1746 Output nets */
wire t_5131,   t_5132,   t_5133;
/* u2_1747 Output nets */
wire t_5134,   t_5135,   t_5136;
/* u2_1748 Output nets */
wire t_5137,   t_5138,   t_5139;
/* u2_1749 Output nets */
wire t_5140,   t_5141,   t_5142;
/* u2_1750 Output nets */
wire t_5143,   t_5144,   t_5145;
/* u2_1751 Output nets */
wire t_5146,   t_5147,   t_5148;
/* u2_1752 Output nets */
wire t_5149,   t_5150,   t_5151;
/* u2_1753 Output nets */
wire t_5152,   t_5153,   t_5154;
/* u2_1754 Output nets */
wire t_5155,   t_5156,   t_5157;
/* u2_1755 Output nets */
wire t_5158,   t_5159,   t_5160;
/* u2_1756 Output nets */
wire t_5161,   t_5162,   t_5163;
/* u2_1757 Output nets */
wire t_5164,   t_5165,   t_5166;
/* u2_1758 Output nets */
wire t_5167,   t_5168,   t_5169;
/* u2_1759 Output nets */
wire t_5170,   t_5171,   t_5172;
/* u2_1760 Output nets */
wire t_5173,   t_5174,   t_5175;
/* u2_1761 Output nets */
wire t_5176,   t_5177,   t_5178;
/* u2_1762 Output nets */
wire t_5179,   t_5180,   t_5181;
/* u2_1763 Output nets */
wire t_5182,   t_5183,   t_5184;
/* u2_1764 Output nets */
wire t_5185,   t_5186,   t_5187;
/* u2_1765 Output nets */
wire t_5188,   t_5189,   t_5190;
/* u2_1766 Output nets */
wire t_5191,   t_5192,   t_5193;
/* u2_1767 Output nets */
wire t_5194,   t_5195,   t_5196;
/* u2_1768 Output nets */
wire t_5197,   t_5198,   t_5199;
/* u2_1769 Output nets */
wire t_5200,   t_5201,   t_5202;
/* u1_1770 Output nets */
wire t_5203,   t_5204;
/* u2_1771 Output nets */
wire t_5205,   t_5206,   t_5207;
/* u2_1772 Output nets */
wire t_5208,   t_5209,   t_5210;
/* u2_1773 Output nets */
wire t_5211,   t_5212,   t_5213;
/* u2_1774 Output nets */
wire t_5214,   t_5215,   t_5216;
/* u2_1775 Output nets */
wire t_5217,   t_5218,   t_5219;
/* u2_1776 Output nets */
wire t_5220,   t_5221,   t_5222;
/* u2_1777 Output nets */
wire t_5223,   t_5224,   t_5225;
/* u2_1778 Output nets */
wire t_5226,   t_5227,   t_5228;
/* u2_1779 Output nets */
wire t_5229,   t_5230,   t_5231;
/* u1_1780 Output nets */
wire t_5232,   t_5233;
/* u2_1781 Output nets */
wire t_5234,   t_5235,   t_5236;
/* u2_1782 Output nets */
wire t_5237,   t_5238,   t_5239;
/* u2_1783 Output nets */
wire t_5240,   t_5241,   t_5242;
/* u2_1784 Output nets */
wire t_5243,   t_5244,   t_5245;
/* u2_1785 Output nets */
wire t_5246,   t_5247,   t_5248;
/* u2_1786 Output nets */
wire t_5249,   t_5250,   t_5251;
/* u2_1787 Output nets */
wire t_5252,   t_5253,   t_5254;
/* u2_1788 Output nets */
wire t_5255,   t_5256,   t_5257;
/* u2_1789 Output nets */
wire t_5258,   t_5259,   t_5260;
/* u0_1790 Output nets */
wire t_5261,   t_5262;
/* u2_1791 Output nets */
wire t_5263,   t_5264,   t_5265;
/* u2_1792 Output nets */
wire t_5266,   t_5267,   t_5268;
/* u2_1793 Output nets */
wire t_5269,   t_5270,   t_5271;
/* u2_1794 Output nets */
wire t_5272,   t_5273,   t_5274;
/* u2_1795 Output nets */
wire t_5275,   t_5276,   t_5277;
/* u2_1796 Output nets */
wire t_5278,   t_5279,   t_5280;
/* u2_1797 Output nets */
wire t_5281,   t_5282,   t_5283;
/* u2_1798 Output nets */
wire t_5284,   t_5285,   t_5286;
/* u2_1799 Output nets */
wire t_5287,   t_5288,   t_5289;
/* u0_1800 Output nets */
wire t_5290,   t_5291;
/* u2_1801 Output nets */
wire t_5292,   t_5293,   t_5294;
/* u2_1802 Output nets */
wire t_5295,   t_5296,   t_5297;
/* u2_1803 Output nets */
wire t_5298,   t_5299,   t_5300;
/* u2_1804 Output nets */
wire t_5301,   t_5302,   t_5303;
/* u2_1805 Output nets */
wire t_5304,   t_5305,   t_5306;
/* u2_1806 Output nets */
wire t_5307,   t_5308,   t_5309;
/* u2_1807 Output nets */
wire t_5310,   t_5311,   t_5312;
/* u2_1808 Output nets */
wire t_5313,   t_5314,   t_5315;
/* u2_1809 Output nets */
wire t_5316,   t_5317,   t_5318;
/* u2_1810 Output nets */
wire t_5319,   t_5320,   t_5321;
/* u2_1811 Output nets */
wire t_5322,   t_5323,   t_5324;
/* u2_1812 Output nets */
wire t_5325,   t_5326,   t_5327;
/* u2_1813 Output nets */
wire t_5328,   t_5329,   t_5330;
/* u2_1814 Output nets */
wire t_5331,   t_5332,   t_5333;
/* u2_1815 Output nets */
wire t_5334,   t_5335,   t_5336;
/* u2_1816 Output nets */
wire t_5337,   t_5338,   t_5339;
/* u2_1817 Output nets */
wire t_5340,   t_5341,   t_5342;
/* u2_1818 Output nets */
wire t_5343,   t_5344,   t_5345;
/* u2_1819 Output nets */
wire t_5346,   t_5347,   t_5348;
/* u2_1820 Output nets */
wire t_5349,   t_5350,   t_5351;
/* u2_1821 Output nets */
wire t_5352,   t_5353,   t_5354;
/* u2_1822 Output nets */
wire t_5355,   t_5356,   t_5357;
/* u2_1823 Output nets */
wire t_5358,   t_5359,   t_5360;
/* u2_1824 Output nets */
wire t_5361,   t_5362,   t_5363;
/* u2_1825 Output nets */
wire t_5364,   t_5365,   t_5366;
/* u2_1826 Output nets */
wire t_5367,   t_5368,   t_5369;
/* u2_1827 Output nets */
wire t_5370,   t_5371,   t_5372;
/* u2_1828 Output nets */
wire t_5373,   t_5374,   t_5375;
/* u2_1829 Output nets */
wire t_5376,   t_5377,   t_5378;
/* u2_1830 Output nets */
wire t_5379,   t_5380,   t_5381;
/* u2_1831 Output nets */
wire t_5382,   t_5383,   t_5384;
/* u2_1832 Output nets */
wire t_5385,   t_5386,   t_5387;
/* u2_1833 Output nets */
wire t_5388,   t_5389,   t_5390;
/* u2_1834 Output nets */
wire t_5391,   t_5392,   t_5393;
/* u2_1835 Output nets */
wire t_5394,   t_5395,   t_5396;
/* u2_1836 Output nets */
wire t_5397,   t_5398,   t_5399;
/* u2_1837 Output nets */
wire t_5400,   t_5401,   t_5402;
/* u2_1838 Output nets */
wire t_5403,   t_5404,   t_5405;
/* u2_1839 Output nets */
wire t_5406,   t_5407,   t_5408;
/* u2_1840 Output nets */
wire t_5409,   t_5410,   t_5411;
/* u2_1841 Output nets */
wire t_5412,   t_5413,   t_5414;
/* u2_1842 Output nets */
wire t_5415,   t_5416,   t_5417;
/* u2_1843 Output nets */
wire t_5418,   t_5419,   t_5420;
/* u2_1844 Output nets */
wire t_5421,   t_5422,   t_5423;
/* u1_1845 Output nets */
wire t_5424,   t_5425;
/* u2_1846 Output nets */
wire t_5426,   t_5427,   t_5428;
/* u2_1847 Output nets */
wire t_5429,   t_5430,   t_5431;
/* u2_1848 Output nets */
wire t_5432,   t_5433,   t_5434;
/* u2_1849 Output nets */
wire t_5435,   t_5436,   t_5437;
/* u2_1850 Output nets */
wire t_5438,   t_5439,   t_5440;
/* u2_1851 Output nets */
wire t_5441,   t_5442,   t_5443;
/* u2_1852 Output nets */
wire t_5444,   t_5445,   t_5446;
/* u2_1853 Output nets */
wire t_5447,   t_5448,   t_5449;
/* u1_1854 Output nets */
wire t_5450,   t_5451;
/* u2_1855 Output nets */
wire t_5452,   t_5453,   t_5454;
/* u2_1856 Output nets */
wire t_5455,   t_5456,   t_5457;
/* u2_1857 Output nets */
wire t_5458,   t_5459,   t_5460;
/* u2_1858 Output nets */
wire t_5461,   t_5462,   t_5463;
/* u2_1859 Output nets */
wire t_5464,   t_5465,   t_5466;
/* u2_1860 Output nets */
wire t_5467,   t_5468,   t_5469;
/* u2_1861 Output nets */
wire t_5470,   t_5471,   t_5472;
/* u2_1862 Output nets */
wire t_5473,   t_5474,   t_5475;
/* u0_1863 Output nets */
wire t_5476,   t_5477;
/* u2_1864 Output nets */
wire t_5478,   t_5479,   t_5480;
/* u2_1865 Output nets */
wire t_5481,   t_5482,   t_5483;
/* u2_1866 Output nets */
wire t_5484,   t_5485,   t_5486;
/* u2_1867 Output nets */
wire t_5487,   t_5488,   t_5489;
/* u2_1868 Output nets */
wire t_5490,   t_5491,   t_5492;
/* u2_1869 Output nets */
wire t_5493,   t_5494,   t_5495;
/* u2_1870 Output nets */
wire t_5496,   t_5497,   t_5498;
/* u2_1871 Output nets */
wire t_5499,   t_5500,   t_5501;
/* u0_1872 Output nets */
wire t_5502,   t_5503;
/* u2_1873 Output nets */
wire t_5504,   t_5505,   t_5506;
/* u2_1874 Output nets */
wire t_5507,   t_5508,   t_5509;
/* u2_1875 Output nets */
wire t_5510,   t_5511,   t_5512;
/* u2_1876 Output nets */
wire t_5513,   t_5514,   t_5515;
/* u2_1877 Output nets */
wire t_5516,   t_5517,   t_5518;
/* u2_1878 Output nets */
wire t_5519,   t_5520,   t_5521;
/* u2_1879 Output nets */
wire t_5522,   t_5523,   t_5524;
/* u2_1880 Output nets */
wire t_5525,   t_5526,   t_5527;
/* u2_1881 Output nets */
wire t_5528,   t_5529,   t_5530;
/* u2_1882 Output nets */
wire t_5531,   t_5532,   t_5533;
/* u2_1883 Output nets */
wire t_5534,   t_5535,   t_5536;
/* u2_1884 Output nets */
wire t_5537,   t_5538,   t_5539;
/* u2_1885 Output nets */
wire t_5540,   t_5541,   t_5542;
/* u2_1886 Output nets */
wire t_5543,   t_5544,   t_5545;
/* u2_1887 Output nets */
wire t_5546,   t_5547,   t_5548;
/* u2_1888 Output nets */
wire t_5549,   t_5550,   t_5551;
/* u2_1889 Output nets */
wire t_5552,   t_5553,   t_5554;
/* u2_1890 Output nets */
wire t_5555,   t_5556,   t_5557;
/* u2_1891 Output nets */
wire t_5558,   t_5559,   t_5560;
/* u2_1892 Output nets */
wire t_5561,   t_5562,   t_5563;
/* u2_1893 Output nets */
wire t_5564,   t_5565,   t_5566;
/* u2_1894 Output nets */
wire t_5567,   t_5568,   t_5569;
/* u2_1895 Output nets */
wire t_5570,   t_5571,   t_5572;
/* u2_1896 Output nets */
wire t_5573,   t_5574,   t_5575;
/* u2_1897 Output nets */
wire t_5576,   t_5577,   t_5578;
/* u2_1898 Output nets */
wire t_5579,   t_5580,   t_5581;
/* u2_1899 Output nets */
wire t_5582,   t_5583,   t_5584;
/* u2_1900 Output nets */
wire t_5585,   t_5586,   t_5587;
/* u2_1901 Output nets */
wire t_5588,   t_5589,   t_5590;
/* u2_1902 Output nets */
wire t_5591,   t_5592,   t_5593;
/* u2_1903 Output nets */
wire t_5594,   t_5595,   t_5596;
/* u2_1904 Output nets */
wire t_5597,   t_5598,   t_5599;
/* u2_1905 Output nets */
wire t_5600,   t_5601,   t_5602;
/* u2_1906 Output nets */
wire t_5603,   t_5604,   t_5605;
/* u2_1907 Output nets */
wire t_5606,   t_5607,   t_5608;
/* u2_1908 Output nets */
wire t_5609,   t_5610,   t_5611;
/* u2_1909 Output nets */
wire t_5612,   t_5613,   t_5614;
/* u2_1910 Output nets */
wire t_5615,   t_5616,   t_5617;
/* u2_1911 Output nets */
wire t_5618,   t_5619,   t_5620;
/* u1_1912 Output nets */
wire t_5621,   t_5622;
/* u2_1913 Output nets */
wire t_5623,   t_5624,   t_5625;
/* u2_1914 Output nets */
wire t_5626,   t_5627,   t_5628;
/* u2_1915 Output nets */
wire t_5629,   t_5630,   t_5631;
/* u2_1916 Output nets */
wire t_5632,   t_5633,   t_5634;
/* u2_1917 Output nets */
wire t_5635,   t_5636,   t_5637;
/* u2_1918 Output nets */
wire t_5638,   t_5639,   t_5640;
/* u2_1919 Output nets */
wire t_5641,   t_5642,   t_5643;
/* u1_1920 Output nets */
wire t_5644,   t_5645;
/* u2_1921 Output nets */
wire t_5646,   t_5647,   t_5648;
/* u2_1922 Output nets */
wire t_5649,   t_5650,   t_5651;
/* u2_1923 Output nets */
wire t_5652,   t_5653,   t_5654;
/* u2_1924 Output nets */
wire t_5655,   t_5656,   t_5657;
/* u2_1925 Output nets */
wire t_5658,   t_5659,   t_5660;
/* u2_1926 Output nets */
wire t_5661,   t_5662,   t_5663;
/* u2_1927 Output nets */
wire t_5664,   t_5665,   t_5666;
/* u0_1928 Output nets */
wire t_5667,   t_5668;
/* u2_1929 Output nets */
wire t_5669,   t_5670,   t_5671;
/* u2_1930 Output nets */
wire t_5672,   t_5673,   t_5674;
/* u2_1931 Output nets */
wire t_5675,   t_5676,   t_5677;
/* u2_1932 Output nets */
wire t_5678,   t_5679,   t_5680;
/* u2_1933 Output nets */
wire t_5681,   t_5682,   t_5683;
/* u2_1934 Output nets */
wire t_5684,   t_5685,   t_5686;
/* u2_1935 Output nets */
wire t_5687,   t_5688,   t_5689;
/* u0_1936 Output nets */
wire t_5690,   t_5691;
/* u2_1937 Output nets */
wire t_5692,   t_5693,   t_5694;
/* u2_1938 Output nets */
wire t_5695,   t_5696,   t_5697;
/* u2_1939 Output nets */
wire t_5698,   t_5699,   t_5700;
/* u2_1940 Output nets */
wire t_5701,   t_5702,   t_5703;
/* u2_1941 Output nets */
wire t_5704,   t_5705,   t_5706;
/* u2_1942 Output nets */
wire t_5707,   t_5708,   t_5709;
/* u2_1943 Output nets */
wire t_5710,   t_5711,   t_5712;
/* u2_1944 Output nets */
wire t_5713,   t_5714,   t_5715;
/* u2_1945 Output nets */
wire t_5716,   t_5717,   t_5718;
/* u2_1946 Output nets */
wire t_5719,   t_5720,   t_5721;
/* u2_1947 Output nets */
wire t_5722,   t_5723,   t_5724;
/* u2_1948 Output nets */
wire t_5725,   t_5726,   t_5727;
/* u2_1949 Output nets */
wire t_5728,   t_5729,   t_5730;
/* u2_1950 Output nets */
wire t_5731,   t_5732,   t_5733;
/* u2_1951 Output nets */
wire t_5734,   t_5735,   t_5736;
/* u2_1952 Output nets */
wire t_5737,   t_5738,   t_5739;
/* u2_1953 Output nets */
wire t_5740,   t_5741,   t_5742;
/* u2_1954 Output nets */
wire t_5743,   t_5744,   t_5745;
/* u2_1955 Output nets */
wire t_5746,   t_5747,   t_5748;
/* u2_1956 Output nets */
wire t_5749,   t_5750,   t_5751;
/* u2_1957 Output nets */
wire t_5752,   t_5753,   t_5754;
/* u2_1958 Output nets */
wire t_5755,   t_5756,   t_5757;
/* u2_1959 Output nets */
wire t_5758,   t_5759,   t_5760;
/* u2_1960 Output nets */
wire t_5761,   t_5762,   t_5763;
/* u2_1961 Output nets */
wire t_5764,   t_5765,   t_5766;
/* u2_1962 Output nets */
wire t_5767,   t_5768,   t_5769;
/* u2_1963 Output nets */
wire t_5770,   t_5771,   t_5772;
/* u2_1964 Output nets */
wire t_5773,   t_5774,   t_5775;
/* u2_1965 Output nets */
wire t_5776,   t_5777,   t_5778;
/* u2_1966 Output nets */
wire t_5779,   t_5780,   t_5781;
/* u2_1967 Output nets */
wire t_5782,   t_5783,   t_5784;
/* u2_1968 Output nets */
wire t_5785,   t_5786,   t_5787;
/* u2_1969 Output nets */
wire t_5788,   t_5789,   t_5790;
/* u2_1970 Output nets */
wire t_5791,   t_5792,   t_5793;
/* u1_1971 Output nets */
wire t_5794,   t_5795;
/* u2_1972 Output nets */
wire t_5796,   t_5797,   t_5798;
/* u2_1973 Output nets */
wire t_5799,   t_5800,   t_5801;
/* u2_1974 Output nets */
wire t_5802,   t_5803,   t_5804;
/* u2_1975 Output nets */
wire t_5805,   t_5806,   t_5807;
/* u2_1976 Output nets */
wire t_5808,   t_5809,   t_5810;
/* u2_1977 Output nets */
wire t_5811,   t_5812,   t_5813;
/* u1_1978 Output nets */
wire t_5814,   t_5815;
/* u2_1979 Output nets */
wire t_5816,   t_5817,   t_5818;
/* u2_1980 Output nets */
wire t_5819,   t_5820,   t_5821;
/* u2_1981 Output nets */
wire t_5822,   t_5823,   t_5824;
/* u2_1982 Output nets */
wire t_5825,   t_5826,   t_5827;
/* u2_1983 Output nets */
wire t_5828,   t_5829,   t_5830;
/* u2_1984 Output nets */
wire t_5831,   t_5832,   t_5833;
/* u0_1985 Output nets */
wire t_5834,   t_5835;
/* u2_1986 Output nets */
wire t_5836,   t_5837,   t_5838;
/* u2_1987 Output nets */
wire t_5839,   t_5840,   t_5841;
/* u2_1988 Output nets */
wire t_5842,   t_5843,   t_5844;
/* u2_1989 Output nets */
wire t_5845,   t_5846,   t_5847;
/* u2_1990 Output nets */
wire t_5848,   t_5849,   t_5850;
/* u2_1991 Output nets */
wire t_5851,   t_5852,   t_5853;
/* u0_1992 Output nets */
wire t_5854,   t_5855;
/* u2_1993 Output nets */
wire t_5856,   t_5857,   t_5858;
/* u2_1994 Output nets */
wire t_5859,   t_5860,   t_5861;
/* u2_1995 Output nets */
wire t_5862,   t_5863,   t_5864;
/* u2_1996 Output nets */
wire t_5865,   t_5866,   t_5867;
/* u2_1997 Output nets */
wire t_5868,   t_5869,   t_5870;
/* u2_1998 Output nets */
wire t_5871,   t_5872,   t_5873;
/* u2_1999 Output nets */
wire t_5874,   t_5875,   t_5876;
/* u2_2000 Output nets */
wire t_5877,   t_5878,   t_5879;
/* u2_2001 Output nets */
wire t_5880,   t_5881,   t_5882;
/* u2_2002 Output nets */
wire t_5883,   t_5884,   t_5885;
/* u2_2003 Output nets */
wire t_5886,   t_5887,   t_5888;
/* u2_2004 Output nets */
wire t_5889,   t_5890,   t_5891;
/* u2_2005 Output nets */
wire t_5892,   t_5893,   t_5894;
/* u2_2006 Output nets */
wire t_5895,   t_5896,   t_5897;
/* u2_2007 Output nets */
wire t_5898,   t_5899,   t_5900;
/* u2_2008 Output nets */
wire t_5901,   t_5902,   t_5903;
/* u2_2009 Output nets */
wire t_5904,   t_5905,   t_5906;
/* u2_2010 Output nets */
wire t_5907,   t_5908,   t_5909;
/* u2_2011 Output nets */
wire t_5910,   t_5911,   t_5912;
/* u2_2012 Output nets */
wire t_5913,   t_5914,   t_5915;
/* u2_2013 Output nets */
wire t_5916,   t_5917,   t_5918;
/* u2_2014 Output nets */
wire t_5919,   t_5920,   t_5921;
/* u2_2015 Output nets */
wire t_5922,   t_5923,   t_5924;
/* u2_2016 Output nets */
wire t_5925,   t_5926,   t_5927;
/* u2_2017 Output nets */
wire t_5928,   t_5929,   t_5930;
/* u2_2018 Output nets */
wire t_5931,   t_5932,   t_5933;
/* u2_2019 Output nets */
wire t_5934,   t_5935,   t_5936;
/* u2_2020 Output nets */
wire t_5937,   t_5938,   t_5939;
/* u2_2021 Output nets */
wire t_5940,   t_5941,   t_5942;
/* u1_2022 Output nets */
wire t_5943,   t_5944;
/* u2_2023 Output nets */
wire t_5945,   t_5946,   t_5947;
/* u2_2024 Output nets */
wire t_5948,   t_5949,   t_5950;
/* u2_2025 Output nets */
wire t_5951,   t_5952,   t_5953;
/* u2_2026 Output nets */
wire t_5954,   t_5955,   t_5956;
/* u2_2027 Output nets */
wire t_5957,   t_5958,   t_5959;
/* u1_2028 Output nets */
wire t_5960,   t_5961;
/* u2_2029 Output nets */
wire t_5962,   t_5963,   t_5964;
/* u2_2030 Output nets */
wire t_5965,   t_5966,   t_5967;
/* u2_2031 Output nets */
wire t_5968,   t_5969,   t_5970;
/* u2_2032 Output nets */
wire t_5971,   t_5972,   t_5973;
/* u2_2033 Output nets */
wire t_5974,   t_5975,   t_5976;
/* u0_2034 Output nets */
wire t_5977,   t_5978;
/* u2_2035 Output nets */
wire t_5979,   t_5980,   t_5981;
/* u2_2036 Output nets */
wire t_5982,   t_5983,   t_5984;
/* u2_2037 Output nets */
wire t_5985,   t_5986,   t_5987;
/* u2_2038 Output nets */
wire t_5988,   t_5989,   t_5990;
/* u2_2039 Output nets */
wire t_5991,   t_5992,   t_5993;
/* u0_2040 Output nets */
wire t_5994,   t_5995;
/* u2_2041 Output nets */
wire t_5996,   t_5997,   t_5998;
/* u2_2042 Output nets */
wire t_5999,   t_6000,   t_6001;
/* u2_2043 Output nets */
wire t_6002,   t_6003,   t_6004;
/* u2_2044 Output nets */
wire t_6005,   t_6006,   t_6007;
/* u2_2045 Output nets */
wire t_6008,   t_6009,   t_6010;
/* u2_2046 Output nets */
wire t_6011,   t_6012,   t_6013;
/* u2_2047 Output nets */
wire t_6014,   t_6015,   t_6016;
/* u2_2048 Output nets */
wire t_6017,   t_6018,   t_6019;
/* u2_2049 Output nets */
wire t_6020,   t_6021,   t_6022;
/* u2_2050 Output nets */
wire t_6023,   t_6024,   t_6025;
/* u2_2051 Output nets */
wire t_6026,   t_6027,   t_6028;
/* u2_2052 Output nets */
wire t_6029,   t_6030,   t_6031;
/* u2_2053 Output nets */
wire t_6032,   t_6033,   t_6034;
/* u2_2054 Output nets */
wire t_6035,   t_6036,   t_6037;
/* u2_2055 Output nets */
wire t_6038,   t_6039,   t_6040;
/* u2_2056 Output nets */
wire t_6041,   t_6042,   t_6043;
/* u2_2057 Output nets */
wire t_6044,   t_6045,   t_6046;
/* u2_2058 Output nets */
wire t_6047,   t_6048,   t_6049;
/* u2_2059 Output nets */
wire t_6050,   t_6051,   t_6052;
/* u2_2060 Output nets */
wire t_6053,   t_6054,   t_6055;
/* u2_2061 Output nets */
wire t_6056,   t_6057,   t_6058;
/* u2_2062 Output nets */
wire t_6059,   t_6060,   t_6061;
/* u2_2063 Output nets */
wire t_6062,   t_6063,   t_6064;
/* u2_2064 Output nets */
wire t_6065,   t_6066,   t_6067;
/* u1_2065 Output nets */
wire t_6068,   t_6069;
/* u2_2066 Output nets */
wire t_6070,   t_6071,   t_6072;
/* u2_2067 Output nets */
wire t_6073,   t_6074,   t_6075;
/* u2_2068 Output nets */
wire t_6076,   t_6077,   t_6078;
/* u2_2069 Output nets */
wire t_6079,   t_6080,   t_6081;
/* u1_2070 Output nets */
wire t_6082,   t_6083;
/* u2_2071 Output nets */
wire t_6084,   t_6085,   t_6086;
/* u2_2072 Output nets */
wire t_6087,   t_6088,   t_6089;
/* u2_2073 Output nets */
wire t_6090,   t_6091,   t_6092;
/* u2_2074 Output nets */
wire t_6093,   t_6094,   t_6095;
/* u0_2075 Output nets */
wire t_6096,   t_6097;
/* u2_2076 Output nets */
wire t_6098,   t_6099,   t_6100;
/* u2_2077 Output nets */
wire t_6101,   t_6102,   t_6103;
/* u2_2078 Output nets */
wire t_6104,   t_6105,   t_6106;
/* u2_2079 Output nets */
wire t_6107,   t_6108,   t_6109;
/* u0_2080 Output nets */
wire t_6110,   t_6111;
/* u2_2081 Output nets */
wire t_6112,   t_6113,   t_6114;
/* u2_2082 Output nets */
wire t_6115,   t_6116,   t_6117;
/* u2_2083 Output nets */
wire t_6118,   t_6119,   t_6120;
/* u2_2084 Output nets */
wire t_6121,   t_6122,   t_6123;
/* u2_2085 Output nets */
wire t_6124,   t_6125,   t_6126;
/* u2_2086 Output nets */
wire t_6127,   t_6128,   t_6129;
/* u2_2087 Output nets */
wire t_6130,   t_6131,   t_6132;
/* u2_2088 Output nets */
wire t_6133,   t_6134,   t_6135;
/* u2_2089 Output nets */
wire t_6136,   t_6137,   t_6138;
/* u2_2090 Output nets */
wire t_6139,   t_6140,   t_6141;
/* u2_2091 Output nets */
wire t_6142,   t_6143,   t_6144;
/* u2_2092 Output nets */
wire t_6145,   t_6146,   t_6147;
/* u2_2093 Output nets */
wire t_6148,   t_6149,   t_6150;
/* u2_2094 Output nets */
wire t_6151,   t_6152,   t_6153;
/* u2_2095 Output nets */
wire t_6154,   t_6155,   t_6156;
/* u2_2096 Output nets */
wire t_6157,   t_6158,   t_6159;
/* u2_2097 Output nets */
wire t_6160,   t_6161,   t_6162;
/* u2_2098 Output nets */
wire t_6163,   t_6164,   t_6165;
/* u2_2099 Output nets */
wire t_6166,   t_6167,   t_6168;
/* u1_2100 Output nets */
wire t_6169,   t_6170;
/* u2_2101 Output nets */
wire t_6171,   t_6172,   t_6173;
/* u2_2102 Output nets */
wire t_6174,   t_6175,   t_6176;
/* u2_2103 Output nets */
wire t_6177,   t_6178,   t_6179;
/* u1_2104 Output nets */
wire t_6180,   t_6181;
/* u2_2105 Output nets */
wire t_6182,   t_6183,   t_6184;
/* u2_2106 Output nets */
wire t_6185,   t_6186,   t_6187;
/* u2_2107 Output nets */
wire t_6188,   t_6189,   t_6190;
/* u0_2108 Output nets */
wire t_6191,   t_6192;
/* u2_2109 Output nets */
wire t_6193,   t_6194,   t_6195;
/* u2_2110 Output nets */
wire t_6196,   t_6197,   t_6198;
/* u2_2111 Output nets */
wire t_6199,   t_6200,   t_6201;
/* u0_2112 Output nets */
wire t_6202,   t_6203;
/* u2_2113 Output nets */
wire t_6204,   t_6205,   t_6206;
/* u2_2114 Output nets */
wire t_6207,   t_6208,   t_6209;
/* u2_2115 Output nets */
wire t_6210,   t_6211,   t_6212;
/* u2_2116 Output nets */
wire t_6213,   t_6214,   t_6215;
/* u2_2117 Output nets */
wire t_6216,   t_6217,   t_6218;
/* u2_2118 Output nets */
wire t_6219,   t_6220,   t_6221;
/* u2_2119 Output nets */
wire t_6222,   t_6223,   t_6224;
/* u2_2120 Output nets */
wire t_6225,   t_6226,   t_6227;
/* u2_2121 Output nets */
wire t_6228,   t_6229,   t_6230;
/* u2_2122 Output nets */
wire t_6231,   t_6232,   t_6233;
/* u2_2123 Output nets */
wire t_6234,   t_6235,   t_6236;
/* u2_2124 Output nets */
wire t_6237,   t_6238,   t_6239;
/* u2_2125 Output nets */
wire t_6240,   t_6241,   t_6242;
/* u2_2126 Output nets */
wire t_6243,   t_6244,   t_6245;
/* u1_2127 Output nets */
wire t_6246,   t_6247;
/* u2_2128 Output nets */
wire t_6248,   t_6249,   t_6250;
/* u2_2129 Output nets */
wire t_6251,   t_6252,   t_6253;
/* u1_2130 Output nets */
wire t_6254,   t_6255;
/* u2_2131 Output nets */
wire t_6256,   t_6257,   t_6258;
/* u2_2132 Output nets */
wire t_6259,   t_6260,   t_6261;
/* u0_2133 Output nets */
wire t_6262,   t_6263;
/* u2_2134 Output nets */
wire t_6264,   t_6265,   t_6266;
/* u2_2135 Output nets */
wire t_6267,   t_6268,   t_6269;
/* u0_2136 Output nets */
wire t_6270,   t_6271;
/* u2_2137 Output nets */
wire t_6272,   t_6273,   t_6274;
/* u2_2138 Output nets */
wire t_6275,   t_6276,   t_6277;
/* u2_2139 Output nets */
wire t_6278,   t_6279,   t_6280;
/* u2_2140 Output nets */
wire t_6281,   t_6282,   t_6283;
/* u2_2141 Output nets */
wire t_6284,   t_6285,   t_6286;
/* u2_2142 Output nets */
wire t_6287,   t_6288,   t_6289;
/* u2_2143 Output nets */
wire t_6290,   t_6291,   t_6292;
/* u2_2144 Output nets */
wire t_6293,   t_6294,   t_6295;
/* u2_2145 Output nets */
wire t_6296,   t_6297,   t_6298;
/* u1_2146 Output nets */
wire t_6299,   t_6300;
/* u2_2147 Output nets */
wire t_6301,   t_6302,   t_6303;
/* u1_2148 Output nets */
wire t_6304,   t_6305;
/* u2_2149 Output nets */
wire t_6306,   t_6307,   t_6308;
/* u0_2150 Output nets */
wire t_6309,   t_6310;
/* u2_2151 Output nets */
wire t_6311,   t_6312,   t_6313;
/* u0_2152 Output nets */
wire t_6314,   t_6315;
/* u2_2153 Output nets */
wire t_6316,   t_6317,   t_6318;
/* u2_2154 Output nets */
wire t_6319,   t_6320,   t_6321;
/* u2_2155 Output nets */
wire t_6322,   t_6323,   t_6324;
/* u2_2156 Output nets */
wire t_6325,   t_6326,   t_6327;
/* u1_2157 Output nets */
wire t_6328,   t_6329;
/* u1_2158 Output nets */
wire t_6330,   t_6331;
/* u0_2159 Output nets */
wire t_6332,   t_6333;
/* u0_2160 Output nets */
wire t_6334;

/* compress stage 1 */
half_adder u0_1(.a(s_0_1), .b(s_0_0), .o(t_0), .cout(t_1));
compressor_3_2 u1_2(.a(s_2_2), .b(s_2_1), .cin(s_2_0), .o(t_2), .cout(t_3));
half_adder u0_3(.a(s_3_1), .b(s_3_0), .o(t_4), .cout(t_5));
compressor_3_2 u1_4(.a(s_4_2), .b(s_4_1), .cin(s_4_0), .o(t_6), .cout(t_7));
compressor_3_2 u1_5(.a(s_5_2), .b(s_5_1), .cin(s_5_0), .o(t_8), .cout(t_9));
compressor_4_2 u2_6(.a(s_6_4), .b(s_6_3), .c(s_6_2), .d(s_6_1), .cin(s_6_0), .o(t_10), .co(t_11), .cout(t_12));
compressor_4_2 u2_7(.a(s_7_3), .b(s_7_2), .c(s_7_1), .d(s_7_0), .cin(t_12), .o(t_13), .co(t_14), .cout(t_15));
compressor_4_2 u2_8(.a(s_8_3), .b(s_8_2), .c(s_8_1), .d(s_8_0), .cin(t_15), .o(t_16), .co(t_17), .cout(t_18));
half_adder u0_9(.a(s_8_5), .b(s_8_4), .o(t_19), .cout(t_20));
compressor_4_2 u2_10(.a(s_9_3), .b(s_9_2), .c(s_9_1), .d(s_9_0), .cin(t_18), .o(t_21), .co(t_22), .cout(t_23));
compressor_4_2 u2_11(.a(s_10_3), .b(s_10_2), .c(s_10_1), .d(s_10_0), .cin(t_23), .o(t_24), .co(t_25), .cout(t_26));
compressor_3_2 u1_12(.a(s_10_6), .b(s_10_5), .cin(s_10_4), .o(t_27), .cout(t_28));
compressor_4_2 u2_13(.a(s_11_3), .b(s_11_2), .c(s_11_1), .d(s_11_0), .cin(t_26), .o(t_29), .co(t_30), .cout(t_31));
half_adder u0_14(.a(s_11_5), .b(s_11_4), .o(t_32), .cout(t_33));
compressor_4_2 u2_15(.a(s_12_3), .b(s_12_2), .c(s_12_1), .d(s_12_0), .cin(t_31), .o(t_34), .co(t_35), .cout(t_36));
compressor_3_2 u1_16(.a(s_12_6), .b(s_12_5), .cin(s_12_4), .o(t_37), .cout(t_38));
compressor_4_2 u2_17(.a(s_13_3), .b(s_13_2), .c(s_13_1), .d(s_13_0), .cin(t_36), .o(t_39), .co(t_40), .cout(t_41));
compressor_3_2 u1_18(.a(s_13_6), .b(s_13_5), .cin(s_13_4), .o(t_42), .cout(t_43));
compressor_4_2 u2_19(.a(s_14_3), .b(s_14_2), .c(s_14_1), .d(s_14_0), .cin(t_41), .o(t_44), .co(t_45), .cout(t_46));
compressor_4_2 u2_20(.a(s_14_8), .b(s_14_7), .c(s_14_6), .d(s_14_5), .cin(s_14_4), .o(t_47), .co(t_48), .cout(t_49));
compressor_4_2 u2_21(.a(s_15_3), .b(s_15_2), .c(s_15_1), .d(s_15_0), .cin(t_46), .o(t_50), .co(t_51), .cout(t_52));
compressor_4_2 u2_22(.a(s_15_7), .b(s_15_6), .c(s_15_5), .d(s_15_4), .cin(t_49), .o(t_53), .co(t_54), .cout(t_55));
compressor_4_2 u2_23(.a(s_16_3), .b(s_16_2), .c(s_16_1), .d(s_16_0), .cin(t_52), .o(t_56), .co(t_57), .cout(t_58));
compressor_4_2 u2_24(.a(s_16_7), .b(s_16_6), .c(s_16_5), .d(s_16_4), .cin(t_55), .o(t_59), .co(t_60), .cout(t_61));
half_adder u0_25(.a(s_16_9), .b(s_16_8), .o(t_62), .cout(t_63));
compressor_4_2 u2_26(.a(s_17_3), .b(s_17_2), .c(s_17_1), .d(s_17_0), .cin(t_58), .o(t_64), .co(t_65), .cout(t_66));
compressor_4_2 u2_27(.a(s_17_7), .b(s_17_6), .c(s_17_5), .d(s_17_4), .cin(t_61), .o(t_67), .co(t_68), .cout(t_69));
compressor_4_2 u2_28(.a(s_18_3), .b(s_18_2), .c(s_18_1), .d(s_18_0), .cin(t_66), .o(t_70), .co(t_71), .cout(t_72));
compressor_4_2 u2_29(.a(s_18_7), .b(s_18_6), .c(s_18_5), .d(s_18_4), .cin(t_69), .o(t_73), .co(t_74), .cout(t_75));
compressor_3_2 u1_30(.a(s_18_10), .b(s_18_9), .cin(s_18_8), .o(t_76), .cout(t_77));
compressor_4_2 u2_31(.a(s_19_3), .b(s_19_2), .c(s_19_1), .d(s_19_0), .cin(t_72), .o(t_78), .co(t_79), .cout(t_80));
compressor_4_2 u2_32(.a(s_19_7), .b(s_19_6), .c(s_19_5), .d(s_19_4), .cin(t_75), .o(t_81), .co(t_82), .cout(t_83));
half_adder u0_33(.a(s_19_9), .b(s_19_8), .o(t_84), .cout(t_85));
compressor_4_2 u2_34(.a(s_20_3), .b(s_20_2), .c(s_20_1), .d(s_20_0), .cin(t_80), .o(t_86), .co(t_87), .cout(t_88));
compressor_4_2 u2_35(.a(s_20_7), .b(s_20_6), .c(s_20_5), .d(s_20_4), .cin(t_83), .o(t_89), .co(t_90), .cout(t_91));
compressor_3_2 u1_36(.a(s_20_10), .b(s_20_9), .cin(s_20_8), .o(t_92), .cout(t_93));
compressor_4_2 u2_37(.a(s_21_3), .b(s_21_2), .c(s_21_1), .d(s_21_0), .cin(t_88), .o(t_94), .co(t_95), .cout(t_96));
compressor_4_2 u2_38(.a(s_21_7), .b(s_21_6), .c(s_21_5), .d(s_21_4), .cin(t_91), .o(t_97), .co(t_98), .cout(t_99));
compressor_3_2 u1_39(.a(s_21_10), .b(s_21_9), .cin(s_21_8), .o(t_100), .cout(t_101));
compressor_4_2 u2_40(.a(s_22_3), .b(s_22_2), .c(s_22_1), .d(s_22_0), .cin(t_96), .o(t_102), .co(t_103), .cout(t_104));
compressor_4_2 u2_41(.a(s_22_7), .b(s_22_6), .c(s_22_5), .d(s_22_4), .cin(t_99), .o(t_105), .co(t_106), .cout(t_107));
compressor_4_2 u2_42(.a(s_22_12), .b(s_22_11), .c(s_22_10), .d(s_22_9), .cin(s_22_8), .o(t_108), .co(t_109), .cout(t_110));
compressor_4_2 u2_43(.a(s_23_3), .b(s_23_2), .c(s_23_1), .d(s_23_0), .cin(t_104), .o(t_111), .co(t_112), .cout(t_113));
compressor_4_2 u2_44(.a(s_23_7), .b(s_23_6), .c(s_23_5), .d(s_23_4), .cin(t_107), .o(t_114), .co(t_115), .cout(t_116));
compressor_4_2 u2_45(.a(s_23_11), .b(s_23_10), .c(s_23_9), .d(s_23_8), .cin(t_110), .o(t_117), .co(t_118), .cout(t_119));
compressor_4_2 u2_46(.a(s_24_3), .b(s_24_2), .c(s_24_1), .d(s_24_0), .cin(t_113), .o(t_120), .co(t_121), .cout(t_122));
compressor_4_2 u2_47(.a(s_24_7), .b(s_24_6), .c(s_24_5), .d(s_24_4), .cin(t_116), .o(t_123), .co(t_124), .cout(t_125));
compressor_4_2 u2_48(.a(s_24_11), .b(s_24_10), .c(s_24_9), .d(s_24_8), .cin(t_119), .o(t_126), .co(t_127), .cout(t_128));
half_adder u0_49(.a(s_24_13), .b(s_24_12), .o(t_129), .cout(t_130));
compressor_4_2 u2_50(.a(s_25_3), .b(s_25_2), .c(s_25_1), .d(s_25_0), .cin(t_122), .o(t_131), .co(t_132), .cout(t_133));
compressor_4_2 u2_51(.a(s_25_7), .b(s_25_6), .c(s_25_5), .d(s_25_4), .cin(t_125), .o(t_134), .co(t_135), .cout(t_136));
compressor_4_2 u2_52(.a(s_25_11), .b(s_25_10), .c(s_25_9), .d(s_25_8), .cin(t_128), .o(t_137), .co(t_138), .cout(t_139));
compressor_4_2 u2_53(.a(s_26_3), .b(s_26_2), .c(s_26_1), .d(s_26_0), .cin(t_133), .o(t_140), .co(t_141), .cout(t_142));
compressor_4_2 u2_54(.a(s_26_7), .b(s_26_6), .c(s_26_5), .d(s_26_4), .cin(t_136), .o(t_143), .co(t_144), .cout(t_145));
compressor_4_2 u2_55(.a(s_26_11), .b(s_26_10), .c(s_26_9), .d(s_26_8), .cin(t_139), .o(t_146), .co(t_147), .cout(t_148));
compressor_3_2 u1_56(.a(s_26_14), .b(s_26_13), .cin(s_26_12), .o(t_149), .cout(t_150));
compressor_4_2 u2_57(.a(s_27_3), .b(s_27_2), .c(s_27_1), .d(s_27_0), .cin(t_142), .o(t_151), .co(t_152), .cout(t_153));
compressor_4_2 u2_58(.a(s_27_7), .b(s_27_6), .c(s_27_5), .d(s_27_4), .cin(t_145), .o(t_154), .co(t_155), .cout(t_156));
compressor_4_2 u2_59(.a(s_27_11), .b(s_27_10), .c(s_27_9), .d(s_27_8), .cin(t_148), .o(t_157), .co(t_158), .cout(t_159));
half_adder u0_60(.a(s_27_13), .b(s_27_12), .o(t_160), .cout(t_161));
compressor_4_2 u2_61(.a(s_28_3), .b(s_28_2), .c(s_28_1), .d(s_28_0), .cin(t_153), .o(t_162), .co(t_163), .cout(t_164));
compressor_4_2 u2_62(.a(s_28_7), .b(s_28_6), .c(s_28_5), .d(s_28_4), .cin(t_156), .o(t_165), .co(t_166), .cout(t_167));
compressor_4_2 u2_63(.a(s_28_11), .b(s_28_10), .c(s_28_9), .d(s_28_8), .cin(t_159), .o(t_168), .co(t_169), .cout(t_170));
compressor_3_2 u1_64(.a(s_28_14), .b(s_28_13), .cin(s_28_12), .o(t_171), .cout(t_172));
compressor_4_2 u2_65(.a(s_29_3), .b(s_29_2), .c(s_29_1), .d(s_29_0), .cin(t_164), .o(t_173), .co(t_174), .cout(t_175));
compressor_4_2 u2_66(.a(s_29_7), .b(s_29_6), .c(s_29_5), .d(s_29_4), .cin(t_167), .o(t_176), .co(t_177), .cout(t_178));
compressor_4_2 u2_67(.a(s_29_11), .b(s_29_10), .c(s_29_9), .d(s_29_8), .cin(t_170), .o(t_179), .co(t_180), .cout(t_181));
compressor_3_2 u1_68(.a(s_29_14), .b(s_29_13), .cin(s_29_12), .o(t_182), .cout(t_183));
compressor_4_2 u2_69(.a(s_30_3), .b(s_30_2), .c(s_30_1), .d(s_30_0), .cin(t_175), .o(t_184), .co(t_185), .cout(t_186));
compressor_4_2 u2_70(.a(s_30_7), .b(s_30_6), .c(s_30_5), .d(s_30_4), .cin(t_178), .o(t_187), .co(t_188), .cout(t_189));
compressor_4_2 u2_71(.a(s_30_11), .b(s_30_10), .c(s_30_9), .d(s_30_8), .cin(t_181), .o(t_190), .co(t_191), .cout(t_192));
compressor_4_2 u2_72(.a(s_30_16), .b(s_30_15), .c(s_30_14), .d(s_30_13), .cin(s_30_12), .o(t_193), .co(t_194), .cout(t_195));
compressor_4_2 u2_73(.a(s_31_3), .b(s_31_2), .c(s_31_1), .d(s_31_0), .cin(t_186), .o(t_196), .co(t_197), .cout(t_198));
compressor_4_2 u2_74(.a(s_31_7), .b(s_31_6), .c(s_31_5), .d(s_31_4), .cin(t_189), .o(t_199), .co(t_200), .cout(t_201));
compressor_4_2 u2_75(.a(s_31_11), .b(s_31_10), .c(s_31_9), .d(s_31_8), .cin(t_192), .o(t_202), .co(t_203), .cout(t_204));
compressor_4_2 u2_76(.a(s_31_15), .b(s_31_14), .c(s_31_13), .d(s_31_12), .cin(t_195), .o(t_205), .co(t_206), .cout(t_207));
compressor_4_2 u2_77(.a(s_32_3), .b(s_32_2), .c(s_32_1), .d(s_32_0), .cin(t_198), .o(t_208), .co(t_209), .cout(t_210));
compressor_4_2 u2_78(.a(s_32_7), .b(s_32_6), .c(s_32_5), .d(s_32_4), .cin(t_201), .o(t_211), .co(t_212), .cout(t_213));
compressor_4_2 u2_79(.a(s_32_11), .b(s_32_10), .c(s_32_9), .d(s_32_8), .cin(t_204), .o(t_214), .co(t_215), .cout(t_216));
compressor_4_2 u2_80(.a(s_32_15), .b(s_32_14), .c(s_32_13), .d(s_32_12), .cin(t_207), .o(t_217), .co(t_218), .cout(t_219));
half_adder u0_81(.a(s_32_17), .b(s_32_16), .o(t_220), .cout(t_221));
compressor_4_2 u2_82(.a(s_33_3), .b(s_33_2), .c(s_33_1), .d(s_33_0), .cin(t_210), .o(t_222), .co(t_223), .cout(t_224));
compressor_4_2 u2_83(.a(s_33_7), .b(s_33_6), .c(s_33_5), .d(s_33_4), .cin(t_213), .o(t_225), .co(t_226), .cout(t_227));
compressor_4_2 u2_84(.a(s_33_11), .b(s_33_10), .c(s_33_9), .d(s_33_8), .cin(t_216), .o(t_228), .co(t_229), .cout(t_230));
compressor_4_2 u2_85(.a(s_33_15), .b(s_33_14), .c(s_33_13), .d(s_33_12), .cin(t_219), .o(t_231), .co(t_232), .cout(t_233));
compressor_4_2 u2_86(.a(s_34_3), .b(s_34_2), .c(s_34_1), .d(s_34_0), .cin(t_224), .o(t_234), .co(t_235), .cout(t_236));
compressor_4_2 u2_87(.a(s_34_7), .b(s_34_6), .c(s_34_5), .d(s_34_4), .cin(t_227), .o(t_237), .co(t_238), .cout(t_239));
compressor_4_2 u2_88(.a(s_34_11), .b(s_34_10), .c(s_34_9), .d(s_34_8), .cin(t_230), .o(t_240), .co(t_241), .cout(t_242));
compressor_4_2 u2_89(.a(s_34_15), .b(s_34_14), .c(s_34_13), .d(s_34_12), .cin(t_233), .o(t_243), .co(t_244), .cout(t_245));
compressor_3_2 u1_90(.a(s_34_18), .b(s_34_17), .cin(s_34_16), .o(t_246), .cout(t_247));
compressor_4_2 u2_91(.a(s_35_3), .b(s_35_2), .c(s_35_1), .d(s_35_0), .cin(t_236), .o(t_248), .co(t_249), .cout(t_250));
compressor_4_2 u2_92(.a(s_35_7), .b(s_35_6), .c(s_35_5), .d(s_35_4), .cin(t_239), .o(t_251), .co(t_252), .cout(t_253));
compressor_4_2 u2_93(.a(s_35_11), .b(s_35_10), .c(s_35_9), .d(s_35_8), .cin(t_242), .o(t_254), .co(t_255), .cout(t_256));
compressor_4_2 u2_94(.a(s_35_15), .b(s_35_14), .c(s_35_13), .d(s_35_12), .cin(t_245), .o(t_257), .co(t_258), .cout(t_259));
half_adder u0_95(.a(s_35_17), .b(s_35_16), .o(t_260), .cout(t_261));
compressor_4_2 u2_96(.a(s_36_3), .b(s_36_2), .c(s_36_1), .d(s_36_0), .cin(t_250), .o(t_262), .co(t_263), .cout(t_264));
compressor_4_2 u2_97(.a(s_36_7), .b(s_36_6), .c(s_36_5), .d(s_36_4), .cin(t_253), .o(t_265), .co(t_266), .cout(t_267));
compressor_4_2 u2_98(.a(s_36_11), .b(s_36_10), .c(s_36_9), .d(s_36_8), .cin(t_256), .o(t_268), .co(t_269), .cout(t_270));
compressor_4_2 u2_99(.a(s_36_15), .b(s_36_14), .c(s_36_13), .d(s_36_12), .cin(t_259), .o(t_271), .co(t_272), .cout(t_273));
compressor_3_2 u1_100(.a(s_36_18), .b(s_36_17), .cin(s_36_16), .o(t_274), .cout(t_275));
compressor_4_2 u2_101(.a(s_37_3), .b(s_37_2), .c(s_37_1), .d(s_37_0), .cin(t_264), .o(t_276), .co(t_277), .cout(t_278));
compressor_4_2 u2_102(.a(s_37_7), .b(s_37_6), .c(s_37_5), .d(s_37_4), .cin(t_267), .o(t_279), .co(t_280), .cout(t_281));
compressor_4_2 u2_103(.a(s_37_11), .b(s_37_10), .c(s_37_9), .d(s_37_8), .cin(t_270), .o(t_282), .co(t_283), .cout(t_284));
compressor_4_2 u2_104(.a(s_37_15), .b(s_37_14), .c(s_37_13), .d(s_37_12), .cin(t_273), .o(t_285), .co(t_286), .cout(t_287));
compressor_3_2 u1_105(.a(s_37_18), .b(s_37_17), .cin(s_37_16), .o(t_288), .cout(t_289));
compressor_4_2 u2_106(.a(s_38_3), .b(s_38_2), .c(s_38_1), .d(s_38_0), .cin(t_278), .o(t_290), .co(t_291), .cout(t_292));
compressor_4_2 u2_107(.a(s_38_7), .b(s_38_6), .c(s_38_5), .d(s_38_4), .cin(t_281), .o(t_293), .co(t_294), .cout(t_295));
compressor_4_2 u2_108(.a(s_38_11), .b(s_38_10), .c(s_38_9), .d(s_38_8), .cin(t_284), .o(t_296), .co(t_297), .cout(t_298));
compressor_4_2 u2_109(.a(s_38_15), .b(s_38_14), .c(s_38_13), .d(s_38_12), .cin(t_287), .o(t_299), .co(t_300), .cout(t_301));
compressor_4_2 u2_110(.a(s_38_20), .b(s_38_19), .c(s_38_18), .d(s_38_17), .cin(s_38_16), .o(t_302), .co(t_303), .cout(t_304));
compressor_4_2 u2_111(.a(s_39_3), .b(s_39_2), .c(s_39_1), .d(s_39_0), .cin(t_292), .o(t_305), .co(t_306), .cout(t_307));
compressor_4_2 u2_112(.a(s_39_7), .b(s_39_6), .c(s_39_5), .d(s_39_4), .cin(t_295), .o(t_308), .co(t_309), .cout(t_310));
compressor_4_2 u2_113(.a(s_39_11), .b(s_39_10), .c(s_39_9), .d(s_39_8), .cin(t_298), .o(t_311), .co(t_312), .cout(t_313));
compressor_4_2 u2_114(.a(s_39_15), .b(s_39_14), .c(s_39_13), .d(s_39_12), .cin(t_301), .o(t_314), .co(t_315), .cout(t_316));
compressor_4_2 u2_115(.a(s_39_19), .b(s_39_18), .c(s_39_17), .d(s_39_16), .cin(t_304), .o(t_317), .co(t_318), .cout(t_319));
compressor_4_2 u2_116(.a(s_40_3), .b(s_40_2), .c(s_40_1), .d(s_40_0), .cin(t_307), .o(t_320), .co(t_321), .cout(t_322));
compressor_4_2 u2_117(.a(s_40_7), .b(s_40_6), .c(s_40_5), .d(s_40_4), .cin(t_310), .o(t_323), .co(t_324), .cout(t_325));
compressor_4_2 u2_118(.a(s_40_11), .b(s_40_10), .c(s_40_9), .d(s_40_8), .cin(t_313), .o(t_326), .co(t_327), .cout(t_328));
compressor_4_2 u2_119(.a(s_40_15), .b(s_40_14), .c(s_40_13), .d(s_40_12), .cin(t_316), .o(t_329), .co(t_330), .cout(t_331));
compressor_4_2 u2_120(.a(s_40_19), .b(s_40_18), .c(s_40_17), .d(s_40_16), .cin(t_319), .o(t_332), .co(t_333), .cout(t_334));
half_adder u0_121(.a(s_40_21), .b(s_40_20), .o(t_335), .cout(t_336));
compressor_4_2 u2_122(.a(s_41_3), .b(s_41_2), .c(s_41_1), .d(s_41_0), .cin(t_322), .o(t_337), .co(t_338), .cout(t_339));
compressor_4_2 u2_123(.a(s_41_7), .b(s_41_6), .c(s_41_5), .d(s_41_4), .cin(t_325), .o(t_340), .co(t_341), .cout(t_342));
compressor_4_2 u2_124(.a(s_41_11), .b(s_41_10), .c(s_41_9), .d(s_41_8), .cin(t_328), .o(t_343), .co(t_344), .cout(t_345));
compressor_4_2 u2_125(.a(s_41_15), .b(s_41_14), .c(s_41_13), .d(s_41_12), .cin(t_331), .o(t_346), .co(t_347), .cout(t_348));
compressor_4_2 u2_126(.a(s_41_19), .b(s_41_18), .c(s_41_17), .d(s_41_16), .cin(t_334), .o(t_349), .co(t_350), .cout(t_351));
compressor_4_2 u2_127(.a(s_42_3), .b(s_42_2), .c(s_42_1), .d(s_42_0), .cin(t_339), .o(t_352), .co(t_353), .cout(t_354));
compressor_4_2 u2_128(.a(s_42_7), .b(s_42_6), .c(s_42_5), .d(s_42_4), .cin(t_342), .o(t_355), .co(t_356), .cout(t_357));
compressor_4_2 u2_129(.a(s_42_11), .b(s_42_10), .c(s_42_9), .d(s_42_8), .cin(t_345), .o(t_358), .co(t_359), .cout(t_360));
compressor_4_2 u2_130(.a(s_42_15), .b(s_42_14), .c(s_42_13), .d(s_42_12), .cin(t_348), .o(t_361), .co(t_362), .cout(t_363));
compressor_4_2 u2_131(.a(s_42_19), .b(s_42_18), .c(s_42_17), .d(s_42_16), .cin(t_351), .o(t_364), .co(t_365), .cout(t_366));
compressor_3_2 u1_132(.a(s_42_22), .b(s_42_21), .cin(s_42_20), .o(t_367), .cout(t_368));
compressor_4_2 u2_133(.a(s_43_3), .b(s_43_2), .c(s_43_1), .d(s_43_0), .cin(t_354), .o(t_369), .co(t_370), .cout(t_371));
compressor_4_2 u2_134(.a(s_43_7), .b(s_43_6), .c(s_43_5), .d(s_43_4), .cin(t_357), .o(t_372), .co(t_373), .cout(t_374));
compressor_4_2 u2_135(.a(s_43_11), .b(s_43_10), .c(s_43_9), .d(s_43_8), .cin(t_360), .o(t_375), .co(t_376), .cout(t_377));
compressor_4_2 u2_136(.a(s_43_15), .b(s_43_14), .c(s_43_13), .d(s_43_12), .cin(t_363), .o(t_378), .co(t_379), .cout(t_380));
compressor_4_2 u2_137(.a(s_43_19), .b(s_43_18), .c(s_43_17), .d(s_43_16), .cin(t_366), .o(t_381), .co(t_382), .cout(t_383));
half_adder u0_138(.a(s_43_21), .b(s_43_20), .o(t_384), .cout(t_385));
compressor_4_2 u2_139(.a(s_44_3), .b(s_44_2), .c(s_44_1), .d(s_44_0), .cin(t_371), .o(t_386), .co(t_387), .cout(t_388));
compressor_4_2 u2_140(.a(s_44_7), .b(s_44_6), .c(s_44_5), .d(s_44_4), .cin(t_374), .o(t_389), .co(t_390), .cout(t_391));
compressor_4_2 u2_141(.a(s_44_11), .b(s_44_10), .c(s_44_9), .d(s_44_8), .cin(t_377), .o(t_392), .co(t_393), .cout(t_394));
compressor_4_2 u2_142(.a(s_44_15), .b(s_44_14), .c(s_44_13), .d(s_44_12), .cin(t_380), .o(t_395), .co(t_396), .cout(t_397));
compressor_4_2 u2_143(.a(s_44_19), .b(s_44_18), .c(s_44_17), .d(s_44_16), .cin(t_383), .o(t_398), .co(t_399), .cout(t_400));
compressor_3_2 u1_144(.a(s_44_22), .b(s_44_21), .cin(s_44_20), .o(t_401), .cout(t_402));
compressor_4_2 u2_145(.a(s_45_3), .b(s_45_2), .c(s_45_1), .d(s_45_0), .cin(t_388), .o(t_403), .co(t_404), .cout(t_405));
compressor_4_2 u2_146(.a(s_45_7), .b(s_45_6), .c(s_45_5), .d(s_45_4), .cin(t_391), .o(t_406), .co(t_407), .cout(t_408));
compressor_4_2 u2_147(.a(s_45_11), .b(s_45_10), .c(s_45_9), .d(s_45_8), .cin(t_394), .o(t_409), .co(t_410), .cout(t_411));
compressor_4_2 u2_148(.a(s_45_15), .b(s_45_14), .c(s_45_13), .d(s_45_12), .cin(t_397), .o(t_412), .co(t_413), .cout(t_414));
compressor_4_2 u2_149(.a(s_45_19), .b(s_45_18), .c(s_45_17), .d(s_45_16), .cin(t_400), .o(t_415), .co(t_416), .cout(t_417));
compressor_3_2 u1_150(.a(s_45_22), .b(s_45_21), .cin(s_45_20), .o(t_418), .cout(t_419));
compressor_4_2 u2_151(.a(s_46_3), .b(s_46_2), .c(s_46_1), .d(s_46_0), .cin(t_405), .o(t_420), .co(t_421), .cout(t_422));
compressor_4_2 u2_152(.a(s_46_7), .b(s_46_6), .c(s_46_5), .d(s_46_4), .cin(t_408), .o(t_423), .co(t_424), .cout(t_425));
compressor_4_2 u2_153(.a(s_46_11), .b(s_46_10), .c(s_46_9), .d(s_46_8), .cin(t_411), .o(t_426), .co(t_427), .cout(t_428));
compressor_4_2 u2_154(.a(s_46_15), .b(s_46_14), .c(s_46_13), .d(s_46_12), .cin(t_414), .o(t_429), .co(t_430), .cout(t_431));
compressor_4_2 u2_155(.a(s_46_19), .b(s_46_18), .c(s_46_17), .d(s_46_16), .cin(t_417), .o(t_432), .co(t_433), .cout(t_434));
compressor_4_2 u2_156(.a(s_46_24), .b(s_46_23), .c(s_46_22), .d(s_46_21), .cin(s_46_20), .o(t_435), .co(t_436), .cout(t_437));
compressor_4_2 u2_157(.a(s_47_3), .b(s_47_2), .c(s_47_1), .d(s_47_0), .cin(t_422), .o(t_438), .co(t_439), .cout(t_440));
compressor_4_2 u2_158(.a(s_47_7), .b(s_47_6), .c(s_47_5), .d(s_47_4), .cin(t_425), .o(t_441), .co(t_442), .cout(t_443));
compressor_4_2 u2_159(.a(s_47_11), .b(s_47_10), .c(s_47_9), .d(s_47_8), .cin(t_428), .o(t_444), .co(t_445), .cout(t_446));
compressor_4_2 u2_160(.a(s_47_15), .b(s_47_14), .c(s_47_13), .d(s_47_12), .cin(t_431), .o(t_447), .co(t_448), .cout(t_449));
compressor_4_2 u2_161(.a(s_47_19), .b(s_47_18), .c(s_47_17), .d(s_47_16), .cin(t_434), .o(t_450), .co(t_451), .cout(t_452));
compressor_4_2 u2_162(.a(s_47_23), .b(s_47_22), .c(s_47_21), .d(s_47_20), .cin(t_437), .o(t_453), .co(t_454), .cout(t_455));
compressor_4_2 u2_163(.a(s_48_3), .b(s_48_2), .c(s_48_1), .d(s_48_0), .cin(t_440), .o(t_456), .co(t_457), .cout(t_458));
compressor_4_2 u2_164(.a(s_48_7), .b(s_48_6), .c(s_48_5), .d(s_48_4), .cin(t_443), .o(t_459), .co(t_460), .cout(t_461));
compressor_4_2 u2_165(.a(s_48_11), .b(s_48_10), .c(s_48_9), .d(s_48_8), .cin(t_446), .o(t_462), .co(t_463), .cout(t_464));
compressor_4_2 u2_166(.a(s_48_15), .b(s_48_14), .c(s_48_13), .d(s_48_12), .cin(t_449), .o(t_465), .co(t_466), .cout(t_467));
compressor_4_2 u2_167(.a(s_48_19), .b(s_48_18), .c(s_48_17), .d(s_48_16), .cin(t_452), .o(t_468), .co(t_469), .cout(t_470));
compressor_4_2 u2_168(.a(s_48_23), .b(s_48_22), .c(s_48_21), .d(s_48_20), .cin(t_455), .o(t_471), .co(t_472), .cout(t_473));
half_adder u0_169(.a(s_48_25), .b(s_48_24), .o(t_474), .cout(t_475));
compressor_4_2 u2_170(.a(s_49_3), .b(s_49_2), .c(s_49_1), .d(s_49_0), .cin(t_458), .o(t_476), .co(t_477), .cout(t_478));
compressor_4_2 u2_171(.a(s_49_7), .b(s_49_6), .c(s_49_5), .d(s_49_4), .cin(t_461), .o(t_479), .co(t_480), .cout(t_481));
compressor_4_2 u2_172(.a(s_49_11), .b(s_49_10), .c(s_49_9), .d(s_49_8), .cin(t_464), .o(t_482), .co(t_483), .cout(t_484));
compressor_4_2 u2_173(.a(s_49_15), .b(s_49_14), .c(s_49_13), .d(s_49_12), .cin(t_467), .o(t_485), .co(t_486), .cout(t_487));
compressor_4_2 u2_174(.a(s_49_19), .b(s_49_18), .c(s_49_17), .d(s_49_16), .cin(t_470), .o(t_488), .co(t_489), .cout(t_490));
compressor_4_2 u2_175(.a(s_49_23), .b(s_49_22), .c(s_49_21), .d(s_49_20), .cin(t_473), .o(t_491), .co(t_492), .cout(t_493));
compressor_4_2 u2_176(.a(s_50_3), .b(s_50_2), .c(s_50_1), .d(s_50_0), .cin(t_478), .o(t_494), .co(t_495), .cout(t_496));
compressor_4_2 u2_177(.a(s_50_7), .b(s_50_6), .c(s_50_5), .d(s_50_4), .cin(t_481), .o(t_497), .co(t_498), .cout(t_499));
compressor_4_2 u2_178(.a(s_50_11), .b(s_50_10), .c(s_50_9), .d(s_50_8), .cin(t_484), .o(t_500), .co(t_501), .cout(t_502));
compressor_4_2 u2_179(.a(s_50_15), .b(s_50_14), .c(s_50_13), .d(s_50_12), .cin(t_487), .o(t_503), .co(t_504), .cout(t_505));
compressor_4_2 u2_180(.a(s_50_19), .b(s_50_18), .c(s_50_17), .d(s_50_16), .cin(t_490), .o(t_506), .co(t_507), .cout(t_508));
compressor_4_2 u2_181(.a(s_50_23), .b(s_50_22), .c(s_50_21), .d(s_50_20), .cin(t_493), .o(t_509), .co(t_510), .cout(t_511));
compressor_3_2 u1_182(.a(s_50_26), .b(s_50_25), .cin(s_50_24), .o(t_512), .cout(t_513));
compressor_4_2 u2_183(.a(s_51_3), .b(s_51_2), .c(s_51_1), .d(s_51_0), .cin(t_496), .o(t_514), .co(t_515), .cout(t_516));
compressor_4_2 u2_184(.a(s_51_7), .b(s_51_6), .c(s_51_5), .d(s_51_4), .cin(t_499), .o(t_517), .co(t_518), .cout(t_519));
compressor_4_2 u2_185(.a(s_51_11), .b(s_51_10), .c(s_51_9), .d(s_51_8), .cin(t_502), .o(t_520), .co(t_521), .cout(t_522));
compressor_4_2 u2_186(.a(s_51_15), .b(s_51_14), .c(s_51_13), .d(s_51_12), .cin(t_505), .o(t_523), .co(t_524), .cout(t_525));
compressor_4_2 u2_187(.a(s_51_19), .b(s_51_18), .c(s_51_17), .d(s_51_16), .cin(t_508), .o(t_526), .co(t_527), .cout(t_528));
compressor_4_2 u2_188(.a(s_51_23), .b(s_51_22), .c(s_51_21), .d(s_51_20), .cin(t_511), .o(t_529), .co(t_530), .cout(t_531));
half_adder u0_189(.a(s_51_25), .b(s_51_24), .o(t_532), .cout(t_533));
compressor_4_2 u2_190(.a(s_52_3), .b(s_52_2), .c(s_52_1), .d(s_52_0), .cin(t_516), .o(t_534), .co(t_535), .cout(t_536));
compressor_4_2 u2_191(.a(s_52_7), .b(s_52_6), .c(s_52_5), .d(s_52_4), .cin(t_519), .o(t_537), .co(t_538), .cout(t_539));
compressor_4_2 u2_192(.a(s_52_11), .b(s_52_10), .c(s_52_9), .d(s_52_8), .cin(t_522), .o(t_540), .co(t_541), .cout(t_542));
compressor_4_2 u2_193(.a(s_52_15), .b(s_52_14), .c(s_52_13), .d(s_52_12), .cin(t_525), .o(t_543), .co(t_544), .cout(t_545));
compressor_4_2 u2_194(.a(s_52_19), .b(s_52_18), .c(s_52_17), .d(s_52_16), .cin(t_528), .o(t_546), .co(t_547), .cout(t_548));
compressor_4_2 u2_195(.a(s_52_23), .b(s_52_22), .c(s_52_21), .d(s_52_20), .cin(t_531), .o(t_549), .co(t_550), .cout(t_551));
compressor_3_2 u1_196(.a(s_52_26), .b(s_52_25), .cin(s_52_24), .o(t_552), .cout(t_553));
compressor_4_2 u2_197(.a(s_53_3), .b(s_53_2), .c(s_53_1), .d(s_53_0), .cin(t_536), .o(t_554), .co(t_555), .cout(t_556));
compressor_4_2 u2_198(.a(s_53_7), .b(s_53_6), .c(s_53_5), .d(s_53_4), .cin(t_539), .o(t_557), .co(t_558), .cout(t_559));
compressor_4_2 u2_199(.a(s_53_11), .b(s_53_10), .c(s_53_9), .d(s_53_8), .cin(t_542), .o(t_560), .co(t_561), .cout(t_562));
compressor_4_2 u2_200(.a(s_53_15), .b(s_53_14), .c(s_53_13), .d(s_53_12), .cin(t_545), .o(t_563), .co(t_564), .cout(t_565));
compressor_4_2 u2_201(.a(s_53_19), .b(s_53_18), .c(s_53_17), .d(s_53_16), .cin(t_548), .o(t_566), .co(t_567), .cout(t_568));
compressor_4_2 u2_202(.a(s_53_23), .b(s_53_22), .c(s_53_21), .d(s_53_20), .cin(t_551), .o(t_569), .co(t_570), .cout(t_571));
compressor_3_2 u1_203(.a(s_53_26), .b(s_53_25), .cin(s_53_24), .o(t_572), .cout(t_573));
compressor_4_2 u2_204(.a(s_54_3), .b(s_54_2), .c(s_54_1), .d(s_54_0), .cin(t_556), .o(t_574), .co(t_575), .cout(t_576));
compressor_4_2 u2_205(.a(s_54_7), .b(s_54_6), .c(s_54_5), .d(s_54_4), .cin(t_559), .o(t_577), .co(t_578), .cout(t_579));
compressor_4_2 u2_206(.a(s_54_11), .b(s_54_10), .c(s_54_9), .d(s_54_8), .cin(t_562), .o(t_580), .co(t_581), .cout(t_582));
compressor_4_2 u2_207(.a(s_54_15), .b(s_54_14), .c(s_54_13), .d(s_54_12), .cin(t_565), .o(t_583), .co(t_584), .cout(t_585));
compressor_4_2 u2_208(.a(s_54_19), .b(s_54_18), .c(s_54_17), .d(s_54_16), .cin(t_568), .o(t_586), .co(t_587), .cout(t_588));
compressor_4_2 u2_209(.a(s_54_23), .b(s_54_22), .c(s_54_21), .d(s_54_20), .cin(t_571), .o(t_589), .co(t_590), .cout(t_591));
compressor_4_2 u2_210(.a(s_54_28), .b(s_54_27), .c(s_54_26), .d(s_54_25), .cin(s_54_24), .o(t_592), .co(t_593), .cout(t_594));
compressor_4_2 u2_211(.a(s_55_3), .b(s_55_2), .c(s_55_1), .d(s_55_0), .cin(t_576), .o(t_595), .co(t_596), .cout(t_597));
compressor_4_2 u2_212(.a(s_55_7), .b(s_55_6), .c(s_55_5), .d(s_55_4), .cin(t_579), .o(t_598), .co(t_599), .cout(t_600));
compressor_4_2 u2_213(.a(s_55_11), .b(s_55_10), .c(s_55_9), .d(s_55_8), .cin(t_582), .o(t_601), .co(t_602), .cout(t_603));
compressor_4_2 u2_214(.a(s_55_15), .b(s_55_14), .c(s_55_13), .d(s_55_12), .cin(t_585), .o(t_604), .co(t_605), .cout(t_606));
compressor_4_2 u2_215(.a(s_55_19), .b(s_55_18), .c(s_55_17), .d(s_55_16), .cin(t_588), .o(t_607), .co(t_608), .cout(t_609));
compressor_4_2 u2_216(.a(s_55_23), .b(s_55_22), .c(s_55_21), .d(s_55_20), .cin(t_591), .o(t_610), .co(t_611), .cout(t_612));
compressor_4_2 u2_217(.a(s_55_27), .b(s_55_26), .c(s_55_25), .d(s_55_24), .cin(t_594), .o(t_613), .co(t_614), .cout(t_615));
compressor_4_2 u2_218(.a(s_56_3), .b(s_56_2), .c(s_56_1), .d(s_56_0), .cin(t_597), .o(t_616), .co(t_617), .cout(t_618));
compressor_4_2 u2_219(.a(s_56_7), .b(s_56_6), .c(s_56_5), .d(s_56_4), .cin(t_600), .o(t_619), .co(t_620), .cout(t_621));
compressor_4_2 u2_220(.a(s_56_11), .b(s_56_10), .c(s_56_9), .d(s_56_8), .cin(t_603), .o(t_622), .co(t_623), .cout(t_624));
compressor_4_2 u2_221(.a(s_56_15), .b(s_56_14), .c(s_56_13), .d(s_56_12), .cin(t_606), .o(t_625), .co(t_626), .cout(t_627));
compressor_4_2 u2_222(.a(s_56_19), .b(s_56_18), .c(s_56_17), .d(s_56_16), .cin(t_609), .o(t_628), .co(t_629), .cout(t_630));
compressor_4_2 u2_223(.a(s_56_23), .b(s_56_22), .c(s_56_21), .d(s_56_20), .cin(t_612), .o(t_631), .co(t_632), .cout(t_633));
compressor_4_2 u2_224(.a(s_56_27), .b(s_56_26), .c(s_56_25), .d(s_56_24), .cin(t_615), .o(t_634), .co(t_635), .cout(t_636));
half_adder u0_225(.a(s_56_29), .b(s_56_28), .o(t_637), .cout(t_638));
compressor_4_2 u2_226(.a(s_57_3), .b(s_57_2), .c(s_57_1), .d(s_57_0), .cin(t_618), .o(t_639), .co(t_640), .cout(t_641));
compressor_4_2 u2_227(.a(s_57_7), .b(s_57_6), .c(s_57_5), .d(s_57_4), .cin(t_621), .o(t_642), .co(t_643), .cout(t_644));
compressor_4_2 u2_228(.a(s_57_11), .b(s_57_10), .c(s_57_9), .d(s_57_8), .cin(t_624), .o(t_645), .co(t_646), .cout(t_647));
compressor_4_2 u2_229(.a(s_57_15), .b(s_57_14), .c(s_57_13), .d(s_57_12), .cin(t_627), .o(t_648), .co(t_649), .cout(t_650));
compressor_4_2 u2_230(.a(s_57_19), .b(s_57_18), .c(s_57_17), .d(s_57_16), .cin(t_630), .o(t_651), .co(t_652), .cout(t_653));
compressor_4_2 u2_231(.a(s_57_23), .b(s_57_22), .c(s_57_21), .d(s_57_20), .cin(t_633), .o(t_654), .co(t_655), .cout(t_656));
compressor_4_2 u2_232(.a(s_57_27), .b(s_57_26), .c(s_57_25), .d(s_57_24), .cin(t_636), .o(t_657), .co(t_658), .cout(t_659));
compressor_4_2 u2_233(.a(s_58_3), .b(s_58_2), .c(s_58_1), .d(s_58_0), .cin(t_641), .o(t_660), .co(t_661), .cout(t_662));
compressor_4_2 u2_234(.a(s_58_7), .b(s_58_6), .c(s_58_5), .d(s_58_4), .cin(t_644), .o(t_663), .co(t_664), .cout(t_665));
compressor_4_2 u2_235(.a(s_58_11), .b(s_58_10), .c(s_58_9), .d(s_58_8), .cin(t_647), .o(t_666), .co(t_667), .cout(t_668));
compressor_4_2 u2_236(.a(s_58_15), .b(s_58_14), .c(s_58_13), .d(s_58_12), .cin(t_650), .o(t_669), .co(t_670), .cout(t_671));
compressor_4_2 u2_237(.a(s_58_19), .b(s_58_18), .c(s_58_17), .d(s_58_16), .cin(t_653), .o(t_672), .co(t_673), .cout(t_674));
compressor_4_2 u2_238(.a(s_58_23), .b(s_58_22), .c(s_58_21), .d(s_58_20), .cin(t_656), .o(t_675), .co(t_676), .cout(t_677));
compressor_4_2 u2_239(.a(s_58_27), .b(s_58_26), .c(s_58_25), .d(s_58_24), .cin(t_659), .o(t_678), .co(t_679), .cout(t_680));
compressor_3_2 u1_240(.a(s_58_30), .b(s_58_29), .cin(s_58_28), .o(t_681), .cout(t_682));
compressor_4_2 u2_241(.a(s_59_3), .b(s_59_2), .c(s_59_1), .d(s_59_0), .cin(t_662), .o(t_683), .co(t_684), .cout(t_685));
compressor_4_2 u2_242(.a(s_59_7), .b(s_59_6), .c(s_59_5), .d(s_59_4), .cin(t_665), .o(t_686), .co(t_687), .cout(t_688));
compressor_4_2 u2_243(.a(s_59_11), .b(s_59_10), .c(s_59_9), .d(s_59_8), .cin(t_668), .o(t_689), .co(t_690), .cout(t_691));
compressor_4_2 u2_244(.a(s_59_15), .b(s_59_14), .c(s_59_13), .d(s_59_12), .cin(t_671), .o(t_692), .co(t_693), .cout(t_694));
compressor_4_2 u2_245(.a(s_59_19), .b(s_59_18), .c(s_59_17), .d(s_59_16), .cin(t_674), .o(t_695), .co(t_696), .cout(t_697));
compressor_4_2 u2_246(.a(s_59_23), .b(s_59_22), .c(s_59_21), .d(s_59_20), .cin(t_677), .o(t_698), .co(t_699), .cout(t_700));
compressor_4_2 u2_247(.a(s_59_27), .b(s_59_26), .c(s_59_25), .d(s_59_24), .cin(t_680), .o(t_701), .co(t_702), .cout(t_703));
half_adder u0_248(.a(s_59_29), .b(s_59_28), .o(t_704), .cout(t_705));
compressor_4_2 u2_249(.a(s_60_3), .b(s_60_2), .c(s_60_1), .d(s_60_0), .cin(t_685), .o(t_706), .co(t_707), .cout(t_708));
compressor_4_2 u2_250(.a(s_60_7), .b(s_60_6), .c(s_60_5), .d(s_60_4), .cin(t_688), .o(t_709), .co(t_710), .cout(t_711));
compressor_4_2 u2_251(.a(s_60_11), .b(s_60_10), .c(s_60_9), .d(s_60_8), .cin(t_691), .o(t_712), .co(t_713), .cout(t_714));
compressor_4_2 u2_252(.a(s_60_15), .b(s_60_14), .c(s_60_13), .d(s_60_12), .cin(t_694), .o(t_715), .co(t_716), .cout(t_717));
compressor_4_2 u2_253(.a(s_60_19), .b(s_60_18), .c(s_60_17), .d(s_60_16), .cin(t_697), .o(t_718), .co(t_719), .cout(t_720));
compressor_4_2 u2_254(.a(s_60_23), .b(s_60_22), .c(s_60_21), .d(s_60_20), .cin(t_700), .o(t_721), .co(t_722), .cout(t_723));
compressor_4_2 u2_255(.a(s_60_27), .b(s_60_26), .c(s_60_25), .d(s_60_24), .cin(t_703), .o(t_724), .co(t_725), .cout(t_726));
compressor_3_2 u1_256(.a(s_60_30), .b(s_60_29), .cin(s_60_28), .o(t_727), .cout(t_728));
compressor_4_2 u2_257(.a(s_61_3), .b(s_61_2), .c(s_61_1), .d(s_61_0), .cin(t_708), .o(t_729), .co(t_730), .cout(t_731));
compressor_4_2 u2_258(.a(s_61_7), .b(s_61_6), .c(s_61_5), .d(s_61_4), .cin(t_711), .o(t_732), .co(t_733), .cout(t_734));
compressor_4_2 u2_259(.a(s_61_11), .b(s_61_10), .c(s_61_9), .d(s_61_8), .cin(t_714), .o(t_735), .co(t_736), .cout(t_737));
compressor_4_2 u2_260(.a(s_61_15), .b(s_61_14), .c(s_61_13), .d(s_61_12), .cin(t_717), .o(t_738), .co(t_739), .cout(t_740));
compressor_4_2 u2_261(.a(s_61_19), .b(s_61_18), .c(s_61_17), .d(s_61_16), .cin(t_720), .o(t_741), .co(t_742), .cout(t_743));
compressor_4_2 u2_262(.a(s_61_23), .b(s_61_22), .c(s_61_21), .d(s_61_20), .cin(t_723), .o(t_744), .co(t_745), .cout(t_746));
compressor_4_2 u2_263(.a(s_61_27), .b(s_61_26), .c(s_61_25), .d(s_61_24), .cin(t_726), .o(t_747), .co(t_748), .cout(t_749));
compressor_3_2 u1_264(.a(s_61_30), .b(s_61_29), .cin(s_61_28), .o(t_750), .cout(t_751));
compressor_4_2 u2_265(.a(s_62_3), .b(s_62_2), .c(s_62_1), .d(s_62_0), .cin(t_731), .o(t_752), .co(t_753), .cout(t_754));
compressor_4_2 u2_266(.a(s_62_7), .b(s_62_6), .c(s_62_5), .d(s_62_4), .cin(t_734), .o(t_755), .co(t_756), .cout(t_757));
compressor_4_2 u2_267(.a(s_62_11), .b(s_62_10), .c(s_62_9), .d(s_62_8), .cin(t_737), .o(t_758), .co(t_759), .cout(t_760));
compressor_4_2 u2_268(.a(s_62_15), .b(s_62_14), .c(s_62_13), .d(s_62_12), .cin(t_740), .o(t_761), .co(t_762), .cout(t_763));
compressor_4_2 u2_269(.a(s_62_19), .b(s_62_18), .c(s_62_17), .d(s_62_16), .cin(t_743), .o(t_764), .co(t_765), .cout(t_766));
compressor_4_2 u2_270(.a(s_62_23), .b(s_62_22), .c(s_62_21), .d(s_62_20), .cin(t_746), .o(t_767), .co(t_768), .cout(t_769));
compressor_4_2 u2_271(.a(s_62_27), .b(s_62_26), .c(s_62_25), .d(s_62_24), .cin(t_749), .o(t_770), .co(t_771), .cout(t_772));
compressor_4_2 u2_272(.a(s_62_32), .b(s_62_31), .c(s_62_30), .d(s_62_29), .cin(s_62_28), .o(t_773), .co(t_774), .cout(t_775));
compressor_4_2 u2_273(.a(s_63_3), .b(s_63_2), .c(s_63_1), .d(s_63_0), .cin(t_754), .o(t_776), .co(t_777), .cout(t_778));
compressor_4_2 u2_274(.a(s_63_7), .b(s_63_6), .c(s_63_5), .d(s_63_4), .cin(t_757), .o(t_779), .co(t_780), .cout(t_781));
compressor_4_2 u2_275(.a(s_63_11), .b(s_63_10), .c(s_63_9), .d(s_63_8), .cin(t_760), .o(t_782), .co(t_783), .cout(t_784));
compressor_4_2 u2_276(.a(s_63_15), .b(s_63_14), .c(s_63_13), .d(s_63_12), .cin(t_763), .o(t_785), .co(t_786), .cout(t_787));
compressor_4_2 u2_277(.a(s_63_19), .b(s_63_18), .c(s_63_17), .d(s_63_16), .cin(t_766), .o(t_788), .co(t_789), .cout(t_790));
compressor_4_2 u2_278(.a(s_63_23), .b(s_63_22), .c(s_63_21), .d(s_63_20), .cin(t_769), .o(t_791), .co(t_792), .cout(t_793));
compressor_4_2 u2_279(.a(s_63_27), .b(s_63_26), .c(s_63_25), .d(s_63_24), .cin(t_772), .o(t_794), .co(t_795), .cout(t_796));
compressor_4_2 u2_280(.a(s_63_31), .b(s_63_30), .c(s_63_29), .d(s_63_28), .cin(t_775), .o(t_797), .co(t_798), .cout(t_799));
compressor_4_2 u2_281(.a(s_64_3), .b(s_64_2), .c(s_64_1), .d(s_64_0), .cin(t_778), .o(t_800), .co(t_801), .cout(t_802));
compressor_4_2 u2_282(.a(s_64_7), .b(s_64_6), .c(s_64_5), .d(s_64_4), .cin(t_781), .o(t_803), .co(t_804), .cout(t_805));
compressor_4_2 u2_283(.a(s_64_11), .b(s_64_10), .c(s_64_9), .d(s_64_8), .cin(t_784), .o(t_806), .co(t_807), .cout(t_808));
compressor_4_2 u2_284(.a(s_64_15), .b(s_64_14), .c(s_64_13), .d(s_64_12), .cin(t_787), .o(t_809), .co(t_810), .cout(t_811));
compressor_4_2 u2_285(.a(s_64_19), .b(s_64_18), .c(s_64_17), .d(s_64_16), .cin(t_790), .o(t_812), .co(t_813), .cout(t_814));
compressor_4_2 u2_286(.a(s_64_23), .b(s_64_22), .c(s_64_21), .d(s_64_20), .cin(t_793), .o(t_815), .co(t_816), .cout(t_817));
compressor_4_2 u2_287(.a(s_64_27), .b(s_64_26), .c(s_64_25), .d(s_64_24), .cin(t_796), .o(t_818), .co(t_819), .cout(t_820));
compressor_4_2 u2_288(.a(s_64_31), .b(s_64_30), .c(s_64_29), .d(s_64_28), .cin(t_799), .o(t_821), .co(t_822), .cout(t_823));
half_adder u0_289(.a(s_64_33), .b(s_64_32), .o(t_824), .cout(t_825));
compressor_4_2 u2_290(.a(s_65_3), .b(s_65_2), .c(s_65_1), .d(s_65_0), .cin(t_802), .o(t_826), .co(t_827), .cout(t_828));
compressor_4_2 u2_291(.a(s_65_7), .b(s_65_6), .c(s_65_5), .d(s_65_4), .cin(t_805), .o(t_829), .co(t_830), .cout(t_831));
compressor_4_2 u2_292(.a(s_65_11), .b(s_65_10), .c(s_65_9), .d(s_65_8), .cin(t_808), .o(t_832), .co(t_833), .cout(t_834));
compressor_4_2 u2_293(.a(s_65_15), .b(s_65_14), .c(s_65_13), .d(s_65_12), .cin(t_811), .o(t_835), .co(t_836), .cout(t_837));
compressor_4_2 u2_294(.a(s_65_19), .b(s_65_18), .c(s_65_17), .d(s_65_16), .cin(t_814), .o(t_838), .co(t_839), .cout(t_840));
compressor_4_2 u2_295(.a(s_65_23), .b(s_65_22), .c(s_65_21), .d(s_65_20), .cin(t_817), .o(t_841), .co(t_842), .cout(t_843));
compressor_4_2 u2_296(.a(s_65_27), .b(s_65_26), .c(s_65_25), .d(s_65_24), .cin(t_820), .o(t_844), .co(t_845), .cout(t_846));
compressor_4_2 u2_297(.a(s_65_31), .b(s_65_30), .c(s_65_29), .d(s_65_28), .cin(t_823), .o(t_847), .co(t_848), .cout(t_849));
compressor_4_2 u2_298(.a(s_66_3), .b(s_66_2), .c(s_66_1), .d(s_66_0), .cin(t_828), .o(t_850), .co(t_851), .cout(t_852));
compressor_4_2 u2_299(.a(s_66_7), .b(s_66_6), .c(s_66_5), .d(s_66_4), .cin(t_831), .o(t_853), .co(t_854), .cout(t_855));
compressor_4_2 u2_300(.a(s_66_11), .b(s_66_10), .c(s_66_9), .d(s_66_8), .cin(t_834), .o(t_856), .co(t_857), .cout(t_858));
compressor_4_2 u2_301(.a(s_66_15), .b(s_66_14), .c(s_66_13), .d(s_66_12), .cin(t_837), .o(t_859), .co(t_860), .cout(t_861));
compressor_4_2 u2_302(.a(s_66_19), .b(s_66_18), .c(s_66_17), .d(s_66_16), .cin(t_840), .o(t_862), .co(t_863), .cout(t_864));
compressor_4_2 u2_303(.a(s_66_23), .b(s_66_22), .c(s_66_21), .d(s_66_20), .cin(t_843), .o(t_865), .co(t_866), .cout(t_867));
compressor_4_2 u2_304(.a(s_66_27), .b(s_66_26), .c(s_66_25), .d(s_66_24), .cin(t_846), .o(t_868), .co(t_869), .cout(t_870));
compressor_4_2 u2_305(.a(s_66_31), .b(s_66_30), .c(s_66_29), .d(s_66_28), .cin(t_849), .o(t_871), .co(t_872), .cout(t_873));
compressor_3_2 u1_306(.a(s_66_34), .b(s_66_33), .cin(s_66_32), .o(t_874), .cout(t_875));
compressor_4_2 u2_307(.a(s_67_3), .b(s_67_2), .c(s_67_1), .d(s_67_0), .cin(t_852), .o(t_876), .co(t_877), .cout(t_878));
compressor_4_2 u2_308(.a(s_67_7), .b(s_67_6), .c(s_67_5), .d(s_67_4), .cin(t_855), .o(t_879), .co(t_880), .cout(t_881));
compressor_4_2 u2_309(.a(s_67_11), .b(s_67_10), .c(s_67_9), .d(s_67_8), .cin(t_858), .o(t_882), .co(t_883), .cout(t_884));
compressor_4_2 u2_310(.a(s_67_15), .b(s_67_14), .c(s_67_13), .d(s_67_12), .cin(t_861), .o(t_885), .co(t_886), .cout(t_887));
compressor_4_2 u2_311(.a(s_67_19), .b(s_67_18), .c(s_67_17), .d(s_67_16), .cin(t_864), .o(t_888), .co(t_889), .cout(t_890));
compressor_4_2 u2_312(.a(s_67_23), .b(s_67_22), .c(s_67_21), .d(s_67_20), .cin(t_867), .o(t_891), .co(t_892), .cout(t_893));
compressor_4_2 u2_313(.a(s_67_27), .b(s_67_26), .c(s_67_25), .d(s_67_24), .cin(t_870), .o(t_894), .co(t_895), .cout(t_896));
compressor_4_2 u2_314(.a(s_67_31), .b(s_67_30), .c(s_67_29), .d(s_67_28), .cin(t_873), .o(t_897), .co(t_898), .cout(t_899));
half_adder u0_315(.a(s_67_33), .b(s_67_32), .o(t_900), .cout(t_901));
compressor_4_2 u2_316(.a(s_68_3), .b(s_68_2), .c(s_68_1), .d(s_68_0), .cin(t_878), .o(t_902), .co(t_903), .cout(t_904));
compressor_4_2 u2_317(.a(s_68_7), .b(s_68_6), .c(s_68_5), .d(s_68_4), .cin(t_881), .o(t_905), .co(t_906), .cout(t_907));
compressor_4_2 u2_318(.a(s_68_11), .b(s_68_10), .c(s_68_9), .d(s_68_8), .cin(t_884), .o(t_908), .co(t_909), .cout(t_910));
compressor_4_2 u2_319(.a(s_68_15), .b(s_68_14), .c(s_68_13), .d(s_68_12), .cin(t_887), .o(t_911), .co(t_912), .cout(t_913));
compressor_4_2 u2_320(.a(s_68_19), .b(s_68_18), .c(s_68_17), .d(s_68_16), .cin(t_890), .o(t_914), .co(t_915), .cout(t_916));
compressor_4_2 u2_321(.a(s_68_23), .b(s_68_22), .c(s_68_21), .d(s_68_20), .cin(t_893), .o(t_917), .co(t_918), .cout(t_919));
compressor_4_2 u2_322(.a(s_68_27), .b(s_68_26), .c(s_68_25), .d(s_68_24), .cin(t_896), .o(t_920), .co(t_921), .cout(t_922));
compressor_4_2 u2_323(.a(s_68_31), .b(s_68_30), .c(s_68_29), .d(s_68_28), .cin(t_899), .o(t_923), .co(t_924), .cout(t_925));
compressor_3_2 u1_324(.a(s_68_34), .b(s_68_33), .cin(s_68_32), .o(t_926), .cout(t_927));
compressor_4_2 u2_325(.a(s_69_3), .b(s_69_2), .c(s_69_1), .d(s_69_0), .cin(t_904), .o(t_928), .co(t_929), .cout(t_930));
compressor_4_2 u2_326(.a(s_69_7), .b(s_69_6), .c(s_69_5), .d(s_69_4), .cin(t_907), .o(t_931), .co(t_932), .cout(t_933));
compressor_4_2 u2_327(.a(s_69_11), .b(s_69_10), .c(s_69_9), .d(s_69_8), .cin(t_910), .o(t_934), .co(t_935), .cout(t_936));
compressor_4_2 u2_328(.a(s_69_15), .b(s_69_14), .c(s_69_13), .d(s_69_12), .cin(t_913), .o(t_937), .co(t_938), .cout(t_939));
compressor_4_2 u2_329(.a(s_69_19), .b(s_69_18), .c(s_69_17), .d(s_69_16), .cin(t_916), .o(t_940), .co(t_941), .cout(t_942));
compressor_4_2 u2_330(.a(s_69_23), .b(s_69_22), .c(s_69_21), .d(s_69_20), .cin(t_919), .o(t_943), .co(t_944), .cout(t_945));
compressor_4_2 u2_331(.a(s_69_27), .b(s_69_26), .c(s_69_25), .d(s_69_24), .cin(t_922), .o(t_946), .co(t_947), .cout(t_948));
compressor_4_2 u2_332(.a(s_69_31), .b(s_69_30), .c(s_69_29), .d(s_69_28), .cin(t_925), .o(t_949), .co(t_950), .cout(t_951));
compressor_3_2 u1_333(.a(s_69_34), .b(s_69_33), .cin(s_69_32), .o(t_952), .cout(t_953));
compressor_4_2 u2_334(.a(s_70_3), .b(s_70_2), .c(s_70_1), .d(s_70_0), .cin(t_930), .o(t_954), .co(t_955), .cout(t_956));
compressor_4_2 u2_335(.a(s_70_7), .b(s_70_6), .c(s_70_5), .d(s_70_4), .cin(t_933), .o(t_957), .co(t_958), .cout(t_959));
compressor_4_2 u2_336(.a(s_70_11), .b(s_70_10), .c(s_70_9), .d(s_70_8), .cin(t_936), .o(t_960), .co(t_961), .cout(t_962));
compressor_4_2 u2_337(.a(s_70_15), .b(s_70_14), .c(s_70_13), .d(s_70_12), .cin(t_939), .o(t_963), .co(t_964), .cout(t_965));
compressor_4_2 u2_338(.a(s_70_19), .b(s_70_18), .c(s_70_17), .d(s_70_16), .cin(t_942), .o(t_966), .co(t_967), .cout(t_968));
compressor_4_2 u2_339(.a(s_70_23), .b(s_70_22), .c(s_70_21), .d(s_70_20), .cin(t_945), .o(t_969), .co(t_970), .cout(t_971));
compressor_4_2 u2_340(.a(s_70_27), .b(s_70_26), .c(s_70_25), .d(s_70_24), .cin(t_948), .o(t_972), .co(t_973), .cout(t_974));
compressor_4_2 u2_341(.a(s_70_31), .b(s_70_30), .c(s_70_29), .d(s_70_28), .cin(t_951), .o(t_975), .co(t_976), .cout(t_977));
compressor_4_2 u2_342(.a(s_70_36), .b(s_70_35), .c(s_70_34), .d(s_70_33), .cin(s_70_32), .o(t_978), .co(t_979), .cout(t_980));
compressor_4_2 u2_343(.a(s_71_3), .b(s_71_2), .c(s_71_1), .d(s_71_0), .cin(t_956), .o(t_981), .co(t_982), .cout(t_983));
compressor_4_2 u2_344(.a(s_71_7), .b(s_71_6), .c(s_71_5), .d(s_71_4), .cin(t_959), .o(t_984), .co(t_985), .cout(t_986));
compressor_4_2 u2_345(.a(s_71_11), .b(s_71_10), .c(s_71_9), .d(s_71_8), .cin(t_962), .o(t_987), .co(t_988), .cout(t_989));
compressor_4_2 u2_346(.a(s_71_15), .b(s_71_14), .c(s_71_13), .d(s_71_12), .cin(t_965), .o(t_990), .co(t_991), .cout(t_992));
compressor_4_2 u2_347(.a(s_71_19), .b(s_71_18), .c(s_71_17), .d(s_71_16), .cin(t_968), .o(t_993), .co(t_994), .cout(t_995));
compressor_4_2 u2_348(.a(s_71_23), .b(s_71_22), .c(s_71_21), .d(s_71_20), .cin(t_971), .o(t_996), .co(t_997), .cout(t_998));
compressor_4_2 u2_349(.a(s_71_27), .b(s_71_26), .c(s_71_25), .d(s_71_24), .cin(t_974), .o(t_999), .co(t_1000), .cout(t_1001));
compressor_4_2 u2_350(.a(s_71_31), .b(s_71_30), .c(s_71_29), .d(s_71_28), .cin(t_977), .o(t_1002), .co(t_1003), .cout(t_1004));
compressor_4_2 u2_351(.a(s_71_35), .b(s_71_34), .c(s_71_33), .d(s_71_32), .cin(t_980), .o(t_1005), .co(t_1006), .cout(t_1007));
compressor_4_2 u2_352(.a(s_72_3), .b(s_72_2), .c(s_72_1), .d(s_72_0), .cin(t_983), .o(t_1008), .co(t_1009), .cout(t_1010));
compressor_4_2 u2_353(.a(s_72_7), .b(s_72_6), .c(s_72_5), .d(s_72_4), .cin(t_986), .o(t_1011), .co(t_1012), .cout(t_1013));
compressor_4_2 u2_354(.a(s_72_11), .b(s_72_10), .c(s_72_9), .d(s_72_8), .cin(t_989), .o(t_1014), .co(t_1015), .cout(t_1016));
compressor_4_2 u2_355(.a(s_72_15), .b(s_72_14), .c(s_72_13), .d(s_72_12), .cin(t_992), .o(t_1017), .co(t_1018), .cout(t_1019));
compressor_4_2 u2_356(.a(s_72_19), .b(s_72_18), .c(s_72_17), .d(s_72_16), .cin(t_995), .o(t_1020), .co(t_1021), .cout(t_1022));
compressor_4_2 u2_357(.a(s_72_23), .b(s_72_22), .c(s_72_21), .d(s_72_20), .cin(t_998), .o(t_1023), .co(t_1024), .cout(t_1025));
compressor_4_2 u2_358(.a(s_72_27), .b(s_72_26), .c(s_72_25), .d(s_72_24), .cin(t_1001), .o(t_1026), .co(t_1027), .cout(t_1028));
compressor_4_2 u2_359(.a(s_72_31), .b(s_72_30), .c(s_72_29), .d(s_72_28), .cin(t_1004), .o(t_1029), .co(t_1030), .cout(t_1031));
compressor_4_2 u2_360(.a(s_72_35), .b(s_72_34), .c(s_72_33), .d(s_72_32), .cin(t_1007), .o(t_1032), .co(t_1033), .cout(t_1034));
half_adder u0_361(.a(s_72_37), .b(s_72_36), .o(t_1035), .cout(t_1036));
compressor_4_2 u2_362(.a(s_73_3), .b(s_73_2), .c(s_73_1), .d(s_73_0), .cin(t_1010), .o(t_1037), .co(t_1038), .cout(t_1039));
compressor_4_2 u2_363(.a(s_73_7), .b(s_73_6), .c(s_73_5), .d(s_73_4), .cin(t_1013), .o(t_1040), .co(t_1041), .cout(t_1042));
compressor_4_2 u2_364(.a(s_73_11), .b(s_73_10), .c(s_73_9), .d(s_73_8), .cin(t_1016), .o(t_1043), .co(t_1044), .cout(t_1045));
compressor_4_2 u2_365(.a(s_73_15), .b(s_73_14), .c(s_73_13), .d(s_73_12), .cin(t_1019), .o(t_1046), .co(t_1047), .cout(t_1048));
compressor_4_2 u2_366(.a(s_73_19), .b(s_73_18), .c(s_73_17), .d(s_73_16), .cin(t_1022), .o(t_1049), .co(t_1050), .cout(t_1051));
compressor_4_2 u2_367(.a(s_73_23), .b(s_73_22), .c(s_73_21), .d(s_73_20), .cin(t_1025), .o(t_1052), .co(t_1053), .cout(t_1054));
compressor_4_2 u2_368(.a(s_73_27), .b(s_73_26), .c(s_73_25), .d(s_73_24), .cin(t_1028), .o(t_1055), .co(t_1056), .cout(t_1057));
compressor_4_2 u2_369(.a(s_73_31), .b(s_73_30), .c(s_73_29), .d(s_73_28), .cin(t_1031), .o(t_1058), .co(t_1059), .cout(t_1060));
compressor_4_2 u2_370(.a(s_73_35), .b(s_73_34), .c(s_73_33), .d(s_73_32), .cin(t_1034), .o(t_1061), .co(t_1062), .cout(t_1063));
compressor_4_2 u2_371(.a(s_74_3), .b(s_74_2), .c(s_74_1), .d(s_74_0), .cin(t_1039), .o(t_1064), .co(t_1065), .cout(t_1066));
compressor_4_2 u2_372(.a(s_74_7), .b(s_74_6), .c(s_74_5), .d(s_74_4), .cin(t_1042), .o(t_1067), .co(t_1068), .cout(t_1069));
compressor_4_2 u2_373(.a(s_74_11), .b(s_74_10), .c(s_74_9), .d(s_74_8), .cin(t_1045), .o(t_1070), .co(t_1071), .cout(t_1072));
compressor_4_2 u2_374(.a(s_74_15), .b(s_74_14), .c(s_74_13), .d(s_74_12), .cin(t_1048), .o(t_1073), .co(t_1074), .cout(t_1075));
compressor_4_2 u2_375(.a(s_74_19), .b(s_74_18), .c(s_74_17), .d(s_74_16), .cin(t_1051), .o(t_1076), .co(t_1077), .cout(t_1078));
compressor_4_2 u2_376(.a(s_74_23), .b(s_74_22), .c(s_74_21), .d(s_74_20), .cin(t_1054), .o(t_1079), .co(t_1080), .cout(t_1081));
compressor_4_2 u2_377(.a(s_74_27), .b(s_74_26), .c(s_74_25), .d(s_74_24), .cin(t_1057), .o(t_1082), .co(t_1083), .cout(t_1084));
compressor_4_2 u2_378(.a(s_74_31), .b(s_74_30), .c(s_74_29), .d(s_74_28), .cin(t_1060), .o(t_1085), .co(t_1086), .cout(t_1087));
compressor_4_2 u2_379(.a(s_74_35), .b(s_74_34), .c(s_74_33), .d(s_74_32), .cin(t_1063), .o(t_1088), .co(t_1089), .cout(t_1090));
compressor_3_2 u1_380(.a(s_74_38), .b(s_74_37), .cin(s_74_36), .o(t_1091), .cout(t_1092));
compressor_4_2 u2_381(.a(s_75_3), .b(s_75_2), .c(s_75_1), .d(s_75_0), .cin(t_1066), .o(t_1093), .co(t_1094), .cout(t_1095));
compressor_4_2 u2_382(.a(s_75_7), .b(s_75_6), .c(s_75_5), .d(s_75_4), .cin(t_1069), .o(t_1096), .co(t_1097), .cout(t_1098));
compressor_4_2 u2_383(.a(s_75_11), .b(s_75_10), .c(s_75_9), .d(s_75_8), .cin(t_1072), .o(t_1099), .co(t_1100), .cout(t_1101));
compressor_4_2 u2_384(.a(s_75_15), .b(s_75_14), .c(s_75_13), .d(s_75_12), .cin(t_1075), .o(t_1102), .co(t_1103), .cout(t_1104));
compressor_4_2 u2_385(.a(s_75_19), .b(s_75_18), .c(s_75_17), .d(s_75_16), .cin(t_1078), .o(t_1105), .co(t_1106), .cout(t_1107));
compressor_4_2 u2_386(.a(s_75_23), .b(s_75_22), .c(s_75_21), .d(s_75_20), .cin(t_1081), .o(t_1108), .co(t_1109), .cout(t_1110));
compressor_4_2 u2_387(.a(s_75_27), .b(s_75_26), .c(s_75_25), .d(s_75_24), .cin(t_1084), .o(t_1111), .co(t_1112), .cout(t_1113));
compressor_4_2 u2_388(.a(s_75_31), .b(s_75_30), .c(s_75_29), .d(s_75_28), .cin(t_1087), .o(t_1114), .co(t_1115), .cout(t_1116));
compressor_4_2 u2_389(.a(s_75_35), .b(s_75_34), .c(s_75_33), .d(s_75_32), .cin(t_1090), .o(t_1117), .co(t_1118), .cout(t_1119));
half_adder u0_390(.a(s_75_37), .b(s_75_36), .o(t_1120), .cout(t_1121));
compressor_4_2 u2_391(.a(s_76_3), .b(s_76_2), .c(s_76_1), .d(s_76_0), .cin(t_1095), .o(t_1122), .co(t_1123), .cout(t_1124));
compressor_4_2 u2_392(.a(s_76_7), .b(s_76_6), .c(s_76_5), .d(s_76_4), .cin(t_1098), .o(t_1125), .co(t_1126), .cout(t_1127));
compressor_4_2 u2_393(.a(s_76_11), .b(s_76_10), .c(s_76_9), .d(s_76_8), .cin(t_1101), .o(t_1128), .co(t_1129), .cout(t_1130));
compressor_4_2 u2_394(.a(s_76_15), .b(s_76_14), .c(s_76_13), .d(s_76_12), .cin(t_1104), .o(t_1131), .co(t_1132), .cout(t_1133));
compressor_4_2 u2_395(.a(s_76_19), .b(s_76_18), .c(s_76_17), .d(s_76_16), .cin(t_1107), .o(t_1134), .co(t_1135), .cout(t_1136));
compressor_4_2 u2_396(.a(s_76_23), .b(s_76_22), .c(s_76_21), .d(s_76_20), .cin(t_1110), .o(t_1137), .co(t_1138), .cout(t_1139));
compressor_4_2 u2_397(.a(s_76_27), .b(s_76_26), .c(s_76_25), .d(s_76_24), .cin(t_1113), .o(t_1140), .co(t_1141), .cout(t_1142));
compressor_4_2 u2_398(.a(s_76_31), .b(s_76_30), .c(s_76_29), .d(s_76_28), .cin(t_1116), .o(t_1143), .co(t_1144), .cout(t_1145));
compressor_4_2 u2_399(.a(s_76_35), .b(s_76_34), .c(s_76_33), .d(s_76_32), .cin(t_1119), .o(t_1146), .co(t_1147), .cout(t_1148));
compressor_3_2 u1_400(.a(s_76_38), .b(s_76_37), .cin(s_76_36), .o(t_1149), .cout(t_1150));
compressor_4_2 u2_401(.a(s_77_3), .b(s_77_2), .c(s_77_1), .d(s_77_0), .cin(t_1124), .o(t_1151), .co(t_1152), .cout(t_1153));
compressor_4_2 u2_402(.a(s_77_7), .b(s_77_6), .c(s_77_5), .d(s_77_4), .cin(t_1127), .o(t_1154), .co(t_1155), .cout(t_1156));
compressor_4_2 u2_403(.a(s_77_11), .b(s_77_10), .c(s_77_9), .d(s_77_8), .cin(t_1130), .o(t_1157), .co(t_1158), .cout(t_1159));
compressor_4_2 u2_404(.a(s_77_15), .b(s_77_14), .c(s_77_13), .d(s_77_12), .cin(t_1133), .o(t_1160), .co(t_1161), .cout(t_1162));
compressor_4_2 u2_405(.a(s_77_19), .b(s_77_18), .c(s_77_17), .d(s_77_16), .cin(t_1136), .o(t_1163), .co(t_1164), .cout(t_1165));
compressor_4_2 u2_406(.a(s_77_23), .b(s_77_22), .c(s_77_21), .d(s_77_20), .cin(t_1139), .o(t_1166), .co(t_1167), .cout(t_1168));
compressor_4_2 u2_407(.a(s_77_27), .b(s_77_26), .c(s_77_25), .d(s_77_24), .cin(t_1142), .o(t_1169), .co(t_1170), .cout(t_1171));
compressor_4_2 u2_408(.a(s_77_31), .b(s_77_30), .c(s_77_29), .d(s_77_28), .cin(t_1145), .o(t_1172), .co(t_1173), .cout(t_1174));
compressor_4_2 u2_409(.a(s_77_35), .b(s_77_34), .c(s_77_33), .d(s_77_32), .cin(t_1148), .o(t_1175), .co(t_1176), .cout(t_1177));
compressor_3_2 u1_410(.a(s_77_38), .b(s_77_37), .cin(s_77_36), .o(t_1178), .cout(t_1179));
compressor_4_2 u2_411(.a(s_78_3), .b(s_78_2), .c(s_78_1), .d(s_78_0), .cin(t_1153), .o(t_1180), .co(t_1181), .cout(t_1182));
compressor_4_2 u2_412(.a(s_78_7), .b(s_78_6), .c(s_78_5), .d(s_78_4), .cin(t_1156), .o(t_1183), .co(t_1184), .cout(t_1185));
compressor_4_2 u2_413(.a(s_78_11), .b(s_78_10), .c(s_78_9), .d(s_78_8), .cin(t_1159), .o(t_1186), .co(t_1187), .cout(t_1188));
compressor_4_2 u2_414(.a(s_78_15), .b(s_78_14), .c(s_78_13), .d(s_78_12), .cin(t_1162), .o(t_1189), .co(t_1190), .cout(t_1191));
compressor_4_2 u2_415(.a(s_78_19), .b(s_78_18), .c(s_78_17), .d(s_78_16), .cin(t_1165), .o(t_1192), .co(t_1193), .cout(t_1194));
compressor_4_2 u2_416(.a(s_78_23), .b(s_78_22), .c(s_78_21), .d(s_78_20), .cin(t_1168), .o(t_1195), .co(t_1196), .cout(t_1197));
compressor_4_2 u2_417(.a(s_78_27), .b(s_78_26), .c(s_78_25), .d(s_78_24), .cin(t_1171), .o(t_1198), .co(t_1199), .cout(t_1200));
compressor_4_2 u2_418(.a(s_78_31), .b(s_78_30), .c(s_78_29), .d(s_78_28), .cin(t_1174), .o(t_1201), .co(t_1202), .cout(t_1203));
compressor_4_2 u2_419(.a(s_78_35), .b(s_78_34), .c(s_78_33), .d(s_78_32), .cin(t_1177), .o(t_1204), .co(t_1205), .cout(t_1206));
compressor_4_2 u2_420(.a(s_78_40), .b(s_78_39), .c(s_78_38), .d(s_78_37), .cin(s_78_36), .o(t_1207), .co(t_1208), .cout(t_1209));
compressor_4_2 u2_421(.a(s_79_3), .b(s_79_2), .c(s_79_1), .d(s_79_0), .cin(t_1182), .o(t_1210), .co(t_1211), .cout(t_1212));
compressor_4_2 u2_422(.a(s_79_7), .b(s_79_6), .c(s_79_5), .d(s_79_4), .cin(t_1185), .o(t_1213), .co(t_1214), .cout(t_1215));
compressor_4_2 u2_423(.a(s_79_11), .b(s_79_10), .c(s_79_9), .d(s_79_8), .cin(t_1188), .o(t_1216), .co(t_1217), .cout(t_1218));
compressor_4_2 u2_424(.a(s_79_15), .b(s_79_14), .c(s_79_13), .d(s_79_12), .cin(t_1191), .o(t_1219), .co(t_1220), .cout(t_1221));
compressor_4_2 u2_425(.a(s_79_19), .b(s_79_18), .c(s_79_17), .d(s_79_16), .cin(t_1194), .o(t_1222), .co(t_1223), .cout(t_1224));
compressor_4_2 u2_426(.a(s_79_23), .b(s_79_22), .c(s_79_21), .d(s_79_20), .cin(t_1197), .o(t_1225), .co(t_1226), .cout(t_1227));
compressor_4_2 u2_427(.a(s_79_27), .b(s_79_26), .c(s_79_25), .d(s_79_24), .cin(t_1200), .o(t_1228), .co(t_1229), .cout(t_1230));
compressor_4_2 u2_428(.a(s_79_31), .b(s_79_30), .c(s_79_29), .d(s_79_28), .cin(t_1203), .o(t_1231), .co(t_1232), .cout(t_1233));
compressor_4_2 u2_429(.a(s_79_35), .b(s_79_34), .c(s_79_33), .d(s_79_32), .cin(t_1206), .o(t_1234), .co(t_1235), .cout(t_1236));
compressor_4_2 u2_430(.a(s_79_39), .b(s_79_38), .c(s_79_37), .d(s_79_36), .cin(t_1209), .o(t_1237), .co(t_1238), .cout(t_1239));
compressor_4_2 u2_431(.a(s_80_3), .b(s_80_2), .c(s_80_1), .d(s_80_0), .cin(t_1212), .o(t_1240), .co(t_1241), .cout(t_1242));
compressor_4_2 u2_432(.a(s_80_7), .b(s_80_6), .c(s_80_5), .d(s_80_4), .cin(t_1215), .o(t_1243), .co(t_1244), .cout(t_1245));
compressor_4_2 u2_433(.a(s_80_11), .b(s_80_10), .c(s_80_9), .d(s_80_8), .cin(t_1218), .o(t_1246), .co(t_1247), .cout(t_1248));
compressor_4_2 u2_434(.a(s_80_15), .b(s_80_14), .c(s_80_13), .d(s_80_12), .cin(t_1221), .o(t_1249), .co(t_1250), .cout(t_1251));
compressor_4_2 u2_435(.a(s_80_19), .b(s_80_18), .c(s_80_17), .d(s_80_16), .cin(t_1224), .o(t_1252), .co(t_1253), .cout(t_1254));
compressor_4_2 u2_436(.a(s_80_23), .b(s_80_22), .c(s_80_21), .d(s_80_20), .cin(t_1227), .o(t_1255), .co(t_1256), .cout(t_1257));
compressor_4_2 u2_437(.a(s_80_27), .b(s_80_26), .c(s_80_25), .d(s_80_24), .cin(t_1230), .o(t_1258), .co(t_1259), .cout(t_1260));
compressor_4_2 u2_438(.a(s_80_31), .b(s_80_30), .c(s_80_29), .d(s_80_28), .cin(t_1233), .o(t_1261), .co(t_1262), .cout(t_1263));
compressor_4_2 u2_439(.a(s_80_35), .b(s_80_34), .c(s_80_33), .d(s_80_32), .cin(t_1236), .o(t_1264), .co(t_1265), .cout(t_1266));
compressor_4_2 u2_440(.a(s_80_39), .b(s_80_38), .c(s_80_37), .d(s_80_36), .cin(t_1239), .o(t_1267), .co(t_1268), .cout(t_1269));
half_adder u0_441(.a(s_80_41), .b(s_80_40), .o(t_1270), .cout(t_1271));
compressor_4_2 u2_442(.a(s_81_3), .b(s_81_2), .c(s_81_1), .d(s_81_0), .cin(t_1242), .o(t_1272), .co(t_1273), .cout(t_1274));
compressor_4_2 u2_443(.a(s_81_7), .b(s_81_6), .c(s_81_5), .d(s_81_4), .cin(t_1245), .o(t_1275), .co(t_1276), .cout(t_1277));
compressor_4_2 u2_444(.a(s_81_11), .b(s_81_10), .c(s_81_9), .d(s_81_8), .cin(t_1248), .o(t_1278), .co(t_1279), .cout(t_1280));
compressor_4_2 u2_445(.a(s_81_15), .b(s_81_14), .c(s_81_13), .d(s_81_12), .cin(t_1251), .o(t_1281), .co(t_1282), .cout(t_1283));
compressor_4_2 u2_446(.a(s_81_19), .b(s_81_18), .c(s_81_17), .d(s_81_16), .cin(t_1254), .o(t_1284), .co(t_1285), .cout(t_1286));
compressor_4_2 u2_447(.a(s_81_23), .b(s_81_22), .c(s_81_21), .d(s_81_20), .cin(t_1257), .o(t_1287), .co(t_1288), .cout(t_1289));
compressor_4_2 u2_448(.a(s_81_27), .b(s_81_26), .c(s_81_25), .d(s_81_24), .cin(t_1260), .o(t_1290), .co(t_1291), .cout(t_1292));
compressor_4_2 u2_449(.a(s_81_31), .b(s_81_30), .c(s_81_29), .d(s_81_28), .cin(t_1263), .o(t_1293), .co(t_1294), .cout(t_1295));
compressor_4_2 u2_450(.a(s_81_35), .b(s_81_34), .c(s_81_33), .d(s_81_32), .cin(t_1266), .o(t_1296), .co(t_1297), .cout(t_1298));
compressor_4_2 u2_451(.a(s_81_39), .b(s_81_38), .c(s_81_37), .d(s_81_36), .cin(t_1269), .o(t_1299), .co(t_1300), .cout(t_1301));
compressor_4_2 u2_452(.a(s_82_3), .b(s_82_2), .c(s_82_1), .d(s_82_0), .cin(t_1274), .o(t_1302), .co(t_1303), .cout(t_1304));
compressor_4_2 u2_453(.a(s_82_7), .b(s_82_6), .c(s_82_5), .d(s_82_4), .cin(t_1277), .o(t_1305), .co(t_1306), .cout(t_1307));
compressor_4_2 u2_454(.a(s_82_11), .b(s_82_10), .c(s_82_9), .d(s_82_8), .cin(t_1280), .o(t_1308), .co(t_1309), .cout(t_1310));
compressor_4_2 u2_455(.a(s_82_15), .b(s_82_14), .c(s_82_13), .d(s_82_12), .cin(t_1283), .o(t_1311), .co(t_1312), .cout(t_1313));
compressor_4_2 u2_456(.a(s_82_19), .b(s_82_18), .c(s_82_17), .d(s_82_16), .cin(t_1286), .o(t_1314), .co(t_1315), .cout(t_1316));
compressor_4_2 u2_457(.a(s_82_23), .b(s_82_22), .c(s_82_21), .d(s_82_20), .cin(t_1289), .o(t_1317), .co(t_1318), .cout(t_1319));
compressor_4_2 u2_458(.a(s_82_27), .b(s_82_26), .c(s_82_25), .d(s_82_24), .cin(t_1292), .o(t_1320), .co(t_1321), .cout(t_1322));
compressor_4_2 u2_459(.a(s_82_31), .b(s_82_30), .c(s_82_29), .d(s_82_28), .cin(t_1295), .o(t_1323), .co(t_1324), .cout(t_1325));
compressor_4_2 u2_460(.a(s_82_35), .b(s_82_34), .c(s_82_33), .d(s_82_32), .cin(t_1298), .o(t_1326), .co(t_1327), .cout(t_1328));
compressor_4_2 u2_461(.a(s_82_39), .b(s_82_38), .c(s_82_37), .d(s_82_36), .cin(t_1301), .o(t_1329), .co(t_1330), .cout(t_1331));
compressor_3_2 u1_462(.a(s_82_42), .b(s_82_41), .cin(s_82_40), .o(t_1332), .cout(t_1333));
compressor_4_2 u2_463(.a(s_83_3), .b(s_83_2), .c(s_83_1), .d(s_83_0), .cin(t_1304), .o(t_1334), .co(t_1335), .cout(t_1336));
compressor_4_2 u2_464(.a(s_83_7), .b(s_83_6), .c(s_83_5), .d(s_83_4), .cin(t_1307), .o(t_1337), .co(t_1338), .cout(t_1339));
compressor_4_2 u2_465(.a(s_83_11), .b(s_83_10), .c(s_83_9), .d(s_83_8), .cin(t_1310), .o(t_1340), .co(t_1341), .cout(t_1342));
compressor_4_2 u2_466(.a(s_83_15), .b(s_83_14), .c(s_83_13), .d(s_83_12), .cin(t_1313), .o(t_1343), .co(t_1344), .cout(t_1345));
compressor_4_2 u2_467(.a(s_83_19), .b(s_83_18), .c(s_83_17), .d(s_83_16), .cin(t_1316), .o(t_1346), .co(t_1347), .cout(t_1348));
compressor_4_2 u2_468(.a(s_83_23), .b(s_83_22), .c(s_83_21), .d(s_83_20), .cin(t_1319), .o(t_1349), .co(t_1350), .cout(t_1351));
compressor_4_2 u2_469(.a(s_83_27), .b(s_83_26), .c(s_83_25), .d(s_83_24), .cin(t_1322), .o(t_1352), .co(t_1353), .cout(t_1354));
compressor_4_2 u2_470(.a(s_83_31), .b(s_83_30), .c(s_83_29), .d(s_83_28), .cin(t_1325), .o(t_1355), .co(t_1356), .cout(t_1357));
compressor_4_2 u2_471(.a(s_83_35), .b(s_83_34), .c(s_83_33), .d(s_83_32), .cin(t_1328), .o(t_1358), .co(t_1359), .cout(t_1360));
compressor_4_2 u2_472(.a(s_83_39), .b(s_83_38), .c(s_83_37), .d(s_83_36), .cin(t_1331), .o(t_1361), .co(t_1362), .cout(t_1363));
half_adder u0_473(.a(s_83_41), .b(s_83_40), .o(t_1364), .cout(t_1365));
compressor_4_2 u2_474(.a(s_84_3), .b(s_84_2), .c(s_84_1), .d(s_84_0), .cin(t_1336), .o(t_1366), .co(t_1367), .cout(t_1368));
compressor_4_2 u2_475(.a(s_84_7), .b(s_84_6), .c(s_84_5), .d(s_84_4), .cin(t_1339), .o(t_1369), .co(t_1370), .cout(t_1371));
compressor_4_2 u2_476(.a(s_84_11), .b(s_84_10), .c(s_84_9), .d(s_84_8), .cin(t_1342), .o(t_1372), .co(t_1373), .cout(t_1374));
compressor_4_2 u2_477(.a(s_84_15), .b(s_84_14), .c(s_84_13), .d(s_84_12), .cin(t_1345), .o(t_1375), .co(t_1376), .cout(t_1377));
compressor_4_2 u2_478(.a(s_84_19), .b(s_84_18), .c(s_84_17), .d(s_84_16), .cin(t_1348), .o(t_1378), .co(t_1379), .cout(t_1380));
compressor_4_2 u2_479(.a(s_84_23), .b(s_84_22), .c(s_84_21), .d(s_84_20), .cin(t_1351), .o(t_1381), .co(t_1382), .cout(t_1383));
compressor_4_2 u2_480(.a(s_84_27), .b(s_84_26), .c(s_84_25), .d(s_84_24), .cin(t_1354), .o(t_1384), .co(t_1385), .cout(t_1386));
compressor_4_2 u2_481(.a(s_84_31), .b(s_84_30), .c(s_84_29), .d(s_84_28), .cin(t_1357), .o(t_1387), .co(t_1388), .cout(t_1389));
compressor_4_2 u2_482(.a(s_84_35), .b(s_84_34), .c(s_84_33), .d(s_84_32), .cin(t_1360), .o(t_1390), .co(t_1391), .cout(t_1392));
compressor_4_2 u2_483(.a(s_84_39), .b(s_84_38), .c(s_84_37), .d(s_84_36), .cin(t_1363), .o(t_1393), .co(t_1394), .cout(t_1395));
compressor_3_2 u1_484(.a(s_84_42), .b(s_84_41), .cin(s_84_40), .o(t_1396), .cout(t_1397));
compressor_4_2 u2_485(.a(s_85_3), .b(s_85_2), .c(s_85_1), .d(s_85_0), .cin(t_1368), .o(t_1398), .co(t_1399), .cout(t_1400));
compressor_4_2 u2_486(.a(s_85_7), .b(s_85_6), .c(s_85_5), .d(s_85_4), .cin(t_1371), .o(t_1401), .co(t_1402), .cout(t_1403));
compressor_4_2 u2_487(.a(s_85_11), .b(s_85_10), .c(s_85_9), .d(s_85_8), .cin(t_1374), .o(t_1404), .co(t_1405), .cout(t_1406));
compressor_4_2 u2_488(.a(s_85_15), .b(s_85_14), .c(s_85_13), .d(s_85_12), .cin(t_1377), .o(t_1407), .co(t_1408), .cout(t_1409));
compressor_4_2 u2_489(.a(s_85_19), .b(s_85_18), .c(s_85_17), .d(s_85_16), .cin(t_1380), .o(t_1410), .co(t_1411), .cout(t_1412));
compressor_4_2 u2_490(.a(s_85_23), .b(s_85_22), .c(s_85_21), .d(s_85_20), .cin(t_1383), .o(t_1413), .co(t_1414), .cout(t_1415));
compressor_4_2 u2_491(.a(s_85_27), .b(s_85_26), .c(s_85_25), .d(s_85_24), .cin(t_1386), .o(t_1416), .co(t_1417), .cout(t_1418));
compressor_4_2 u2_492(.a(s_85_31), .b(s_85_30), .c(s_85_29), .d(s_85_28), .cin(t_1389), .o(t_1419), .co(t_1420), .cout(t_1421));
compressor_4_2 u2_493(.a(s_85_35), .b(s_85_34), .c(s_85_33), .d(s_85_32), .cin(t_1392), .o(t_1422), .co(t_1423), .cout(t_1424));
compressor_4_2 u2_494(.a(s_85_39), .b(s_85_38), .c(s_85_37), .d(s_85_36), .cin(t_1395), .o(t_1425), .co(t_1426), .cout(t_1427));
compressor_3_2 u1_495(.a(s_85_42), .b(s_85_41), .cin(s_85_40), .o(t_1428), .cout(t_1429));
compressor_4_2 u2_496(.a(s_86_3), .b(s_86_2), .c(s_86_1), .d(s_86_0), .cin(t_1400), .o(t_1430), .co(t_1431), .cout(t_1432));
compressor_4_2 u2_497(.a(s_86_7), .b(s_86_6), .c(s_86_5), .d(s_86_4), .cin(t_1403), .o(t_1433), .co(t_1434), .cout(t_1435));
compressor_4_2 u2_498(.a(s_86_11), .b(s_86_10), .c(s_86_9), .d(s_86_8), .cin(t_1406), .o(t_1436), .co(t_1437), .cout(t_1438));
compressor_4_2 u2_499(.a(s_86_15), .b(s_86_14), .c(s_86_13), .d(s_86_12), .cin(t_1409), .o(t_1439), .co(t_1440), .cout(t_1441));
compressor_4_2 u2_500(.a(s_86_19), .b(s_86_18), .c(s_86_17), .d(s_86_16), .cin(t_1412), .o(t_1442), .co(t_1443), .cout(t_1444));
compressor_4_2 u2_501(.a(s_86_23), .b(s_86_22), .c(s_86_21), .d(s_86_20), .cin(t_1415), .o(t_1445), .co(t_1446), .cout(t_1447));
compressor_4_2 u2_502(.a(s_86_27), .b(s_86_26), .c(s_86_25), .d(s_86_24), .cin(t_1418), .o(t_1448), .co(t_1449), .cout(t_1450));
compressor_4_2 u2_503(.a(s_86_31), .b(s_86_30), .c(s_86_29), .d(s_86_28), .cin(t_1421), .o(t_1451), .co(t_1452), .cout(t_1453));
compressor_4_2 u2_504(.a(s_86_35), .b(s_86_34), .c(s_86_33), .d(s_86_32), .cin(t_1424), .o(t_1454), .co(t_1455), .cout(t_1456));
compressor_4_2 u2_505(.a(s_86_39), .b(s_86_38), .c(s_86_37), .d(s_86_36), .cin(t_1427), .o(t_1457), .co(t_1458), .cout(t_1459));
compressor_4_2 u2_506(.a(s_86_44), .b(s_86_43), .c(s_86_42), .d(s_86_41), .cin(s_86_40), .o(t_1460), .co(t_1461), .cout(t_1462));
compressor_4_2 u2_507(.a(s_87_3), .b(s_87_2), .c(s_87_1), .d(s_87_0), .cin(t_1432), .o(t_1463), .co(t_1464), .cout(t_1465));
compressor_4_2 u2_508(.a(s_87_7), .b(s_87_6), .c(s_87_5), .d(s_87_4), .cin(t_1435), .o(t_1466), .co(t_1467), .cout(t_1468));
compressor_4_2 u2_509(.a(s_87_11), .b(s_87_10), .c(s_87_9), .d(s_87_8), .cin(t_1438), .o(t_1469), .co(t_1470), .cout(t_1471));
compressor_4_2 u2_510(.a(s_87_15), .b(s_87_14), .c(s_87_13), .d(s_87_12), .cin(t_1441), .o(t_1472), .co(t_1473), .cout(t_1474));
compressor_4_2 u2_511(.a(s_87_19), .b(s_87_18), .c(s_87_17), .d(s_87_16), .cin(t_1444), .o(t_1475), .co(t_1476), .cout(t_1477));
compressor_4_2 u2_512(.a(s_87_23), .b(s_87_22), .c(s_87_21), .d(s_87_20), .cin(t_1447), .o(t_1478), .co(t_1479), .cout(t_1480));
compressor_4_2 u2_513(.a(s_87_27), .b(s_87_26), .c(s_87_25), .d(s_87_24), .cin(t_1450), .o(t_1481), .co(t_1482), .cout(t_1483));
compressor_4_2 u2_514(.a(s_87_31), .b(s_87_30), .c(s_87_29), .d(s_87_28), .cin(t_1453), .o(t_1484), .co(t_1485), .cout(t_1486));
compressor_4_2 u2_515(.a(s_87_35), .b(s_87_34), .c(s_87_33), .d(s_87_32), .cin(t_1456), .o(t_1487), .co(t_1488), .cout(t_1489));
compressor_4_2 u2_516(.a(s_87_39), .b(s_87_38), .c(s_87_37), .d(s_87_36), .cin(t_1459), .o(t_1490), .co(t_1491), .cout(t_1492));
compressor_4_2 u2_517(.a(s_87_43), .b(s_87_42), .c(s_87_41), .d(s_87_40), .cin(t_1462), .o(t_1493), .co(t_1494), .cout(t_1495));
compressor_4_2 u2_518(.a(s_88_3), .b(s_88_2), .c(s_88_1), .d(s_88_0), .cin(t_1465), .o(t_1496), .co(t_1497), .cout(t_1498));
compressor_4_2 u2_519(.a(s_88_7), .b(s_88_6), .c(s_88_5), .d(s_88_4), .cin(t_1468), .o(t_1499), .co(t_1500), .cout(t_1501));
compressor_4_2 u2_520(.a(s_88_11), .b(s_88_10), .c(s_88_9), .d(s_88_8), .cin(t_1471), .o(t_1502), .co(t_1503), .cout(t_1504));
compressor_4_2 u2_521(.a(s_88_15), .b(s_88_14), .c(s_88_13), .d(s_88_12), .cin(t_1474), .o(t_1505), .co(t_1506), .cout(t_1507));
compressor_4_2 u2_522(.a(s_88_19), .b(s_88_18), .c(s_88_17), .d(s_88_16), .cin(t_1477), .o(t_1508), .co(t_1509), .cout(t_1510));
compressor_4_2 u2_523(.a(s_88_23), .b(s_88_22), .c(s_88_21), .d(s_88_20), .cin(t_1480), .o(t_1511), .co(t_1512), .cout(t_1513));
compressor_4_2 u2_524(.a(s_88_27), .b(s_88_26), .c(s_88_25), .d(s_88_24), .cin(t_1483), .o(t_1514), .co(t_1515), .cout(t_1516));
compressor_4_2 u2_525(.a(s_88_31), .b(s_88_30), .c(s_88_29), .d(s_88_28), .cin(t_1486), .o(t_1517), .co(t_1518), .cout(t_1519));
compressor_4_2 u2_526(.a(s_88_35), .b(s_88_34), .c(s_88_33), .d(s_88_32), .cin(t_1489), .o(t_1520), .co(t_1521), .cout(t_1522));
compressor_4_2 u2_527(.a(s_88_39), .b(s_88_38), .c(s_88_37), .d(s_88_36), .cin(t_1492), .o(t_1523), .co(t_1524), .cout(t_1525));
compressor_4_2 u2_528(.a(s_88_43), .b(s_88_42), .c(s_88_41), .d(s_88_40), .cin(t_1495), .o(t_1526), .co(t_1527), .cout(t_1528));
half_adder u0_529(.a(s_88_45), .b(s_88_44), .o(t_1529), .cout(t_1530));
compressor_4_2 u2_530(.a(s_89_3), .b(s_89_2), .c(s_89_1), .d(s_89_0), .cin(t_1498), .o(t_1531), .co(t_1532), .cout(t_1533));
compressor_4_2 u2_531(.a(s_89_7), .b(s_89_6), .c(s_89_5), .d(s_89_4), .cin(t_1501), .o(t_1534), .co(t_1535), .cout(t_1536));
compressor_4_2 u2_532(.a(s_89_11), .b(s_89_10), .c(s_89_9), .d(s_89_8), .cin(t_1504), .o(t_1537), .co(t_1538), .cout(t_1539));
compressor_4_2 u2_533(.a(s_89_15), .b(s_89_14), .c(s_89_13), .d(s_89_12), .cin(t_1507), .o(t_1540), .co(t_1541), .cout(t_1542));
compressor_4_2 u2_534(.a(s_89_19), .b(s_89_18), .c(s_89_17), .d(s_89_16), .cin(t_1510), .o(t_1543), .co(t_1544), .cout(t_1545));
compressor_4_2 u2_535(.a(s_89_23), .b(s_89_22), .c(s_89_21), .d(s_89_20), .cin(t_1513), .o(t_1546), .co(t_1547), .cout(t_1548));
compressor_4_2 u2_536(.a(s_89_27), .b(s_89_26), .c(s_89_25), .d(s_89_24), .cin(t_1516), .o(t_1549), .co(t_1550), .cout(t_1551));
compressor_4_2 u2_537(.a(s_89_31), .b(s_89_30), .c(s_89_29), .d(s_89_28), .cin(t_1519), .o(t_1552), .co(t_1553), .cout(t_1554));
compressor_4_2 u2_538(.a(s_89_35), .b(s_89_34), .c(s_89_33), .d(s_89_32), .cin(t_1522), .o(t_1555), .co(t_1556), .cout(t_1557));
compressor_4_2 u2_539(.a(s_89_39), .b(s_89_38), .c(s_89_37), .d(s_89_36), .cin(t_1525), .o(t_1558), .co(t_1559), .cout(t_1560));
compressor_4_2 u2_540(.a(s_89_43), .b(s_89_42), .c(s_89_41), .d(s_89_40), .cin(t_1528), .o(t_1561), .co(t_1562), .cout(t_1563));
compressor_4_2 u2_541(.a(s_90_3), .b(s_90_2), .c(s_90_1), .d(s_90_0), .cin(t_1533), .o(t_1564), .co(t_1565), .cout(t_1566));
compressor_4_2 u2_542(.a(s_90_7), .b(s_90_6), .c(s_90_5), .d(s_90_4), .cin(t_1536), .o(t_1567), .co(t_1568), .cout(t_1569));
compressor_4_2 u2_543(.a(s_90_11), .b(s_90_10), .c(s_90_9), .d(s_90_8), .cin(t_1539), .o(t_1570), .co(t_1571), .cout(t_1572));
compressor_4_2 u2_544(.a(s_90_15), .b(s_90_14), .c(s_90_13), .d(s_90_12), .cin(t_1542), .o(t_1573), .co(t_1574), .cout(t_1575));
compressor_4_2 u2_545(.a(s_90_19), .b(s_90_18), .c(s_90_17), .d(s_90_16), .cin(t_1545), .o(t_1576), .co(t_1577), .cout(t_1578));
compressor_4_2 u2_546(.a(s_90_23), .b(s_90_22), .c(s_90_21), .d(s_90_20), .cin(t_1548), .o(t_1579), .co(t_1580), .cout(t_1581));
compressor_4_2 u2_547(.a(s_90_27), .b(s_90_26), .c(s_90_25), .d(s_90_24), .cin(t_1551), .o(t_1582), .co(t_1583), .cout(t_1584));
compressor_4_2 u2_548(.a(s_90_31), .b(s_90_30), .c(s_90_29), .d(s_90_28), .cin(t_1554), .o(t_1585), .co(t_1586), .cout(t_1587));
compressor_4_2 u2_549(.a(s_90_35), .b(s_90_34), .c(s_90_33), .d(s_90_32), .cin(t_1557), .o(t_1588), .co(t_1589), .cout(t_1590));
compressor_4_2 u2_550(.a(s_90_39), .b(s_90_38), .c(s_90_37), .d(s_90_36), .cin(t_1560), .o(t_1591), .co(t_1592), .cout(t_1593));
compressor_4_2 u2_551(.a(s_90_43), .b(s_90_42), .c(s_90_41), .d(s_90_40), .cin(t_1563), .o(t_1594), .co(t_1595), .cout(t_1596));
compressor_3_2 u1_552(.a(s_90_46), .b(s_90_45), .cin(s_90_44), .o(t_1597), .cout(t_1598));
compressor_4_2 u2_553(.a(s_91_3), .b(s_91_2), .c(s_91_1), .d(s_91_0), .cin(t_1566), .o(t_1599), .co(t_1600), .cout(t_1601));
compressor_4_2 u2_554(.a(s_91_7), .b(s_91_6), .c(s_91_5), .d(s_91_4), .cin(t_1569), .o(t_1602), .co(t_1603), .cout(t_1604));
compressor_4_2 u2_555(.a(s_91_11), .b(s_91_10), .c(s_91_9), .d(s_91_8), .cin(t_1572), .o(t_1605), .co(t_1606), .cout(t_1607));
compressor_4_2 u2_556(.a(s_91_15), .b(s_91_14), .c(s_91_13), .d(s_91_12), .cin(t_1575), .o(t_1608), .co(t_1609), .cout(t_1610));
compressor_4_2 u2_557(.a(s_91_19), .b(s_91_18), .c(s_91_17), .d(s_91_16), .cin(t_1578), .o(t_1611), .co(t_1612), .cout(t_1613));
compressor_4_2 u2_558(.a(s_91_23), .b(s_91_22), .c(s_91_21), .d(s_91_20), .cin(t_1581), .o(t_1614), .co(t_1615), .cout(t_1616));
compressor_4_2 u2_559(.a(s_91_27), .b(s_91_26), .c(s_91_25), .d(s_91_24), .cin(t_1584), .o(t_1617), .co(t_1618), .cout(t_1619));
compressor_4_2 u2_560(.a(s_91_31), .b(s_91_30), .c(s_91_29), .d(s_91_28), .cin(t_1587), .o(t_1620), .co(t_1621), .cout(t_1622));
compressor_4_2 u2_561(.a(s_91_35), .b(s_91_34), .c(s_91_33), .d(s_91_32), .cin(t_1590), .o(t_1623), .co(t_1624), .cout(t_1625));
compressor_4_2 u2_562(.a(s_91_39), .b(s_91_38), .c(s_91_37), .d(s_91_36), .cin(t_1593), .o(t_1626), .co(t_1627), .cout(t_1628));
compressor_4_2 u2_563(.a(s_91_43), .b(s_91_42), .c(s_91_41), .d(s_91_40), .cin(t_1596), .o(t_1629), .co(t_1630), .cout(t_1631));
half_adder u0_564(.a(s_91_45), .b(s_91_44), .o(t_1632), .cout(t_1633));
compressor_4_2 u2_565(.a(s_92_3), .b(s_92_2), .c(s_92_1), .d(s_92_0), .cin(t_1601), .o(t_1634), .co(t_1635), .cout(t_1636));
compressor_4_2 u2_566(.a(s_92_7), .b(s_92_6), .c(s_92_5), .d(s_92_4), .cin(t_1604), .o(t_1637), .co(t_1638), .cout(t_1639));
compressor_4_2 u2_567(.a(s_92_11), .b(s_92_10), .c(s_92_9), .d(s_92_8), .cin(t_1607), .o(t_1640), .co(t_1641), .cout(t_1642));
compressor_4_2 u2_568(.a(s_92_15), .b(s_92_14), .c(s_92_13), .d(s_92_12), .cin(t_1610), .o(t_1643), .co(t_1644), .cout(t_1645));
compressor_4_2 u2_569(.a(s_92_19), .b(s_92_18), .c(s_92_17), .d(s_92_16), .cin(t_1613), .o(t_1646), .co(t_1647), .cout(t_1648));
compressor_4_2 u2_570(.a(s_92_23), .b(s_92_22), .c(s_92_21), .d(s_92_20), .cin(t_1616), .o(t_1649), .co(t_1650), .cout(t_1651));
compressor_4_2 u2_571(.a(s_92_27), .b(s_92_26), .c(s_92_25), .d(s_92_24), .cin(t_1619), .o(t_1652), .co(t_1653), .cout(t_1654));
compressor_4_2 u2_572(.a(s_92_31), .b(s_92_30), .c(s_92_29), .d(s_92_28), .cin(t_1622), .o(t_1655), .co(t_1656), .cout(t_1657));
compressor_4_2 u2_573(.a(s_92_35), .b(s_92_34), .c(s_92_33), .d(s_92_32), .cin(t_1625), .o(t_1658), .co(t_1659), .cout(t_1660));
compressor_4_2 u2_574(.a(s_92_39), .b(s_92_38), .c(s_92_37), .d(s_92_36), .cin(t_1628), .o(t_1661), .co(t_1662), .cout(t_1663));
compressor_4_2 u2_575(.a(s_92_43), .b(s_92_42), .c(s_92_41), .d(s_92_40), .cin(t_1631), .o(t_1664), .co(t_1665), .cout(t_1666));
compressor_3_2 u1_576(.a(s_92_46), .b(s_92_45), .cin(s_92_44), .o(t_1667), .cout(t_1668));
compressor_4_2 u2_577(.a(s_93_3), .b(s_93_2), .c(s_93_1), .d(s_93_0), .cin(t_1636), .o(t_1669), .co(t_1670), .cout(t_1671));
compressor_4_2 u2_578(.a(s_93_7), .b(s_93_6), .c(s_93_5), .d(s_93_4), .cin(t_1639), .o(t_1672), .co(t_1673), .cout(t_1674));
compressor_4_2 u2_579(.a(s_93_11), .b(s_93_10), .c(s_93_9), .d(s_93_8), .cin(t_1642), .o(t_1675), .co(t_1676), .cout(t_1677));
compressor_4_2 u2_580(.a(s_93_15), .b(s_93_14), .c(s_93_13), .d(s_93_12), .cin(t_1645), .o(t_1678), .co(t_1679), .cout(t_1680));
compressor_4_2 u2_581(.a(s_93_19), .b(s_93_18), .c(s_93_17), .d(s_93_16), .cin(t_1648), .o(t_1681), .co(t_1682), .cout(t_1683));
compressor_4_2 u2_582(.a(s_93_23), .b(s_93_22), .c(s_93_21), .d(s_93_20), .cin(t_1651), .o(t_1684), .co(t_1685), .cout(t_1686));
compressor_4_2 u2_583(.a(s_93_27), .b(s_93_26), .c(s_93_25), .d(s_93_24), .cin(t_1654), .o(t_1687), .co(t_1688), .cout(t_1689));
compressor_4_2 u2_584(.a(s_93_31), .b(s_93_30), .c(s_93_29), .d(s_93_28), .cin(t_1657), .o(t_1690), .co(t_1691), .cout(t_1692));
compressor_4_2 u2_585(.a(s_93_35), .b(s_93_34), .c(s_93_33), .d(s_93_32), .cin(t_1660), .o(t_1693), .co(t_1694), .cout(t_1695));
compressor_4_2 u2_586(.a(s_93_39), .b(s_93_38), .c(s_93_37), .d(s_93_36), .cin(t_1663), .o(t_1696), .co(t_1697), .cout(t_1698));
compressor_4_2 u2_587(.a(s_93_43), .b(s_93_42), .c(s_93_41), .d(s_93_40), .cin(t_1666), .o(t_1699), .co(t_1700), .cout(t_1701));
compressor_3_2 u1_588(.a(s_93_46), .b(s_93_45), .cin(s_93_44), .o(t_1702), .cout(t_1703));
compressor_4_2 u2_589(.a(s_94_3), .b(s_94_2), .c(s_94_1), .d(s_94_0), .cin(t_1671), .o(t_1704), .co(t_1705), .cout(t_1706));
compressor_4_2 u2_590(.a(s_94_7), .b(s_94_6), .c(s_94_5), .d(s_94_4), .cin(t_1674), .o(t_1707), .co(t_1708), .cout(t_1709));
compressor_4_2 u2_591(.a(s_94_11), .b(s_94_10), .c(s_94_9), .d(s_94_8), .cin(t_1677), .o(t_1710), .co(t_1711), .cout(t_1712));
compressor_4_2 u2_592(.a(s_94_15), .b(s_94_14), .c(s_94_13), .d(s_94_12), .cin(t_1680), .o(t_1713), .co(t_1714), .cout(t_1715));
compressor_4_2 u2_593(.a(s_94_19), .b(s_94_18), .c(s_94_17), .d(s_94_16), .cin(t_1683), .o(t_1716), .co(t_1717), .cout(t_1718));
compressor_4_2 u2_594(.a(s_94_23), .b(s_94_22), .c(s_94_21), .d(s_94_20), .cin(t_1686), .o(t_1719), .co(t_1720), .cout(t_1721));
compressor_4_2 u2_595(.a(s_94_27), .b(s_94_26), .c(s_94_25), .d(s_94_24), .cin(t_1689), .o(t_1722), .co(t_1723), .cout(t_1724));
compressor_4_2 u2_596(.a(s_94_31), .b(s_94_30), .c(s_94_29), .d(s_94_28), .cin(t_1692), .o(t_1725), .co(t_1726), .cout(t_1727));
compressor_4_2 u2_597(.a(s_94_35), .b(s_94_34), .c(s_94_33), .d(s_94_32), .cin(t_1695), .o(t_1728), .co(t_1729), .cout(t_1730));
compressor_4_2 u2_598(.a(s_94_39), .b(s_94_38), .c(s_94_37), .d(s_94_36), .cin(t_1698), .o(t_1731), .co(t_1732), .cout(t_1733));
compressor_4_2 u2_599(.a(s_94_43), .b(s_94_42), .c(s_94_41), .d(s_94_40), .cin(t_1701), .o(t_1734), .co(t_1735), .cout(t_1736));
compressor_4_2 u2_600(.a(s_94_48), .b(s_94_47), .c(s_94_46), .d(s_94_45), .cin(s_94_44), .o(t_1737), .co(t_1738), .cout(t_1739));
compressor_4_2 u2_601(.a(s_95_3), .b(s_95_2), .c(s_95_1), .d(s_95_0), .cin(t_1706), .o(t_1740), .co(t_1741), .cout(t_1742));
compressor_4_2 u2_602(.a(s_95_7), .b(s_95_6), .c(s_95_5), .d(s_95_4), .cin(t_1709), .o(t_1743), .co(t_1744), .cout(t_1745));
compressor_4_2 u2_603(.a(s_95_11), .b(s_95_10), .c(s_95_9), .d(s_95_8), .cin(t_1712), .o(t_1746), .co(t_1747), .cout(t_1748));
compressor_4_2 u2_604(.a(s_95_15), .b(s_95_14), .c(s_95_13), .d(s_95_12), .cin(t_1715), .o(t_1749), .co(t_1750), .cout(t_1751));
compressor_4_2 u2_605(.a(s_95_19), .b(s_95_18), .c(s_95_17), .d(s_95_16), .cin(t_1718), .o(t_1752), .co(t_1753), .cout(t_1754));
compressor_4_2 u2_606(.a(s_95_23), .b(s_95_22), .c(s_95_21), .d(s_95_20), .cin(t_1721), .o(t_1755), .co(t_1756), .cout(t_1757));
compressor_4_2 u2_607(.a(s_95_27), .b(s_95_26), .c(s_95_25), .d(s_95_24), .cin(t_1724), .o(t_1758), .co(t_1759), .cout(t_1760));
compressor_4_2 u2_608(.a(s_95_31), .b(s_95_30), .c(s_95_29), .d(s_95_28), .cin(t_1727), .o(t_1761), .co(t_1762), .cout(t_1763));
compressor_4_2 u2_609(.a(s_95_35), .b(s_95_34), .c(s_95_33), .d(s_95_32), .cin(t_1730), .o(t_1764), .co(t_1765), .cout(t_1766));
compressor_4_2 u2_610(.a(s_95_39), .b(s_95_38), .c(s_95_37), .d(s_95_36), .cin(t_1733), .o(t_1767), .co(t_1768), .cout(t_1769));
compressor_4_2 u2_611(.a(s_95_43), .b(s_95_42), .c(s_95_41), .d(s_95_40), .cin(t_1736), .o(t_1770), .co(t_1771), .cout(t_1772));
compressor_4_2 u2_612(.a(s_95_47), .b(s_95_46), .c(s_95_45), .d(s_95_44), .cin(t_1739), .o(t_1773), .co(t_1774), .cout(t_1775));
compressor_4_2 u2_613(.a(s_96_3), .b(s_96_2), .c(s_96_1), .d(s_96_0), .cin(t_1742), .o(t_1776), .co(t_1777), .cout(t_1778));
compressor_4_2 u2_614(.a(s_96_7), .b(s_96_6), .c(s_96_5), .d(s_96_4), .cin(t_1745), .o(t_1779), .co(t_1780), .cout(t_1781));
compressor_4_2 u2_615(.a(s_96_11), .b(s_96_10), .c(s_96_9), .d(s_96_8), .cin(t_1748), .o(t_1782), .co(t_1783), .cout(t_1784));
compressor_4_2 u2_616(.a(s_96_15), .b(s_96_14), .c(s_96_13), .d(s_96_12), .cin(t_1751), .o(t_1785), .co(t_1786), .cout(t_1787));
compressor_4_2 u2_617(.a(s_96_19), .b(s_96_18), .c(s_96_17), .d(s_96_16), .cin(t_1754), .o(t_1788), .co(t_1789), .cout(t_1790));
compressor_4_2 u2_618(.a(s_96_23), .b(s_96_22), .c(s_96_21), .d(s_96_20), .cin(t_1757), .o(t_1791), .co(t_1792), .cout(t_1793));
compressor_4_2 u2_619(.a(s_96_27), .b(s_96_26), .c(s_96_25), .d(s_96_24), .cin(t_1760), .o(t_1794), .co(t_1795), .cout(t_1796));
compressor_4_2 u2_620(.a(s_96_31), .b(s_96_30), .c(s_96_29), .d(s_96_28), .cin(t_1763), .o(t_1797), .co(t_1798), .cout(t_1799));
compressor_4_2 u2_621(.a(s_96_35), .b(s_96_34), .c(s_96_33), .d(s_96_32), .cin(t_1766), .o(t_1800), .co(t_1801), .cout(t_1802));
compressor_4_2 u2_622(.a(s_96_39), .b(s_96_38), .c(s_96_37), .d(s_96_36), .cin(t_1769), .o(t_1803), .co(t_1804), .cout(t_1805));
compressor_4_2 u2_623(.a(s_96_43), .b(s_96_42), .c(s_96_41), .d(s_96_40), .cin(t_1772), .o(t_1806), .co(t_1807), .cout(t_1808));
compressor_4_2 u2_624(.a(s_96_47), .b(s_96_46), .c(s_96_45), .d(s_96_44), .cin(t_1775), .o(t_1809), .co(t_1810), .cout(t_1811));
half_adder u0_625(.a(s_96_49), .b(s_96_48), .o(t_1812), .cout(t_1813));
compressor_4_2 u2_626(.a(s_97_3), .b(s_97_2), .c(s_97_1), .d(s_97_0), .cin(t_1778), .o(t_1814), .co(t_1815), .cout(t_1816));
compressor_4_2 u2_627(.a(s_97_7), .b(s_97_6), .c(s_97_5), .d(s_97_4), .cin(t_1781), .o(t_1817), .co(t_1818), .cout(t_1819));
compressor_4_2 u2_628(.a(s_97_11), .b(s_97_10), .c(s_97_9), .d(s_97_8), .cin(t_1784), .o(t_1820), .co(t_1821), .cout(t_1822));
compressor_4_2 u2_629(.a(s_97_15), .b(s_97_14), .c(s_97_13), .d(s_97_12), .cin(t_1787), .o(t_1823), .co(t_1824), .cout(t_1825));
compressor_4_2 u2_630(.a(s_97_19), .b(s_97_18), .c(s_97_17), .d(s_97_16), .cin(t_1790), .o(t_1826), .co(t_1827), .cout(t_1828));
compressor_4_2 u2_631(.a(s_97_23), .b(s_97_22), .c(s_97_21), .d(s_97_20), .cin(t_1793), .o(t_1829), .co(t_1830), .cout(t_1831));
compressor_4_2 u2_632(.a(s_97_27), .b(s_97_26), .c(s_97_25), .d(s_97_24), .cin(t_1796), .o(t_1832), .co(t_1833), .cout(t_1834));
compressor_4_2 u2_633(.a(s_97_31), .b(s_97_30), .c(s_97_29), .d(s_97_28), .cin(t_1799), .o(t_1835), .co(t_1836), .cout(t_1837));
compressor_4_2 u2_634(.a(s_97_35), .b(s_97_34), .c(s_97_33), .d(s_97_32), .cin(t_1802), .o(t_1838), .co(t_1839), .cout(t_1840));
compressor_4_2 u2_635(.a(s_97_39), .b(s_97_38), .c(s_97_37), .d(s_97_36), .cin(t_1805), .o(t_1841), .co(t_1842), .cout(t_1843));
compressor_4_2 u2_636(.a(s_97_43), .b(s_97_42), .c(s_97_41), .d(s_97_40), .cin(t_1808), .o(t_1844), .co(t_1845), .cout(t_1846));
compressor_4_2 u2_637(.a(s_97_47), .b(s_97_46), .c(s_97_45), .d(s_97_44), .cin(t_1811), .o(t_1847), .co(t_1848), .cout(t_1849));
compressor_4_2 u2_638(.a(s_98_3), .b(s_98_2), .c(s_98_1), .d(s_98_0), .cin(t_1816), .o(t_1850), .co(t_1851), .cout(t_1852));
compressor_4_2 u2_639(.a(s_98_7), .b(s_98_6), .c(s_98_5), .d(s_98_4), .cin(t_1819), .o(t_1853), .co(t_1854), .cout(t_1855));
compressor_4_2 u2_640(.a(s_98_11), .b(s_98_10), .c(s_98_9), .d(s_98_8), .cin(t_1822), .o(t_1856), .co(t_1857), .cout(t_1858));
compressor_4_2 u2_641(.a(s_98_15), .b(s_98_14), .c(s_98_13), .d(s_98_12), .cin(t_1825), .o(t_1859), .co(t_1860), .cout(t_1861));
compressor_4_2 u2_642(.a(s_98_19), .b(s_98_18), .c(s_98_17), .d(s_98_16), .cin(t_1828), .o(t_1862), .co(t_1863), .cout(t_1864));
compressor_4_2 u2_643(.a(s_98_23), .b(s_98_22), .c(s_98_21), .d(s_98_20), .cin(t_1831), .o(t_1865), .co(t_1866), .cout(t_1867));
compressor_4_2 u2_644(.a(s_98_27), .b(s_98_26), .c(s_98_25), .d(s_98_24), .cin(t_1834), .o(t_1868), .co(t_1869), .cout(t_1870));
compressor_4_2 u2_645(.a(s_98_31), .b(s_98_30), .c(s_98_29), .d(s_98_28), .cin(t_1837), .o(t_1871), .co(t_1872), .cout(t_1873));
compressor_4_2 u2_646(.a(s_98_35), .b(s_98_34), .c(s_98_33), .d(s_98_32), .cin(t_1840), .o(t_1874), .co(t_1875), .cout(t_1876));
compressor_4_2 u2_647(.a(s_98_39), .b(s_98_38), .c(s_98_37), .d(s_98_36), .cin(t_1843), .o(t_1877), .co(t_1878), .cout(t_1879));
compressor_4_2 u2_648(.a(s_98_43), .b(s_98_42), .c(s_98_41), .d(s_98_40), .cin(t_1846), .o(t_1880), .co(t_1881), .cout(t_1882));
compressor_4_2 u2_649(.a(s_98_47), .b(s_98_46), .c(s_98_45), .d(s_98_44), .cin(t_1849), .o(t_1883), .co(t_1884), .cout(t_1885));
compressor_3_2 u1_650(.a(s_98_50), .b(s_98_49), .cin(s_98_48), .o(t_1886), .cout(t_1887));
compressor_4_2 u2_651(.a(s_99_3), .b(s_99_2), .c(s_99_1), .d(s_99_0), .cin(t_1852), .o(t_1888), .co(t_1889), .cout(t_1890));
compressor_4_2 u2_652(.a(s_99_7), .b(s_99_6), .c(s_99_5), .d(s_99_4), .cin(t_1855), .o(t_1891), .co(t_1892), .cout(t_1893));
compressor_4_2 u2_653(.a(s_99_11), .b(s_99_10), .c(s_99_9), .d(s_99_8), .cin(t_1858), .o(t_1894), .co(t_1895), .cout(t_1896));
compressor_4_2 u2_654(.a(s_99_15), .b(s_99_14), .c(s_99_13), .d(s_99_12), .cin(t_1861), .o(t_1897), .co(t_1898), .cout(t_1899));
compressor_4_2 u2_655(.a(s_99_19), .b(s_99_18), .c(s_99_17), .d(s_99_16), .cin(t_1864), .o(t_1900), .co(t_1901), .cout(t_1902));
compressor_4_2 u2_656(.a(s_99_23), .b(s_99_22), .c(s_99_21), .d(s_99_20), .cin(t_1867), .o(t_1903), .co(t_1904), .cout(t_1905));
compressor_4_2 u2_657(.a(s_99_27), .b(s_99_26), .c(s_99_25), .d(s_99_24), .cin(t_1870), .o(t_1906), .co(t_1907), .cout(t_1908));
compressor_4_2 u2_658(.a(s_99_31), .b(s_99_30), .c(s_99_29), .d(s_99_28), .cin(t_1873), .o(t_1909), .co(t_1910), .cout(t_1911));
compressor_4_2 u2_659(.a(s_99_35), .b(s_99_34), .c(s_99_33), .d(s_99_32), .cin(t_1876), .o(t_1912), .co(t_1913), .cout(t_1914));
compressor_4_2 u2_660(.a(s_99_39), .b(s_99_38), .c(s_99_37), .d(s_99_36), .cin(t_1879), .o(t_1915), .co(t_1916), .cout(t_1917));
compressor_4_2 u2_661(.a(s_99_43), .b(s_99_42), .c(s_99_41), .d(s_99_40), .cin(t_1882), .o(t_1918), .co(t_1919), .cout(t_1920));
compressor_4_2 u2_662(.a(s_99_47), .b(s_99_46), .c(s_99_45), .d(s_99_44), .cin(t_1885), .o(t_1921), .co(t_1922), .cout(t_1923));
half_adder u0_663(.a(s_99_49), .b(s_99_48), .o(t_1924), .cout(t_1925));
compressor_4_2 u2_664(.a(s_100_3), .b(s_100_2), .c(s_100_1), .d(s_100_0), .cin(t_1890), .o(t_1926), .co(t_1927), .cout(t_1928));
compressor_4_2 u2_665(.a(s_100_7), .b(s_100_6), .c(s_100_5), .d(s_100_4), .cin(t_1893), .o(t_1929), .co(t_1930), .cout(t_1931));
compressor_4_2 u2_666(.a(s_100_11), .b(s_100_10), .c(s_100_9), .d(s_100_8), .cin(t_1896), .o(t_1932), .co(t_1933), .cout(t_1934));
compressor_4_2 u2_667(.a(s_100_15), .b(s_100_14), .c(s_100_13), .d(s_100_12), .cin(t_1899), .o(t_1935), .co(t_1936), .cout(t_1937));
compressor_4_2 u2_668(.a(s_100_19), .b(s_100_18), .c(s_100_17), .d(s_100_16), .cin(t_1902), .o(t_1938), .co(t_1939), .cout(t_1940));
compressor_4_2 u2_669(.a(s_100_23), .b(s_100_22), .c(s_100_21), .d(s_100_20), .cin(t_1905), .o(t_1941), .co(t_1942), .cout(t_1943));
compressor_4_2 u2_670(.a(s_100_27), .b(s_100_26), .c(s_100_25), .d(s_100_24), .cin(t_1908), .o(t_1944), .co(t_1945), .cout(t_1946));
compressor_4_2 u2_671(.a(s_100_31), .b(s_100_30), .c(s_100_29), .d(s_100_28), .cin(t_1911), .o(t_1947), .co(t_1948), .cout(t_1949));
compressor_4_2 u2_672(.a(s_100_35), .b(s_100_34), .c(s_100_33), .d(s_100_32), .cin(t_1914), .o(t_1950), .co(t_1951), .cout(t_1952));
compressor_4_2 u2_673(.a(s_100_39), .b(s_100_38), .c(s_100_37), .d(s_100_36), .cin(t_1917), .o(t_1953), .co(t_1954), .cout(t_1955));
compressor_4_2 u2_674(.a(s_100_43), .b(s_100_42), .c(s_100_41), .d(s_100_40), .cin(t_1920), .o(t_1956), .co(t_1957), .cout(t_1958));
compressor_4_2 u2_675(.a(s_100_47), .b(s_100_46), .c(s_100_45), .d(s_100_44), .cin(t_1923), .o(t_1959), .co(t_1960), .cout(t_1961));
compressor_3_2 u1_676(.a(s_100_50), .b(s_100_49), .cin(s_100_48), .o(t_1962), .cout(t_1963));
compressor_4_2 u2_677(.a(s_101_3), .b(s_101_2), .c(s_101_1), .d(s_101_0), .cin(t_1928), .o(t_1964), .co(t_1965), .cout(t_1966));
compressor_4_2 u2_678(.a(s_101_7), .b(s_101_6), .c(s_101_5), .d(s_101_4), .cin(t_1931), .o(t_1967), .co(t_1968), .cout(t_1969));
compressor_4_2 u2_679(.a(s_101_11), .b(s_101_10), .c(s_101_9), .d(s_101_8), .cin(t_1934), .o(t_1970), .co(t_1971), .cout(t_1972));
compressor_4_2 u2_680(.a(s_101_15), .b(s_101_14), .c(s_101_13), .d(s_101_12), .cin(t_1937), .o(t_1973), .co(t_1974), .cout(t_1975));
compressor_4_2 u2_681(.a(s_101_19), .b(s_101_18), .c(s_101_17), .d(s_101_16), .cin(t_1940), .o(t_1976), .co(t_1977), .cout(t_1978));
compressor_4_2 u2_682(.a(s_101_23), .b(s_101_22), .c(s_101_21), .d(s_101_20), .cin(t_1943), .o(t_1979), .co(t_1980), .cout(t_1981));
compressor_4_2 u2_683(.a(s_101_27), .b(s_101_26), .c(s_101_25), .d(s_101_24), .cin(t_1946), .o(t_1982), .co(t_1983), .cout(t_1984));
compressor_4_2 u2_684(.a(s_101_31), .b(s_101_30), .c(s_101_29), .d(s_101_28), .cin(t_1949), .o(t_1985), .co(t_1986), .cout(t_1987));
compressor_4_2 u2_685(.a(s_101_35), .b(s_101_34), .c(s_101_33), .d(s_101_32), .cin(t_1952), .o(t_1988), .co(t_1989), .cout(t_1990));
compressor_4_2 u2_686(.a(s_101_39), .b(s_101_38), .c(s_101_37), .d(s_101_36), .cin(t_1955), .o(t_1991), .co(t_1992), .cout(t_1993));
compressor_4_2 u2_687(.a(s_101_43), .b(s_101_42), .c(s_101_41), .d(s_101_40), .cin(t_1958), .o(t_1994), .co(t_1995), .cout(t_1996));
compressor_4_2 u2_688(.a(s_101_47), .b(s_101_46), .c(s_101_45), .d(s_101_44), .cin(t_1961), .o(t_1997), .co(t_1998), .cout(t_1999));
compressor_3_2 u1_689(.a(s_101_50), .b(s_101_49), .cin(s_101_48), .o(t_2000), .cout(t_2001));
compressor_4_2 u2_690(.a(s_102_3), .b(s_102_2), .c(s_102_1), .d(s_102_0), .cin(t_1966), .o(t_2002), .co(t_2003), .cout(t_2004));
compressor_4_2 u2_691(.a(s_102_7), .b(s_102_6), .c(s_102_5), .d(s_102_4), .cin(t_1969), .o(t_2005), .co(t_2006), .cout(t_2007));
compressor_4_2 u2_692(.a(s_102_11), .b(s_102_10), .c(s_102_9), .d(s_102_8), .cin(t_1972), .o(t_2008), .co(t_2009), .cout(t_2010));
compressor_4_2 u2_693(.a(s_102_15), .b(s_102_14), .c(s_102_13), .d(s_102_12), .cin(t_1975), .o(t_2011), .co(t_2012), .cout(t_2013));
compressor_4_2 u2_694(.a(s_102_19), .b(s_102_18), .c(s_102_17), .d(s_102_16), .cin(t_1978), .o(t_2014), .co(t_2015), .cout(t_2016));
compressor_4_2 u2_695(.a(s_102_23), .b(s_102_22), .c(s_102_21), .d(s_102_20), .cin(t_1981), .o(t_2017), .co(t_2018), .cout(t_2019));
compressor_4_2 u2_696(.a(s_102_27), .b(s_102_26), .c(s_102_25), .d(s_102_24), .cin(t_1984), .o(t_2020), .co(t_2021), .cout(t_2022));
compressor_4_2 u2_697(.a(s_102_31), .b(s_102_30), .c(s_102_29), .d(s_102_28), .cin(t_1987), .o(t_2023), .co(t_2024), .cout(t_2025));
compressor_4_2 u2_698(.a(s_102_35), .b(s_102_34), .c(s_102_33), .d(s_102_32), .cin(t_1990), .o(t_2026), .co(t_2027), .cout(t_2028));
compressor_4_2 u2_699(.a(s_102_39), .b(s_102_38), .c(s_102_37), .d(s_102_36), .cin(t_1993), .o(t_2029), .co(t_2030), .cout(t_2031));
compressor_4_2 u2_700(.a(s_102_43), .b(s_102_42), .c(s_102_41), .d(s_102_40), .cin(t_1996), .o(t_2032), .co(t_2033), .cout(t_2034));
compressor_4_2 u2_701(.a(s_102_47), .b(s_102_46), .c(s_102_45), .d(s_102_44), .cin(t_1999), .o(t_2035), .co(t_2036), .cout(t_2037));
compressor_4_2 u2_702(.a(s_102_52), .b(s_102_51), .c(s_102_50), .d(s_102_49), .cin(s_102_48), .o(t_2038), .co(t_2039), .cout(t_2040));
compressor_4_2 u2_703(.a(s_103_3), .b(s_103_2), .c(s_103_1), .d(s_103_0), .cin(t_2004), .o(t_2041), .co(t_2042), .cout(t_2043));
compressor_4_2 u2_704(.a(s_103_7), .b(s_103_6), .c(s_103_5), .d(s_103_4), .cin(t_2007), .o(t_2044), .co(t_2045), .cout(t_2046));
compressor_4_2 u2_705(.a(s_103_11), .b(s_103_10), .c(s_103_9), .d(s_103_8), .cin(t_2010), .o(t_2047), .co(t_2048), .cout(t_2049));
compressor_4_2 u2_706(.a(s_103_15), .b(s_103_14), .c(s_103_13), .d(s_103_12), .cin(t_2013), .o(t_2050), .co(t_2051), .cout(t_2052));
compressor_4_2 u2_707(.a(s_103_19), .b(s_103_18), .c(s_103_17), .d(s_103_16), .cin(t_2016), .o(t_2053), .co(t_2054), .cout(t_2055));
compressor_4_2 u2_708(.a(s_103_23), .b(s_103_22), .c(s_103_21), .d(s_103_20), .cin(t_2019), .o(t_2056), .co(t_2057), .cout(t_2058));
compressor_4_2 u2_709(.a(s_103_27), .b(s_103_26), .c(s_103_25), .d(s_103_24), .cin(t_2022), .o(t_2059), .co(t_2060), .cout(t_2061));
compressor_4_2 u2_710(.a(s_103_31), .b(s_103_30), .c(s_103_29), .d(s_103_28), .cin(t_2025), .o(t_2062), .co(t_2063), .cout(t_2064));
compressor_4_2 u2_711(.a(s_103_35), .b(s_103_34), .c(s_103_33), .d(s_103_32), .cin(t_2028), .o(t_2065), .co(t_2066), .cout(t_2067));
compressor_4_2 u2_712(.a(s_103_39), .b(s_103_38), .c(s_103_37), .d(s_103_36), .cin(t_2031), .o(t_2068), .co(t_2069), .cout(t_2070));
compressor_4_2 u2_713(.a(s_103_43), .b(s_103_42), .c(s_103_41), .d(s_103_40), .cin(t_2034), .o(t_2071), .co(t_2072), .cout(t_2073));
compressor_4_2 u2_714(.a(s_103_47), .b(s_103_46), .c(s_103_45), .d(s_103_44), .cin(t_2037), .o(t_2074), .co(t_2075), .cout(t_2076));
compressor_4_2 u2_715(.a(s_103_51), .b(s_103_50), .c(s_103_49), .d(s_103_48), .cin(t_2040), .o(t_2077), .co(t_2078), .cout(t_2079));
compressor_4_2 u2_716(.a(s_104_3), .b(s_104_2), .c(s_104_1), .d(s_104_0), .cin(t_2043), .o(t_2080), .co(t_2081), .cout(t_2082));
compressor_4_2 u2_717(.a(s_104_7), .b(s_104_6), .c(s_104_5), .d(s_104_4), .cin(t_2046), .o(t_2083), .co(t_2084), .cout(t_2085));
compressor_4_2 u2_718(.a(s_104_11), .b(s_104_10), .c(s_104_9), .d(s_104_8), .cin(t_2049), .o(t_2086), .co(t_2087), .cout(t_2088));
compressor_4_2 u2_719(.a(s_104_15), .b(s_104_14), .c(s_104_13), .d(s_104_12), .cin(t_2052), .o(t_2089), .co(t_2090), .cout(t_2091));
compressor_4_2 u2_720(.a(s_104_19), .b(s_104_18), .c(s_104_17), .d(s_104_16), .cin(t_2055), .o(t_2092), .co(t_2093), .cout(t_2094));
compressor_4_2 u2_721(.a(s_104_23), .b(s_104_22), .c(s_104_21), .d(s_104_20), .cin(t_2058), .o(t_2095), .co(t_2096), .cout(t_2097));
compressor_4_2 u2_722(.a(s_104_27), .b(s_104_26), .c(s_104_25), .d(s_104_24), .cin(t_2061), .o(t_2098), .co(t_2099), .cout(t_2100));
compressor_4_2 u2_723(.a(s_104_31), .b(s_104_30), .c(s_104_29), .d(s_104_28), .cin(t_2064), .o(t_2101), .co(t_2102), .cout(t_2103));
compressor_4_2 u2_724(.a(s_104_35), .b(s_104_34), .c(s_104_33), .d(s_104_32), .cin(t_2067), .o(t_2104), .co(t_2105), .cout(t_2106));
compressor_4_2 u2_725(.a(s_104_39), .b(s_104_38), .c(s_104_37), .d(s_104_36), .cin(t_2070), .o(t_2107), .co(t_2108), .cout(t_2109));
compressor_4_2 u2_726(.a(s_104_43), .b(s_104_42), .c(s_104_41), .d(s_104_40), .cin(t_2073), .o(t_2110), .co(t_2111), .cout(t_2112));
compressor_4_2 u2_727(.a(s_104_47), .b(s_104_46), .c(s_104_45), .d(s_104_44), .cin(t_2076), .o(t_2113), .co(t_2114), .cout(t_2115));
compressor_4_2 u2_728(.a(s_104_51), .b(s_104_50), .c(s_104_49), .d(s_104_48), .cin(t_2079), .o(t_2116), .co(t_2117), .cout(t_2118));
half_adder u0_729(.a(s_104_53), .b(s_104_52), .o(t_2119), .cout(t_2120));
compressor_4_2 u2_730(.a(s_105_3), .b(s_105_2), .c(s_105_1), .d(s_105_0), .cin(t_2082), .o(t_2121), .co(t_2122), .cout(t_2123));
compressor_4_2 u2_731(.a(s_105_7), .b(s_105_6), .c(s_105_5), .d(s_105_4), .cin(t_2085), .o(t_2124), .co(t_2125), .cout(t_2126));
compressor_4_2 u2_732(.a(s_105_11), .b(s_105_10), .c(s_105_9), .d(s_105_8), .cin(t_2088), .o(t_2127), .co(t_2128), .cout(t_2129));
compressor_4_2 u2_733(.a(s_105_15), .b(s_105_14), .c(s_105_13), .d(s_105_12), .cin(t_2091), .o(t_2130), .co(t_2131), .cout(t_2132));
compressor_4_2 u2_734(.a(s_105_19), .b(s_105_18), .c(s_105_17), .d(s_105_16), .cin(t_2094), .o(t_2133), .co(t_2134), .cout(t_2135));
compressor_4_2 u2_735(.a(s_105_23), .b(s_105_22), .c(s_105_21), .d(s_105_20), .cin(t_2097), .o(t_2136), .co(t_2137), .cout(t_2138));
compressor_4_2 u2_736(.a(s_105_27), .b(s_105_26), .c(s_105_25), .d(s_105_24), .cin(t_2100), .o(t_2139), .co(t_2140), .cout(t_2141));
compressor_4_2 u2_737(.a(s_105_31), .b(s_105_30), .c(s_105_29), .d(s_105_28), .cin(t_2103), .o(t_2142), .co(t_2143), .cout(t_2144));
compressor_4_2 u2_738(.a(s_105_35), .b(s_105_34), .c(s_105_33), .d(s_105_32), .cin(t_2106), .o(t_2145), .co(t_2146), .cout(t_2147));
compressor_4_2 u2_739(.a(s_105_39), .b(s_105_38), .c(s_105_37), .d(s_105_36), .cin(t_2109), .o(t_2148), .co(t_2149), .cout(t_2150));
compressor_4_2 u2_740(.a(s_105_43), .b(s_105_42), .c(s_105_41), .d(s_105_40), .cin(t_2112), .o(t_2151), .co(t_2152), .cout(t_2153));
compressor_4_2 u2_741(.a(s_105_47), .b(s_105_46), .c(s_105_45), .d(s_105_44), .cin(t_2115), .o(t_2154), .co(t_2155), .cout(t_2156));
compressor_4_2 u2_742(.a(s_105_51), .b(s_105_50), .c(s_105_49), .d(s_105_48), .cin(t_2118), .o(t_2157), .co(t_2158), .cout(t_2159));
compressor_4_2 u2_743(.a(s_106_3), .b(s_106_2), .c(s_106_1), .d(s_106_0), .cin(t_2123), .o(t_2160), .co(t_2161), .cout(t_2162));
compressor_4_2 u2_744(.a(s_106_7), .b(s_106_6), .c(s_106_5), .d(s_106_4), .cin(t_2126), .o(t_2163), .co(t_2164), .cout(t_2165));
compressor_4_2 u2_745(.a(s_106_11), .b(s_106_10), .c(s_106_9), .d(s_106_8), .cin(t_2129), .o(t_2166), .co(t_2167), .cout(t_2168));
compressor_4_2 u2_746(.a(s_106_15), .b(s_106_14), .c(s_106_13), .d(s_106_12), .cin(t_2132), .o(t_2169), .co(t_2170), .cout(t_2171));
compressor_4_2 u2_747(.a(s_106_19), .b(s_106_18), .c(s_106_17), .d(s_106_16), .cin(t_2135), .o(t_2172), .co(t_2173), .cout(t_2174));
compressor_4_2 u2_748(.a(s_106_23), .b(s_106_22), .c(s_106_21), .d(s_106_20), .cin(t_2138), .o(t_2175), .co(t_2176), .cout(t_2177));
compressor_4_2 u2_749(.a(s_106_27), .b(s_106_26), .c(s_106_25), .d(s_106_24), .cin(t_2141), .o(t_2178), .co(t_2179), .cout(t_2180));
compressor_4_2 u2_750(.a(s_106_31), .b(s_106_30), .c(s_106_29), .d(s_106_28), .cin(t_2144), .o(t_2181), .co(t_2182), .cout(t_2183));
compressor_4_2 u2_751(.a(s_106_35), .b(s_106_34), .c(s_106_33), .d(s_106_32), .cin(t_2147), .o(t_2184), .co(t_2185), .cout(t_2186));
compressor_4_2 u2_752(.a(s_106_39), .b(s_106_38), .c(s_106_37), .d(s_106_36), .cin(t_2150), .o(t_2187), .co(t_2188), .cout(t_2189));
compressor_4_2 u2_753(.a(s_106_43), .b(s_106_42), .c(s_106_41), .d(s_106_40), .cin(t_2153), .o(t_2190), .co(t_2191), .cout(t_2192));
compressor_4_2 u2_754(.a(s_106_47), .b(s_106_46), .c(s_106_45), .d(s_106_44), .cin(t_2156), .o(t_2193), .co(t_2194), .cout(t_2195));
compressor_4_2 u2_755(.a(s_106_51), .b(s_106_50), .c(s_106_49), .d(s_106_48), .cin(t_2159), .o(t_2196), .co(t_2197), .cout(t_2198));
compressor_3_2 u1_756(.a(s_106_54), .b(s_106_53), .cin(s_106_52), .o(t_2199), .cout(t_2200));
compressor_4_2 u2_757(.a(s_107_3), .b(s_107_2), .c(s_107_1), .d(s_107_0), .cin(t_2162), .o(t_2201), .co(t_2202), .cout(t_2203));
compressor_4_2 u2_758(.a(s_107_7), .b(s_107_6), .c(s_107_5), .d(s_107_4), .cin(t_2165), .o(t_2204), .co(t_2205), .cout(t_2206));
compressor_4_2 u2_759(.a(s_107_11), .b(s_107_10), .c(s_107_9), .d(s_107_8), .cin(t_2168), .o(t_2207), .co(t_2208), .cout(t_2209));
compressor_4_2 u2_760(.a(s_107_15), .b(s_107_14), .c(s_107_13), .d(s_107_12), .cin(t_2171), .o(t_2210), .co(t_2211), .cout(t_2212));
compressor_4_2 u2_761(.a(s_107_19), .b(s_107_18), .c(s_107_17), .d(s_107_16), .cin(t_2174), .o(t_2213), .co(t_2214), .cout(t_2215));
compressor_4_2 u2_762(.a(s_107_23), .b(s_107_22), .c(s_107_21), .d(s_107_20), .cin(t_2177), .o(t_2216), .co(t_2217), .cout(t_2218));
compressor_4_2 u2_763(.a(s_107_27), .b(s_107_26), .c(s_107_25), .d(s_107_24), .cin(t_2180), .o(t_2219), .co(t_2220), .cout(t_2221));
compressor_4_2 u2_764(.a(s_107_31), .b(s_107_30), .c(s_107_29), .d(s_107_28), .cin(t_2183), .o(t_2222), .co(t_2223), .cout(t_2224));
compressor_4_2 u2_765(.a(s_107_35), .b(s_107_34), .c(s_107_33), .d(s_107_32), .cin(t_2186), .o(t_2225), .co(t_2226), .cout(t_2227));
compressor_4_2 u2_766(.a(s_107_39), .b(s_107_38), .c(s_107_37), .d(s_107_36), .cin(t_2189), .o(t_2228), .co(t_2229), .cout(t_2230));
compressor_4_2 u2_767(.a(s_107_43), .b(s_107_42), .c(s_107_41), .d(s_107_40), .cin(t_2192), .o(t_2231), .co(t_2232), .cout(t_2233));
compressor_4_2 u2_768(.a(s_107_47), .b(s_107_46), .c(s_107_45), .d(s_107_44), .cin(t_2195), .o(t_2234), .co(t_2235), .cout(t_2236));
compressor_4_2 u2_769(.a(s_107_51), .b(s_107_50), .c(s_107_49), .d(s_107_48), .cin(t_2198), .o(t_2237), .co(t_2238), .cout(t_2239));
half_adder u0_770(.a(s_107_53), .b(s_107_52), .o(t_2240), .cout(t_2241));
compressor_4_2 u2_771(.a(s_108_3), .b(s_108_2), .c(s_108_1), .d(s_108_0), .cin(t_2203), .o(t_2242), .co(t_2243), .cout(t_2244));
compressor_4_2 u2_772(.a(s_108_7), .b(s_108_6), .c(s_108_5), .d(s_108_4), .cin(t_2206), .o(t_2245), .co(t_2246), .cout(t_2247));
compressor_4_2 u2_773(.a(s_108_11), .b(s_108_10), .c(s_108_9), .d(s_108_8), .cin(t_2209), .o(t_2248), .co(t_2249), .cout(t_2250));
compressor_4_2 u2_774(.a(s_108_15), .b(s_108_14), .c(s_108_13), .d(s_108_12), .cin(t_2212), .o(t_2251), .co(t_2252), .cout(t_2253));
compressor_4_2 u2_775(.a(s_108_19), .b(s_108_18), .c(s_108_17), .d(s_108_16), .cin(t_2215), .o(t_2254), .co(t_2255), .cout(t_2256));
compressor_4_2 u2_776(.a(s_108_23), .b(s_108_22), .c(s_108_21), .d(s_108_20), .cin(t_2218), .o(t_2257), .co(t_2258), .cout(t_2259));
compressor_4_2 u2_777(.a(s_108_27), .b(s_108_26), .c(s_108_25), .d(s_108_24), .cin(t_2221), .o(t_2260), .co(t_2261), .cout(t_2262));
compressor_4_2 u2_778(.a(s_108_31), .b(s_108_30), .c(s_108_29), .d(s_108_28), .cin(t_2224), .o(t_2263), .co(t_2264), .cout(t_2265));
compressor_4_2 u2_779(.a(s_108_35), .b(s_108_34), .c(s_108_33), .d(s_108_32), .cin(t_2227), .o(t_2266), .co(t_2267), .cout(t_2268));
compressor_4_2 u2_780(.a(s_108_39), .b(s_108_38), .c(s_108_37), .d(s_108_36), .cin(t_2230), .o(t_2269), .co(t_2270), .cout(t_2271));
compressor_4_2 u2_781(.a(s_108_43), .b(s_108_42), .c(s_108_41), .d(s_108_40), .cin(t_2233), .o(t_2272), .co(t_2273), .cout(t_2274));
compressor_4_2 u2_782(.a(s_108_47), .b(s_108_46), .c(s_108_45), .d(s_108_44), .cin(t_2236), .o(t_2275), .co(t_2276), .cout(t_2277));
compressor_4_2 u2_783(.a(s_108_51), .b(s_108_50), .c(s_108_49), .d(s_108_48), .cin(t_2239), .o(t_2278), .co(t_2279), .cout(t_2280));
compressor_3_2 u1_784(.a(s_108_54), .b(s_108_53), .cin(s_108_52), .o(t_2281), .cout(t_2282));
compressor_4_2 u2_785(.a(s_109_3), .b(s_109_2), .c(s_109_1), .d(s_109_0), .cin(t_2244), .o(t_2283), .co(t_2284), .cout(t_2285));
compressor_4_2 u2_786(.a(s_109_7), .b(s_109_6), .c(s_109_5), .d(s_109_4), .cin(t_2247), .o(t_2286), .co(t_2287), .cout(t_2288));
compressor_4_2 u2_787(.a(s_109_11), .b(s_109_10), .c(s_109_9), .d(s_109_8), .cin(t_2250), .o(t_2289), .co(t_2290), .cout(t_2291));
compressor_4_2 u2_788(.a(s_109_15), .b(s_109_14), .c(s_109_13), .d(s_109_12), .cin(t_2253), .o(t_2292), .co(t_2293), .cout(t_2294));
compressor_4_2 u2_789(.a(s_109_19), .b(s_109_18), .c(s_109_17), .d(s_109_16), .cin(t_2256), .o(t_2295), .co(t_2296), .cout(t_2297));
compressor_4_2 u2_790(.a(s_109_23), .b(s_109_22), .c(s_109_21), .d(s_109_20), .cin(t_2259), .o(t_2298), .co(t_2299), .cout(t_2300));
compressor_4_2 u2_791(.a(s_109_27), .b(s_109_26), .c(s_109_25), .d(s_109_24), .cin(t_2262), .o(t_2301), .co(t_2302), .cout(t_2303));
compressor_4_2 u2_792(.a(s_109_31), .b(s_109_30), .c(s_109_29), .d(s_109_28), .cin(t_2265), .o(t_2304), .co(t_2305), .cout(t_2306));
compressor_4_2 u2_793(.a(s_109_35), .b(s_109_34), .c(s_109_33), .d(s_109_32), .cin(t_2268), .o(t_2307), .co(t_2308), .cout(t_2309));
compressor_4_2 u2_794(.a(s_109_39), .b(s_109_38), .c(s_109_37), .d(s_109_36), .cin(t_2271), .o(t_2310), .co(t_2311), .cout(t_2312));
compressor_4_2 u2_795(.a(s_109_43), .b(s_109_42), .c(s_109_41), .d(s_109_40), .cin(t_2274), .o(t_2313), .co(t_2314), .cout(t_2315));
compressor_4_2 u2_796(.a(s_109_47), .b(s_109_46), .c(s_109_45), .d(s_109_44), .cin(t_2277), .o(t_2316), .co(t_2317), .cout(t_2318));
compressor_4_2 u2_797(.a(s_109_51), .b(s_109_50), .c(s_109_49), .d(s_109_48), .cin(t_2280), .o(t_2319), .co(t_2320), .cout(t_2321));
compressor_3_2 u1_798(.a(s_109_54), .b(s_109_53), .cin(s_109_52), .o(t_2322), .cout(t_2323));
compressor_4_2 u2_799(.a(s_110_3), .b(s_110_2), .c(s_110_1), .d(s_110_0), .cin(t_2285), .o(t_2324), .co(t_2325), .cout(t_2326));
compressor_4_2 u2_800(.a(s_110_7), .b(s_110_6), .c(s_110_5), .d(s_110_4), .cin(t_2288), .o(t_2327), .co(t_2328), .cout(t_2329));
compressor_4_2 u2_801(.a(s_110_11), .b(s_110_10), .c(s_110_9), .d(s_110_8), .cin(t_2291), .o(t_2330), .co(t_2331), .cout(t_2332));
compressor_4_2 u2_802(.a(s_110_15), .b(s_110_14), .c(s_110_13), .d(s_110_12), .cin(t_2294), .o(t_2333), .co(t_2334), .cout(t_2335));
compressor_4_2 u2_803(.a(s_110_19), .b(s_110_18), .c(s_110_17), .d(s_110_16), .cin(t_2297), .o(t_2336), .co(t_2337), .cout(t_2338));
compressor_4_2 u2_804(.a(s_110_23), .b(s_110_22), .c(s_110_21), .d(s_110_20), .cin(t_2300), .o(t_2339), .co(t_2340), .cout(t_2341));
compressor_4_2 u2_805(.a(s_110_27), .b(s_110_26), .c(s_110_25), .d(s_110_24), .cin(t_2303), .o(t_2342), .co(t_2343), .cout(t_2344));
compressor_4_2 u2_806(.a(s_110_31), .b(s_110_30), .c(s_110_29), .d(s_110_28), .cin(t_2306), .o(t_2345), .co(t_2346), .cout(t_2347));
compressor_4_2 u2_807(.a(s_110_35), .b(s_110_34), .c(s_110_33), .d(s_110_32), .cin(t_2309), .o(t_2348), .co(t_2349), .cout(t_2350));
compressor_4_2 u2_808(.a(s_110_39), .b(s_110_38), .c(s_110_37), .d(s_110_36), .cin(t_2312), .o(t_2351), .co(t_2352), .cout(t_2353));
compressor_4_2 u2_809(.a(s_110_43), .b(s_110_42), .c(s_110_41), .d(s_110_40), .cin(t_2315), .o(t_2354), .co(t_2355), .cout(t_2356));
compressor_4_2 u2_810(.a(s_110_47), .b(s_110_46), .c(s_110_45), .d(s_110_44), .cin(t_2318), .o(t_2357), .co(t_2358), .cout(t_2359));
compressor_4_2 u2_811(.a(s_110_51), .b(s_110_50), .c(s_110_49), .d(s_110_48), .cin(t_2321), .o(t_2360), .co(t_2361), .cout(t_2362));
compressor_4_2 u2_812(.a(s_110_56), .b(s_110_55), .c(s_110_54), .d(s_110_53), .cin(s_110_52), .o(t_2363), .co(t_2364), .cout(t_2365));
compressor_4_2 u2_813(.a(s_111_3), .b(s_111_2), .c(s_111_1), .d(s_111_0), .cin(t_2326), .o(t_2366), .co(t_2367), .cout(t_2368));
compressor_4_2 u2_814(.a(s_111_7), .b(s_111_6), .c(s_111_5), .d(s_111_4), .cin(t_2329), .o(t_2369), .co(t_2370), .cout(t_2371));
compressor_4_2 u2_815(.a(s_111_11), .b(s_111_10), .c(s_111_9), .d(s_111_8), .cin(t_2332), .o(t_2372), .co(t_2373), .cout(t_2374));
compressor_4_2 u2_816(.a(s_111_15), .b(s_111_14), .c(s_111_13), .d(s_111_12), .cin(t_2335), .o(t_2375), .co(t_2376), .cout(t_2377));
compressor_4_2 u2_817(.a(s_111_19), .b(s_111_18), .c(s_111_17), .d(s_111_16), .cin(t_2338), .o(t_2378), .co(t_2379), .cout(t_2380));
compressor_4_2 u2_818(.a(s_111_23), .b(s_111_22), .c(s_111_21), .d(s_111_20), .cin(t_2341), .o(t_2381), .co(t_2382), .cout(t_2383));
compressor_4_2 u2_819(.a(s_111_27), .b(s_111_26), .c(s_111_25), .d(s_111_24), .cin(t_2344), .o(t_2384), .co(t_2385), .cout(t_2386));
compressor_4_2 u2_820(.a(s_111_31), .b(s_111_30), .c(s_111_29), .d(s_111_28), .cin(t_2347), .o(t_2387), .co(t_2388), .cout(t_2389));
compressor_4_2 u2_821(.a(s_111_35), .b(s_111_34), .c(s_111_33), .d(s_111_32), .cin(t_2350), .o(t_2390), .co(t_2391), .cout(t_2392));
compressor_4_2 u2_822(.a(s_111_39), .b(s_111_38), .c(s_111_37), .d(s_111_36), .cin(t_2353), .o(t_2393), .co(t_2394), .cout(t_2395));
compressor_4_2 u2_823(.a(s_111_43), .b(s_111_42), .c(s_111_41), .d(s_111_40), .cin(t_2356), .o(t_2396), .co(t_2397), .cout(t_2398));
compressor_4_2 u2_824(.a(s_111_47), .b(s_111_46), .c(s_111_45), .d(s_111_44), .cin(t_2359), .o(t_2399), .co(t_2400), .cout(t_2401));
compressor_4_2 u2_825(.a(s_111_51), .b(s_111_50), .c(s_111_49), .d(s_111_48), .cin(t_2362), .o(t_2402), .co(t_2403), .cout(t_2404));
compressor_4_2 u2_826(.a(s_111_55), .b(s_111_54), .c(s_111_53), .d(s_111_52), .cin(t_2365), .o(t_2405), .co(t_2406), .cout(t_2407));
compressor_4_2 u2_827(.a(s_112_3), .b(s_112_2), .c(s_112_1), .d(s_112_0), .cin(t_2368), .o(t_2408), .co(t_2409), .cout(t_2410));
compressor_4_2 u2_828(.a(s_112_7), .b(s_112_6), .c(s_112_5), .d(s_112_4), .cin(t_2371), .o(t_2411), .co(t_2412), .cout(t_2413));
compressor_4_2 u2_829(.a(s_112_11), .b(s_112_10), .c(s_112_9), .d(s_112_8), .cin(t_2374), .o(t_2414), .co(t_2415), .cout(t_2416));
compressor_4_2 u2_830(.a(s_112_15), .b(s_112_14), .c(s_112_13), .d(s_112_12), .cin(t_2377), .o(t_2417), .co(t_2418), .cout(t_2419));
compressor_4_2 u2_831(.a(s_112_19), .b(s_112_18), .c(s_112_17), .d(s_112_16), .cin(t_2380), .o(t_2420), .co(t_2421), .cout(t_2422));
compressor_4_2 u2_832(.a(s_112_23), .b(s_112_22), .c(s_112_21), .d(s_112_20), .cin(t_2383), .o(t_2423), .co(t_2424), .cout(t_2425));
compressor_4_2 u2_833(.a(s_112_27), .b(s_112_26), .c(s_112_25), .d(s_112_24), .cin(t_2386), .o(t_2426), .co(t_2427), .cout(t_2428));
compressor_4_2 u2_834(.a(s_112_31), .b(s_112_30), .c(s_112_29), .d(s_112_28), .cin(t_2389), .o(t_2429), .co(t_2430), .cout(t_2431));
compressor_4_2 u2_835(.a(s_112_35), .b(s_112_34), .c(s_112_33), .d(s_112_32), .cin(t_2392), .o(t_2432), .co(t_2433), .cout(t_2434));
compressor_4_2 u2_836(.a(s_112_39), .b(s_112_38), .c(s_112_37), .d(s_112_36), .cin(t_2395), .o(t_2435), .co(t_2436), .cout(t_2437));
compressor_4_2 u2_837(.a(s_112_43), .b(s_112_42), .c(s_112_41), .d(s_112_40), .cin(t_2398), .o(t_2438), .co(t_2439), .cout(t_2440));
compressor_4_2 u2_838(.a(s_112_47), .b(s_112_46), .c(s_112_45), .d(s_112_44), .cin(t_2401), .o(t_2441), .co(t_2442), .cout(t_2443));
compressor_4_2 u2_839(.a(s_112_51), .b(s_112_50), .c(s_112_49), .d(s_112_48), .cin(t_2404), .o(t_2444), .co(t_2445), .cout(t_2446));
compressor_4_2 u2_840(.a(s_112_55), .b(s_112_54), .c(s_112_53), .d(s_112_52), .cin(t_2407), .o(t_2447), .co(t_2448), .cout(t_2449));
half_adder u0_841(.a(s_112_57), .b(s_112_56), .o(t_2450), .cout(t_2451));
compressor_4_2 u2_842(.a(s_113_3), .b(s_113_2), .c(s_113_1), .d(s_113_0), .cin(t_2410), .o(t_2452), .co(t_2453), .cout(t_2454));
compressor_4_2 u2_843(.a(s_113_7), .b(s_113_6), .c(s_113_5), .d(s_113_4), .cin(t_2413), .o(t_2455), .co(t_2456), .cout(t_2457));
compressor_4_2 u2_844(.a(s_113_11), .b(s_113_10), .c(s_113_9), .d(s_113_8), .cin(t_2416), .o(t_2458), .co(t_2459), .cout(t_2460));
compressor_4_2 u2_845(.a(s_113_15), .b(s_113_14), .c(s_113_13), .d(s_113_12), .cin(t_2419), .o(t_2461), .co(t_2462), .cout(t_2463));
compressor_4_2 u2_846(.a(s_113_19), .b(s_113_18), .c(s_113_17), .d(s_113_16), .cin(t_2422), .o(t_2464), .co(t_2465), .cout(t_2466));
compressor_4_2 u2_847(.a(s_113_23), .b(s_113_22), .c(s_113_21), .d(s_113_20), .cin(t_2425), .o(t_2467), .co(t_2468), .cout(t_2469));
compressor_4_2 u2_848(.a(s_113_27), .b(s_113_26), .c(s_113_25), .d(s_113_24), .cin(t_2428), .o(t_2470), .co(t_2471), .cout(t_2472));
compressor_4_2 u2_849(.a(s_113_31), .b(s_113_30), .c(s_113_29), .d(s_113_28), .cin(t_2431), .o(t_2473), .co(t_2474), .cout(t_2475));
compressor_4_2 u2_850(.a(s_113_35), .b(s_113_34), .c(s_113_33), .d(s_113_32), .cin(t_2434), .o(t_2476), .co(t_2477), .cout(t_2478));
compressor_4_2 u2_851(.a(s_113_39), .b(s_113_38), .c(s_113_37), .d(s_113_36), .cin(t_2437), .o(t_2479), .co(t_2480), .cout(t_2481));
compressor_4_2 u2_852(.a(s_113_43), .b(s_113_42), .c(s_113_41), .d(s_113_40), .cin(t_2440), .o(t_2482), .co(t_2483), .cout(t_2484));
compressor_4_2 u2_853(.a(s_113_47), .b(s_113_46), .c(s_113_45), .d(s_113_44), .cin(t_2443), .o(t_2485), .co(t_2486), .cout(t_2487));
compressor_4_2 u2_854(.a(s_113_51), .b(s_113_50), .c(s_113_49), .d(s_113_48), .cin(t_2446), .o(t_2488), .co(t_2489), .cout(t_2490));
compressor_4_2 u2_855(.a(s_113_55), .b(s_113_54), .c(s_113_53), .d(s_113_52), .cin(t_2449), .o(t_2491), .co(t_2492), .cout(t_2493));
compressor_4_2 u2_856(.a(s_114_3), .b(s_114_2), .c(s_114_1), .d(s_114_0), .cin(t_2454), .o(t_2494), .co(t_2495), .cout(t_2496));
compressor_4_2 u2_857(.a(s_114_7), .b(s_114_6), .c(s_114_5), .d(s_114_4), .cin(t_2457), .o(t_2497), .co(t_2498), .cout(t_2499));
compressor_4_2 u2_858(.a(s_114_11), .b(s_114_10), .c(s_114_9), .d(s_114_8), .cin(t_2460), .o(t_2500), .co(t_2501), .cout(t_2502));
compressor_4_2 u2_859(.a(s_114_15), .b(s_114_14), .c(s_114_13), .d(s_114_12), .cin(t_2463), .o(t_2503), .co(t_2504), .cout(t_2505));
compressor_4_2 u2_860(.a(s_114_19), .b(s_114_18), .c(s_114_17), .d(s_114_16), .cin(t_2466), .o(t_2506), .co(t_2507), .cout(t_2508));
compressor_4_2 u2_861(.a(s_114_23), .b(s_114_22), .c(s_114_21), .d(s_114_20), .cin(t_2469), .o(t_2509), .co(t_2510), .cout(t_2511));
compressor_4_2 u2_862(.a(s_114_27), .b(s_114_26), .c(s_114_25), .d(s_114_24), .cin(t_2472), .o(t_2512), .co(t_2513), .cout(t_2514));
compressor_4_2 u2_863(.a(s_114_31), .b(s_114_30), .c(s_114_29), .d(s_114_28), .cin(t_2475), .o(t_2515), .co(t_2516), .cout(t_2517));
compressor_4_2 u2_864(.a(s_114_35), .b(s_114_34), .c(s_114_33), .d(s_114_32), .cin(t_2478), .o(t_2518), .co(t_2519), .cout(t_2520));
compressor_4_2 u2_865(.a(s_114_39), .b(s_114_38), .c(s_114_37), .d(s_114_36), .cin(t_2481), .o(t_2521), .co(t_2522), .cout(t_2523));
compressor_4_2 u2_866(.a(s_114_43), .b(s_114_42), .c(s_114_41), .d(s_114_40), .cin(t_2484), .o(t_2524), .co(t_2525), .cout(t_2526));
compressor_4_2 u2_867(.a(s_114_47), .b(s_114_46), .c(s_114_45), .d(s_114_44), .cin(t_2487), .o(t_2527), .co(t_2528), .cout(t_2529));
compressor_4_2 u2_868(.a(s_114_51), .b(s_114_50), .c(s_114_49), .d(s_114_48), .cin(t_2490), .o(t_2530), .co(t_2531), .cout(t_2532));
compressor_4_2 u2_869(.a(s_114_55), .b(s_114_54), .c(s_114_53), .d(s_114_52), .cin(t_2493), .o(t_2533), .co(t_2534), .cout(t_2535));
compressor_3_2 u1_870(.a(s_114_58), .b(s_114_57), .cin(s_114_56), .o(t_2536), .cout(t_2537));
compressor_4_2 u2_871(.a(s_115_3), .b(s_115_2), .c(s_115_1), .d(s_115_0), .cin(t_2496), .o(t_2538), .co(t_2539), .cout(t_2540));
compressor_4_2 u2_872(.a(s_115_7), .b(s_115_6), .c(s_115_5), .d(s_115_4), .cin(t_2499), .o(t_2541), .co(t_2542), .cout(t_2543));
compressor_4_2 u2_873(.a(s_115_11), .b(s_115_10), .c(s_115_9), .d(s_115_8), .cin(t_2502), .o(t_2544), .co(t_2545), .cout(t_2546));
compressor_4_2 u2_874(.a(s_115_15), .b(s_115_14), .c(s_115_13), .d(s_115_12), .cin(t_2505), .o(t_2547), .co(t_2548), .cout(t_2549));
compressor_4_2 u2_875(.a(s_115_19), .b(s_115_18), .c(s_115_17), .d(s_115_16), .cin(t_2508), .o(t_2550), .co(t_2551), .cout(t_2552));
compressor_4_2 u2_876(.a(s_115_23), .b(s_115_22), .c(s_115_21), .d(s_115_20), .cin(t_2511), .o(t_2553), .co(t_2554), .cout(t_2555));
compressor_4_2 u2_877(.a(s_115_27), .b(s_115_26), .c(s_115_25), .d(s_115_24), .cin(t_2514), .o(t_2556), .co(t_2557), .cout(t_2558));
compressor_4_2 u2_878(.a(s_115_31), .b(s_115_30), .c(s_115_29), .d(s_115_28), .cin(t_2517), .o(t_2559), .co(t_2560), .cout(t_2561));
compressor_4_2 u2_879(.a(s_115_35), .b(s_115_34), .c(s_115_33), .d(s_115_32), .cin(t_2520), .o(t_2562), .co(t_2563), .cout(t_2564));
compressor_4_2 u2_880(.a(s_115_39), .b(s_115_38), .c(s_115_37), .d(s_115_36), .cin(t_2523), .o(t_2565), .co(t_2566), .cout(t_2567));
compressor_4_2 u2_881(.a(s_115_43), .b(s_115_42), .c(s_115_41), .d(s_115_40), .cin(t_2526), .o(t_2568), .co(t_2569), .cout(t_2570));
compressor_4_2 u2_882(.a(s_115_47), .b(s_115_46), .c(s_115_45), .d(s_115_44), .cin(t_2529), .o(t_2571), .co(t_2572), .cout(t_2573));
compressor_4_2 u2_883(.a(s_115_51), .b(s_115_50), .c(s_115_49), .d(s_115_48), .cin(t_2532), .o(t_2574), .co(t_2575), .cout(t_2576));
compressor_4_2 u2_884(.a(s_115_55), .b(s_115_54), .c(s_115_53), .d(s_115_52), .cin(t_2535), .o(t_2577), .co(t_2578), .cout(t_2579));
half_adder u0_885(.a(s_115_57), .b(s_115_56), .o(t_2580), .cout(t_2581));
compressor_4_2 u2_886(.a(s_116_3), .b(s_116_2), .c(s_116_1), .d(s_116_0), .cin(t_2540), .o(t_2582), .co(t_2583), .cout(t_2584));
compressor_4_2 u2_887(.a(s_116_7), .b(s_116_6), .c(s_116_5), .d(s_116_4), .cin(t_2543), .o(t_2585), .co(t_2586), .cout(t_2587));
compressor_4_2 u2_888(.a(s_116_11), .b(s_116_10), .c(s_116_9), .d(s_116_8), .cin(t_2546), .o(t_2588), .co(t_2589), .cout(t_2590));
compressor_4_2 u2_889(.a(s_116_15), .b(s_116_14), .c(s_116_13), .d(s_116_12), .cin(t_2549), .o(t_2591), .co(t_2592), .cout(t_2593));
compressor_4_2 u2_890(.a(s_116_19), .b(s_116_18), .c(s_116_17), .d(s_116_16), .cin(t_2552), .o(t_2594), .co(t_2595), .cout(t_2596));
compressor_4_2 u2_891(.a(s_116_23), .b(s_116_22), .c(s_116_21), .d(s_116_20), .cin(t_2555), .o(t_2597), .co(t_2598), .cout(t_2599));
compressor_4_2 u2_892(.a(s_116_27), .b(s_116_26), .c(s_116_25), .d(s_116_24), .cin(t_2558), .o(t_2600), .co(t_2601), .cout(t_2602));
compressor_4_2 u2_893(.a(s_116_31), .b(s_116_30), .c(s_116_29), .d(s_116_28), .cin(t_2561), .o(t_2603), .co(t_2604), .cout(t_2605));
compressor_4_2 u2_894(.a(s_116_35), .b(s_116_34), .c(s_116_33), .d(s_116_32), .cin(t_2564), .o(t_2606), .co(t_2607), .cout(t_2608));
compressor_4_2 u2_895(.a(s_116_39), .b(s_116_38), .c(s_116_37), .d(s_116_36), .cin(t_2567), .o(t_2609), .co(t_2610), .cout(t_2611));
compressor_4_2 u2_896(.a(s_116_43), .b(s_116_42), .c(s_116_41), .d(s_116_40), .cin(t_2570), .o(t_2612), .co(t_2613), .cout(t_2614));
compressor_4_2 u2_897(.a(s_116_47), .b(s_116_46), .c(s_116_45), .d(s_116_44), .cin(t_2573), .o(t_2615), .co(t_2616), .cout(t_2617));
compressor_4_2 u2_898(.a(s_116_51), .b(s_116_50), .c(s_116_49), .d(s_116_48), .cin(t_2576), .o(t_2618), .co(t_2619), .cout(t_2620));
compressor_4_2 u2_899(.a(s_116_55), .b(s_116_54), .c(s_116_53), .d(s_116_52), .cin(t_2579), .o(t_2621), .co(t_2622), .cout(t_2623));
compressor_3_2 u1_900(.a(s_116_58), .b(s_116_57), .cin(s_116_56), .o(t_2624), .cout(t_2625));
compressor_4_2 u2_901(.a(s_117_3), .b(s_117_2), .c(s_117_1), .d(s_117_0), .cin(t_2584), .o(t_2626), .co(t_2627), .cout(t_2628));
compressor_4_2 u2_902(.a(s_117_7), .b(s_117_6), .c(s_117_5), .d(s_117_4), .cin(t_2587), .o(t_2629), .co(t_2630), .cout(t_2631));
compressor_4_2 u2_903(.a(s_117_11), .b(s_117_10), .c(s_117_9), .d(s_117_8), .cin(t_2590), .o(t_2632), .co(t_2633), .cout(t_2634));
compressor_4_2 u2_904(.a(s_117_15), .b(s_117_14), .c(s_117_13), .d(s_117_12), .cin(t_2593), .o(t_2635), .co(t_2636), .cout(t_2637));
compressor_4_2 u2_905(.a(s_117_19), .b(s_117_18), .c(s_117_17), .d(s_117_16), .cin(t_2596), .o(t_2638), .co(t_2639), .cout(t_2640));
compressor_4_2 u2_906(.a(s_117_23), .b(s_117_22), .c(s_117_21), .d(s_117_20), .cin(t_2599), .o(t_2641), .co(t_2642), .cout(t_2643));
compressor_4_2 u2_907(.a(s_117_27), .b(s_117_26), .c(s_117_25), .d(s_117_24), .cin(t_2602), .o(t_2644), .co(t_2645), .cout(t_2646));
compressor_4_2 u2_908(.a(s_117_31), .b(s_117_30), .c(s_117_29), .d(s_117_28), .cin(t_2605), .o(t_2647), .co(t_2648), .cout(t_2649));
compressor_4_2 u2_909(.a(s_117_35), .b(s_117_34), .c(s_117_33), .d(s_117_32), .cin(t_2608), .o(t_2650), .co(t_2651), .cout(t_2652));
compressor_4_2 u2_910(.a(s_117_39), .b(s_117_38), .c(s_117_37), .d(s_117_36), .cin(t_2611), .o(t_2653), .co(t_2654), .cout(t_2655));
compressor_4_2 u2_911(.a(s_117_43), .b(s_117_42), .c(s_117_41), .d(s_117_40), .cin(t_2614), .o(t_2656), .co(t_2657), .cout(t_2658));
compressor_4_2 u2_912(.a(s_117_47), .b(s_117_46), .c(s_117_45), .d(s_117_44), .cin(t_2617), .o(t_2659), .co(t_2660), .cout(t_2661));
compressor_4_2 u2_913(.a(s_117_51), .b(s_117_50), .c(s_117_49), .d(s_117_48), .cin(t_2620), .o(t_2662), .co(t_2663), .cout(t_2664));
compressor_4_2 u2_914(.a(s_117_55), .b(s_117_54), .c(s_117_53), .d(s_117_52), .cin(t_2623), .o(t_2665), .co(t_2666), .cout(t_2667));
compressor_3_2 u1_915(.a(s_117_58), .b(s_117_57), .cin(s_117_56), .o(t_2668), .cout(t_2669));
compressor_4_2 u2_916(.a(s_118_3), .b(s_118_2), .c(s_118_1), .d(s_118_0), .cin(t_2628), .o(t_2670), .co(t_2671), .cout(t_2672));
compressor_4_2 u2_917(.a(s_118_7), .b(s_118_6), .c(s_118_5), .d(s_118_4), .cin(t_2631), .o(t_2673), .co(t_2674), .cout(t_2675));
compressor_4_2 u2_918(.a(s_118_11), .b(s_118_10), .c(s_118_9), .d(s_118_8), .cin(t_2634), .o(t_2676), .co(t_2677), .cout(t_2678));
compressor_4_2 u2_919(.a(s_118_15), .b(s_118_14), .c(s_118_13), .d(s_118_12), .cin(t_2637), .o(t_2679), .co(t_2680), .cout(t_2681));
compressor_4_2 u2_920(.a(s_118_19), .b(s_118_18), .c(s_118_17), .d(s_118_16), .cin(t_2640), .o(t_2682), .co(t_2683), .cout(t_2684));
compressor_4_2 u2_921(.a(s_118_23), .b(s_118_22), .c(s_118_21), .d(s_118_20), .cin(t_2643), .o(t_2685), .co(t_2686), .cout(t_2687));
compressor_4_2 u2_922(.a(s_118_27), .b(s_118_26), .c(s_118_25), .d(s_118_24), .cin(t_2646), .o(t_2688), .co(t_2689), .cout(t_2690));
compressor_4_2 u2_923(.a(s_118_31), .b(s_118_30), .c(s_118_29), .d(s_118_28), .cin(t_2649), .o(t_2691), .co(t_2692), .cout(t_2693));
compressor_4_2 u2_924(.a(s_118_35), .b(s_118_34), .c(s_118_33), .d(s_118_32), .cin(t_2652), .o(t_2694), .co(t_2695), .cout(t_2696));
compressor_4_2 u2_925(.a(s_118_39), .b(s_118_38), .c(s_118_37), .d(s_118_36), .cin(t_2655), .o(t_2697), .co(t_2698), .cout(t_2699));
compressor_4_2 u2_926(.a(s_118_43), .b(s_118_42), .c(s_118_41), .d(s_118_40), .cin(t_2658), .o(t_2700), .co(t_2701), .cout(t_2702));
compressor_4_2 u2_927(.a(s_118_47), .b(s_118_46), .c(s_118_45), .d(s_118_44), .cin(t_2661), .o(t_2703), .co(t_2704), .cout(t_2705));
compressor_4_2 u2_928(.a(s_118_51), .b(s_118_50), .c(s_118_49), .d(s_118_48), .cin(t_2664), .o(t_2706), .co(t_2707), .cout(t_2708));
compressor_4_2 u2_929(.a(s_118_55), .b(s_118_54), .c(s_118_53), .d(s_118_52), .cin(t_2667), .o(t_2709), .co(t_2710), .cout(t_2711));
compressor_4_2 u2_930(.a(s_118_60), .b(s_118_59), .c(s_118_58), .d(s_118_57), .cin(s_118_56), .o(t_2712), .co(t_2713), .cout(t_2714));
compressor_4_2 u2_931(.a(s_119_3), .b(s_119_2), .c(s_119_1), .d(s_119_0), .cin(t_2672), .o(t_2715), .co(t_2716), .cout(t_2717));
compressor_4_2 u2_932(.a(s_119_7), .b(s_119_6), .c(s_119_5), .d(s_119_4), .cin(t_2675), .o(t_2718), .co(t_2719), .cout(t_2720));
compressor_4_2 u2_933(.a(s_119_11), .b(s_119_10), .c(s_119_9), .d(s_119_8), .cin(t_2678), .o(t_2721), .co(t_2722), .cout(t_2723));
compressor_4_2 u2_934(.a(s_119_15), .b(s_119_14), .c(s_119_13), .d(s_119_12), .cin(t_2681), .o(t_2724), .co(t_2725), .cout(t_2726));
compressor_4_2 u2_935(.a(s_119_19), .b(s_119_18), .c(s_119_17), .d(s_119_16), .cin(t_2684), .o(t_2727), .co(t_2728), .cout(t_2729));
compressor_4_2 u2_936(.a(s_119_23), .b(s_119_22), .c(s_119_21), .d(s_119_20), .cin(t_2687), .o(t_2730), .co(t_2731), .cout(t_2732));
compressor_4_2 u2_937(.a(s_119_27), .b(s_119_26), .c(s_119_25), .d(s_119_24), .cin(t_2690), .o(t_2733), .co(t_2734), .cout(t_2735));
compressor_4_2 u2_938(.a(s_119_31), .b(s_119_30), .c(s_119_29), .d(s_119_28), .cin(t_2693), .o(t_2736), .co(t_2737), .cout(t_2738));
compressor_4_2 u2_939(.a(s_119_35), .b(s_119_34), .c(s_119_33), .d(s_119_32), .cin(t_2696), .o(t_2739), .co(t_2740), .cout(t_2741));
compressor_4_2 u2_940(.a(s_119_39), .b(s_119_38), .c(s_119_37), .d(s_119_36), .cin(t_2699), .o(t_2742), .co(t_2743), .cout(t_2744));
compressor_4_2 u2_941(.a(s_119_43), .b(s_119_42), .c(s_119_41), .d(s_119_40), .cin(t_2702), .o(t_2745), .co(t_2746), .cout(t_2747));
compressor_4_2 u2_942(.a(s_119_47), .b(s_119_46), .c(s_119_45), .d(s_119_44), .cin(t_2705), .o(t_2748), .co(t_2749), .cout(t_2750));
compressor_4_2 u2_943(.a(s_119_51), .b(s_119_50), .c(s_119_49), .d(s_119_48), .cin(t_2708), .o(t_2751), .co(t_2752), .cout(t_2753));
compressor_4_2 u2_944(.a(s_119_55), .b(s_119_54), .c(s_119_53), .d(s_119_52), .cin(t_2711), .o(t_2754), .co(t_2755), .cout(t_2756));
compressor_4_2 u2_945(.a(s_119_59), .b(s_119_58), .c(s_119_57), .d(s_119_56), .cin(t_2714), .o(t_2757), .co(t_2758), .cout(t_2759));
compressor_4_2 u2_946(.a(s_120_3), .b(s_120_2), .c(s_120_1), .d(s_120_0), .cin(t_2717), .o(t_2760), .co(t_2761), .cout(t_2762));
compressor_4_2 u2_947(.a(s_120_7), .b(s_120_6), .c(s_120_5), .d(s_120_4), .cin(t_2720), .o(t_2763), .co(t_2764), .cout(t_2765));
compressor_4_2 u2_948(.a(s_120_11), .b(s_120_10), .c(s_120_9), .d(s_120_8), .cin(t_2723), .o(t_2766), .co(t_2767), .cout(t_2768));
compressor_4_2 u2_949(.a(s_120_15), .b(s_120_14), .c(s_120_13), .d(s_120_12), .cin(t_2726), .o(t_2769), .co(t_2770), .cout(t_2771));
compressor_4_2 u2_950(.a(s_120_19), .b(s_120_18), .c(s_120_17), .d(s_120_16), .cin(t_2729), .o(t_2772), .co(t_2773), .cout(t_2774));
compressor_4_2 u2_951(.a(s_120_23), .b(s_120_22), .c(s_120_21), .d(s_120_20), .cin(t_2732), .o(t_2775), .co(t_2776), .cout(t_2777));
compressor_4_2 u2_952(.a(s_120_27), .b(s_120_26), .c(s_120_25), .d(s_120_24), .cin(t_2735), .o(t_2778), .co(t_2779), .cout(t_2780));
compressor_4_2 u2_953(.a(s_120_31), .b(s_120_30), .c(s_120_29), .d(s_120_28), .cin(t_2738), .o(t_2781), .co(t_2782), .cout(t_2783));
compressor_4_2 u2_954(.a(s_120_35), .b(s_120_34), .c(s_120_33), .d(s_120_32), .cin(t_2741), .o(t_2784), .co(t_2785), .cout(t_2786));
compressor_4_2 u2_955(.a(s_120_39), .b(s_120_38), .c(s_120_37), .d(s_120_36), .cin(t_2744), .o(t_2787), .co(t_2788), .cout(t_2789));
compressor_4_2 u2_956(.a(s_120_43), .b(s_120_42), .c(s_120_41), .d(s_120_40), .cin(t_2747), .o(t_2790), .co(t_2791), .cout(t_2792));
compressor_4_2 u2_957(.a(s_120_47), .b(s_120_46), .c(s_120_45), .d(s_120_44), .cin(t_2750), .o(t_2793), .co(t_2794), .cout(t_2795));
compressor_4_2 u2_958(.a(s_120_51), .b(s_120_50), .c(s_120_49), .d(s_120_48), .cin(t_2753), .o(t_2796), .co(t_2797), .cout(t_2798));
compressor_4_2 u2_959(.a(s_120_55), .b(s_120_54), .c(s_120_53), .d(s_120_52), .cin(t_2756), .o(t_2799), .co(t_2800), .cout(t_2801));
compressor_4_2 u2_960(.a(s_120_59), .b(s_120_58), .c(s_120_57), .d(s_120_56), .cin(t_2759), .o(t_2802), .co(t_2803), .cout(t_2804));
half_adder u0_961(.a(s_120_61), .b(s_120_60), .o(t_2805), .cout(t_2806));
compressor_4_2 u2_962(.a(s_121_3), .b(s_121_2), .c(s_121_1), .d(s_121_0), .cin(t_2762), .o(t_2807), .co(t_2808), .cout(t_2809));
compressor_4_2 u2_963(.a(s_121_7), .b(s_121_6), .c(s_121_5), .d(s_121_4), .cin(t_2765), .o(t_2810), .co(t_2811), .cout(t_2812));
compressor_4_2 u2_964(.a(s_121_11), .b(s_121_10), .c(s_121_9), .d(s_121_8), .cin(t_2768), .o(t_2813), .co(t_2814), .cout(t_2815));
compressor_4_2 u2_965(.a(s_121_15), .b(s_121_14), .c(s_121_13), .d(s_121_12), .cin(t_2771), .o(t_2816), .co(t_2817), .cout(t_2818));
compressor_4_2 u2_966(.a(s_121_19), .b(s_121_18), .c(s_121_17), .d(s_121_16), .cin(t_2774), .o(t_2819), .co(t_2820), .cout(t_2821));
compressor_4_2 u2_967(.a(s_121_23), .b(s_121_22), .c(s_121_21), .d(s_121_20), .cin(t_2777), .o(t_2822), .co(t_2823), .cout(t_2824));
compressor_4_2 u2_968(.a(s_121_27), .b(s_121_26), .c(s_121_25), .d(s_121_24), .cin(t_2780), .o(t_2825), .co(t_2826), .cout(t_2827));
compressor_4_2 u2_969(.a(s_121_31), .b(s_121_30), .c(s_121_29), .d(s_121_28), .cin(t_2783), .o(t_2828), .co(t_2829), .cout(t_2830));
compressor_4_2 u2_970(.a(s_121_35), .b(s_121_34), .c(s_121_33), .d(s_121_32), .cin(t_2786), .o(t_2831), .co(t_2832), .cout(t_2833));
compressor_4_2 u2_971(.a(s_121_39), .b(s_121_38), .c(s_121_37), .d(s_121_36), .cin(t_2789), .o(t_2834), .co(t_2835), .cout(t_2836));
compressor_4_2 u2_972(.a(s_121_43), .b(s_121_42), .c(s_121_41), .d(s_121_40), .cin(t_2792), .o(t_2837), .co(t_2838), .cout(t_2839));
compressor_4_2 u2_973(.a(s_121_47), .b(s_121_46), .c(s_121_45), .d(s_121_44), .cin(t_2795), .o(t_2840), .co(t_2841), .cout(t_2842));
compressor_4_2 u2_974(.a(s_121_51), .b(s_121_50), .c(s_121_49), .d(s_121_48), .cin(t_2798), .o(t_2843), .co(t_2844), .cout(t_2845));
compressor_4_2 u2_975(.a(s_121_55), .b(s_121_54), .c(s_121_53), .d(s_121_52), .cin(t_2801), .o(t_2846), .co(t_2847), .cout(t_2848));
compressor_4_2 u2_976(.a(s_121_59), .b(s_121_58), .c(s_121_57), .d(s_121_56), .cin(t_2804), .o(t_2849), .co(t_2850), .cout(t_2851));
compressor_4_2 u2_977(.a(s_122_3), .b(s_122_2), .c(s_122_1), .d(s_122_0), .cin(t_2809), .o(t_2852), .co(t_2853), .cout(t_2854));
compressor_4_2 u2_978(.a(s_122_7), .b(s_122_6), .c(s_122_5), .d(s_122_4), .cin(t_2812), .o(t_2855), .co(t_2856), .cout(t_2857));
compressor_4_2 u2_979(.a(s_122_11), .b(s_122_10), .c(s_122_9), .d(s_122_8), .cin(t_2815), .o(t_2858), .co(t_2859), .cout(t_2860));
compressor_4_2 u2_980(.a(s_122_15), .b(s_122_14), .c(s_122_13), .d(s_122_12), .cin(t_2818), .o(t_2861), .co(t_2862), .cout(t_2863));
compressor_4_2 u2_981(.a(s_122_19), .b(s_122_18), .c(s_122_17), .d(s_122_16), .cin(t_2821), .o(t_2864), .co(t_2865), .cout(t_2866));
compressor_4_2 u2_982(.a(s_122_23), .b(s_122_22), .c(s_122_21), .d(s_122_20), .cin(t_2824), .o(t_2867), .co(t_2868), .cout(t_2869));
compressor_4_2 u2_983(.a(s_122_27), .b(s_122_26), .c(s_122_25), .d(s_122_24), .cin(t_2827), .o(t_2870), .co(t_2871), .cout(t_2872));
compressor_4_2 u2_984(.a(s_122_31), .b(s_122_30), .c(s_122_29), .d(s_122_28), .cin(t_2830), .o(t_2873), .co(t_2874), .cout(t_2875));
compressor_4_2 u2_985(.a(s_122_35), .b(s_122_34), .c(s_122_33), .d(s_122_32), .cin(t_2833), .o(t_2876), .co(t_2877), .cout(t_2878));
compressor_4_2 u2_986(.a(s_122_39), .b(s_122_38), .c(s_122_37), .d(s_122_36), .cin(t_2836), .o(t_2879), .co(t_2880), .cout(t_2881));
compressor_4_2 u2_987(.a(s_122_43), .b(s_122_42), .c(s_122_41), .d(s_122_40), .cin(t_2839), .o(t_2882), .co(t_2883), .cout(t_2884));
compressor_4_2 u2_988(.a(s_122_47), .b(s_122_46), .c(s_122_45), .d(s_122_44), .cin(t_2842), .o(t_2885), .co(t_2886), .cout(t_2887));
compressor_4_2 u2_989(.a(s_122_51), .b(s_122_50), .c(s_122_49), .d(s_122_48), .cin(t_2845), .o(t_2888), .co(t_2889), .cout(t_2890));
compressor_4_2 u2_990(.a(s_122_55), .b(s_122_54), .c(s_122_53), .d(s_122_52), .cin(t_2848), .o(t_2891), .co(t_2892), .cout(t_2893));
compressor_4_2 u2_991(.a(s_122_59), .b(s_122_58), .c(s_122_57), .d(s_122_56), .cin(t_2851), .o(t_2894), .co(t_2895), .cout(t_2896));
compressor_3_2 u1_992(.a(s_122_62), .b(s_122_61), .cin(s_122_60), .o(t_2897), .cout(t_2898));
compressor_4_2 u2_993(.a(s_123_3), .b(s_123_2), .c(s_123_1), .d(s_123_0), .cin(t_2854), .o(t_2899), .co(t_2900), .cout(t_2901));
compressor_4_2 u2_994(.a(s_123_7), .b(s_123_6), .c(s_123_5), .d(s_123_4), .cin(t_2857), .o(t_2902), .co(t_2903), .cout(t_2904));
compressor_4_2 u2_995(.a(s_123_11), .b(s_123_10), .c(s_123_9), .d(s_123_8), .cin(t_2860), .o(t_2905), .co(t_2906), .cout(t_2907));
compressor_4_2 u2_996(.a(s_123_15), .b(s_123_14), .c(s_123_13), .d(s_123_12), .cin(t_2863), .o(t_2908), .co(t_2909), .cout(t_2910));
compressor_4_2 u2_997(.a(s_123_19), .b(s_123_18), .c(s_123_17), .d(s_123_16), .cin(t_2866), .o(t_2911), .co(t_2912), .cout(t_2913));
compressor_4_2 u2_998(.a(s_123_23), .b(s_123_22), .c(s_123_21), .d(s_123_20), .cin(t_2869), .o(t_2914), .co(t_2915), .cout(t_2916));
compressor_4_2 u2_999(.a(s_123_27), .b(s_123_26), .c(s_123_25), .d(s_123_24), .cin(t_2872), .o(t_2917), .co(t_2918), .cout(t_2919));
compressor_4_2 u2_1000(.a(s_123_31), .b(s_123_30), .c(s_123_29), .d(s_123_28), .cin(t_2875), .o(t_2920), .co(t_2921), .cout(t_2922));
compressor_4_2 u2_1001(.a(s_123_35), .b(s_123_34), .c(s_123_33), .d(s_123_32), .cin(t_2878), .o(t_2923), .co(t_2924), .cout(t_2925));
compressor_4_2 u2_1002(.a(s_123_39), .b(s_123_38), .c(s_123_37), .d(s_123_36), .cin(t_2881), .o(t_2926), .co(t_2927), .cout(t_2928));
compressor_4_2 u2_1003(.a(s_123_43), .b(s_123_42), .c(s_123_41), .d(s_123_40), .cin(t_2884), .o(t_2929), .co(t_2930), .cout(t_2931));
compressor_4_2 u2_1004(.a(s_123_47), .b(s_123_46), .c(s_123_45), .d(s_123_44), .cin(t_2887), .o(t_2932), .co(t_2933), .cout(t_2934));
compressor_4_2 u2_1005(.a(s_123_51), .b(s_123_50), .c(s_123_49), .d(s_123_48), .cin(t_2890), .o(t_2935), .co(t_2936), .cout(t_2937));
compressor_4_2 u2_1006(.a(s_123_55), .b(s_123_54), .c(s_123_53), .d(s_123_52), .cin(t_2893), .o(t_2938), .co(t_2939), .cout(t_2940));
compressor_4_2 u2_1007(.a(s_123_59), .b(s_123_58), .c(s_123_57), .d(s_123_56), .cin(t_2896), .o(t_2941), .co(t_2942), .cout(t_2943));
half_adder u0_1008(.a(s_123_61), .b(s_123_60), .o(t_2944), .cout(t_2945));
compressor_4_2 u2_1009(.a(s_124_3), .b(s_124_2), .c(s_124_1), .d(s_124_0), .cin(t_2901), .o(t_2946), .co(t_2947), .cout(t_2948));
compressor_4_2 u2_1010(.a(s_124_7), .b(s_124_6), .c(s_124_5), .d(s_124_4), .cin(t_2904), .o(t_2949), .co(t_2950), .cout(t_2951));
compressor_4_2 u2_1011(.a(s_124_11), .b(s_124_10), .c(s_124_9), .d(s_124_8), .cin(t_2907), .o(t_2952), .co(t_2953), .cout(t_2954));
compressor_4_2 u2_1012(.a(s_124_15), .b(s_124_14), .c(s_124_13), .d(s_124_12), .cin(t_2910), .o(t_2955), .co(t_2956), .cout(t_2957));
compressor_4_2 u2_1013(.a(s_124_19), .b(s_124_18), .c(s_124_17), .d(s_124_16), .cin(t_2913), .o(t_2958), .co(t_2959), .cout(t_2960));
compressor_4_2 u2_1014(.a(s_124_23), .b(s_124_22), .c(s_124_21), .d(s_124_20), .cin(t_2916), .o(t_2961), .co(t_2962), .cout(t_2963));
compressor_4_2 u2_1015(.a(s_124_27), .b(s_124_26), .c(s_124_25), .d(s_124_24), .cin(t_2919), .o(t_2964), .co(t_2965), .cout(t_2966));
compressor_4_2 u2_1016(.a(s_124_31), .b(s_124_30), .c(s_124_29), .d(s_124_28), .cin(t_2922), .o(t_2967), .co(t_2968), .cout(t_2969));
compressor_4_2 u2_1017(.a(s_124_35), .b(s_124_34), .c(s_124_33), .d(s_124_32), .cin(t_2925), .o(t_2970), .co(t_2971), .cout(t_2972));
compressor_4_2 u2_1018(.a(s_124_39), .b(s_124_38), .c(s_124_37), .d(s_124_36), .cin(t_2928), .o(t_2973), .co(t_2974), .cout(t_2975));
compressor_4_2 u2_1019(.a(s_124_43), .b(s_124_42), .c(s_124_41), .d(s_124_40), .cin(t_2931), .o(t_2976), .co(t_2977), .cout(t_2978));
compressor_4_2 u2_1020(.a(s_124_47), .b(s_124_46), .c(s_124_45), .d(s_124_44), .cin(t_2934), .o(t_2979), .co(t_2980), .cout(t_2981));
compressor_4_2 u2_1021(.a(s_124_51), .b(s_124_50), .c(s_124_49), .d(s_124_48), .cin(t_2937), .o(t_2982), .co(t_2983), .cout(t_2984));
compressor_4_2 u2_1022(.a(s_124_55), .b(s_124_54), .c(s_124_53), .d(s_124_52), .cin(t_2940), .o(t_2985), .co(t_2986), .cout(t_2987));
compressor_4_2 u2_1023(.a(s_124_59), .b(s_124_58), .c(s_124_57), .d(s_124_56), .cin(t_2943), .o(t_2988), .co(t_2989), .cout(t_2990));
compressor_3_2 u1_1024(.a(s_124_62), .b(s_124_61), .cin(s_124_60), .o(t_2991), .cout(t_2992));
compressor_4_2 u2_1025(.a(s_125_3), .b(s_125_2), .c(s_125_1), .d(s_125_0), .cin(t_2948), .o(t_2993), .co(t_2994), .cout(t_2995));
compressor_4_2 u2_1026(.a(s_125_7), .b(s_125_6), .c(s_125_5), .d(s_125_4), .cin(t_2951), .o(t_2996), .co(t_2997), .cout(t_2998));
compressor_4_2 u2_1027(.a(s_125_11), .b(s_125_10), .c(s_125_9), .d(s_125_8), .cin(t_2954), .o(t_2999), .co(t_3000), .cout(t_3001));
compressor_4_2 u2_1028(.a(s_125_15), .b(s_125_14), .c(s_125_13), .d(s_125_12), .cin(t_2957), .o(t_3002), .co(t_3003), .cout(t_3004));
compressor_4_2 u2_1029(.a(s_125_19), .b(s_125_18), .c(s_125_17), .d(s_125_16), .cin(t_2960), .o(t_3005), .co(t_3006), .cout(t_3007));
compressor_4_2 u2_1030(.a(s_125_23), .b(s_125_22), .c(s_125_21), .d(s_125_20), .cin(t_2963), .o(t_3008), .co(t_3009), .cout(t_3010));
compressor_4_2 u2_1031(.a(s_125_27), .b(s_125_26), .c(s_125_25), .d(s_125_24), .cin(t_2966), .o(t_3011), .co(t_3012), .cout(t_3013));
compressor_4_2 u2_1032(.a(s_125_31), .b(s_125_30), .c(s_125_29), .d(s_125_28), .cin(t_2969), .o(t_3014), .co(t_3015), .cout(t_3016));
compressor_4_2 u2_1033(.a(s_125_35), .b(s_125_34), .c(s_125_33), .d(s_125_32), .cin(t_2972), .o(t_3017), .co(t_3018), .cout(t_3019));
compressor_4_2 u2_1034(.a(s_125_39), .b(s_125_38), .c(s_125_37), .d(s_125_36), .cin(t_2975), .o(t_3020), .co(t_3021), .cout(t_3022));
compressor_4_2 u2_1035(.a(s_125_43), .b(s_125_42), .c(s_125_41), .d(s_125_40), .cin(t_2978), .o(t_3023), .co(t_3024), .cout(t_3025));
compressor_4_2 u2_1036(.a(s_125_47), .b(s_125_46), .c(s_125_45), .d(s_125_44), .cin(t_2981), .o(t_3026), .co(t_3027), .cout(t_3028));
compressor_4_2 u2_1037(.a(s_125_51), .b(s_125_50), .c(s_125_49), .d(s_125_48), .cin(t_2984), .o(t_3029), .co(t_3030), .cout(t_3031));
compressor_4_2 u2_1038(.a(s_125_55), .b(s_125_54), .c(s_125_53), .d(s_125_52), .cin(t_2987), .o(t_3032), .co(t_3033), .cout(t_3034));
compressor_4_2 u2_1039(.a(s_125_59), .b(s_125_58), .c(s_125_57), .d(s_125_56), .cin(t_2990), .o(t_3035), .co(t_3036), .cout(t_3037));
compressor_3_2 u1_1040(.a(s_125_62), .b(s_125_61), .cin(s_125_60), .o(t_3038), .cout(t_3039));
compressor_4_2 u2_1041(.a(s_126_3), .b(s_126_2), .c(s_126_1), .d(s_126_0), .cin(t_2995), .o(t_3040), .co(t_3041), .cout(t_3042));
compressor_4_2 u2_1042(.a(s_126_7), .b(s_126_6), .c(s_126_5), .d(s_126_4), .cin(t_2998), .o(t_3043), .co(t_3044), .cout(t_3045));
compressor_4_2 u2_1043(.a(s_126_11), .b(s_126_10), .c(s_126_9), .d(s_126_8), .cin(t_3001), .o(t_3046), .co(t_3047), .cout(t_3048));
compressor_4_2 u2_1044(.a(s_126_15), .b(s_126_14), .c(s_126_13), .d(s_126_12), .cin(t_3004), .o(t_3049), .co(t_3050), .cout(t_3051));
compressor_4_2 u2_1045(.a(s_126_19), .b(s_126_18), .c(s_126_17), .d(s_126_16), .cin(t_3007), .o(t_3052), .co(t_3053), .cout(t_3054));
compressor_4_2 u2_1046(.a(s_126_23), .b(s_126_22), .c(s_126_21), .d(s_126_20), .cin(t_3010), .o(t_3055), .co(t_3056), .cout(t_3057));
compressor_4_2 u2_1047(.a(s_126_27), .b(s_126_26), .c(s_126_25), .d(s_126_24), .cin(t_3013), .o(t_3058), .co(t_3059), .cout(t_3060));
compressor_4_2 u2_1048(.a(s_126_31), .b(s_126_30), .c(s_126_29), .d(s_126_28), .cin(t_3016), .o(t_3061), .co(t_3062), .cout(t_3063));
compressor_4_2 u2_1049(.a(s_126_35), .b(s_126_34), .c(s_126_33), .d(s_126_32), .cin(t_3019), .o(t_3064), .co(t_3065), .cout(t_3066));
compressor_4_2 u2_1050(.a(s_126_39), .b(s_126_38), .c(s_126_37), .d(s_126_36), .cin(t_3022), .o(t_3067), .co(t_3068), .cout(t_3069));
compressor_4_2 u2_1051(.a(s_126_43), .b(s_126_42), .c(s_126_41), .d(s_126_40), .cin(t_3025), .o(t_3070), .co(t_3071), .cout(t_3072));
compressor_4_2 u2_1052(.a(s_126_47), .b(s_126_46), .c(s_126_45), .d(s_126_44), .cin(t_3028), .o(t_3073), .co(t_3074), .cout(t_3075));
compressor_4_2 u2_1053(.a(s_126_51), .b(s_126_50), .c(s_126_49), .d(s_126_48), .cin(t_3031), .o(t_3076), .co(t_3077), .cout(t_3078));
compressor_4_2 u2_1054(.a(s_126_55), .b(s_126_54), .c(s_126_53), .d(s_126_52), .cin(t_3034), .o(t_3079), .co(t_3080), .cout(t_3081));
compressor_4_2 u2_1055(.a(s_126_59), .b(s_126_58), .c(s_126_57), .d(s_126_56), .cin(t_3037), .o(t_3082), .co(t_3083), .cout(t_3084));
compressor_4_2 u2_1056(.a(s_126_64), .b(s_126_63), .c(s_126_62), .d(s_126_61), .cin(s_126_60), .o(t_3085), .co(t_3086), .cout(t_3087));
compressor_4_2 u2_1057(.a(s_127_3), .b(s_127_2), .c(s_127_1), .d(s_127_0), .cin(t_3042), .o(t_3088), .co(t_3089), .cout(t_3090));
compressor_4_2 u2_1058(.a(s_127_7), .b(s_127_6), .c(s_127_5), .d(s_127_4), .cin(t_3045), .o(t_3091), .co(t_3092), .cout(t_3093));
compressor_4_2 u2_1059(.a(s_127_11), .b(s_127_10), .c(s_127_9), .d(s_127_8), .cin(t_3048), .o(t_3094), .co(t_3095), .cout(t_3096));
compressor_4_2 u2_1060(.a(s_127_15), .b(s_127_14), .c(s_127_13), .d(s_127_12), .cin(t_3051), .o(t_3097), .co(t_3098), .cout(t_3099));
compressor_4_2 u2_1061(.a(s_127_19), .b(s_127_18), .c(s_127_17), .d(s_127_16), .cin(t_3054), .o(t_3100), .co(t_3101), .cout(t_3102));
compressor_4_2 u2_1062(.a(s_127_23), .b(s_127_22), .c(s_127_21), .d(s_127_20), .cin(t_3057), .o(t_3103), .co(t_3104), .cout(t_3105));
compressor_4_2 u2_1063(.a(s_127_27), .b(s_127_26), .c(s_127_25), .d(s_127_24), .cin(t_3060), .o(t_3106), .co(t_3107), .cout(t_3108));
compressor_4_2 u2_1064(.a(s_127_31), .b(s_127_30), .c(s_127_29), .d(s_127_28), .cin(t_3063), .o(t_3109), .co(t_3110), .cout(t_3111));
compressor_4_2 u2_1065(.a(s_127_35), .b(s_127_34), .c(s_127_33), .d(s_127_32), .cin(t_3066), .o(t_3112), .co(t_3113), .cout(t_3114));
compressor_4_2 u2_1066(.a(s_127_39), .b(s_127_38), .c(s_127_37), .d(s_127_36), .cin(t_3069), .o(t_3115), .co(t_3116), .cout(t_3117));
compressor_4_2 u2_1067(.a(s_127_43), .b(s_127_42), .c(s_127_41), .d(s_127_40), .cin(t_3072), .o(t_3118), .co(t_3119), .cout(t_3120));
compressor_4_2 u2_1068(.a(s_127_47), .b(s_127_46), .c(s_127_45), .d(s_127_44), .cin(t_3075), .o(t_3121), .co(t_3122), .cout(t_3123));
compressor_4_2 u2_1069(.a(s_127_51), .b(s_127_50), .c(s_127_49), .d(s_127_48), .cin(t_3078), .o(t_3124), .co(t_3125), .cout(t_3126));
compressor_4_2 u2_1070(.a(s_127_55), .b(s_127_54), .c(s_127_53), .d(s_127_52), .cin(t_3081), .o(t_3127), .co(t_3128), .cout(t_3129));
compressor_4_2 u2_1071(.a(s_127_59), .b(s_127_58), .c(s_127_57), .d(s_127_56), .cin(t_3084), .o(t_3130), .co(t_3131), .cout(t_3132));
compressor_4_2 u2_1072(.a(s_127_63), .b(s_127_62), .c(s_127_61), .d(s_127_60), .cin(t_3087), .o(t_3133), .co(t_3134), .cout(t_3135));
compressor_4_2 u2_1073(.a(s_128_3), .b(s_128_2), .c(s_128_1), .d(s_128_0), .cin(t_3090), .o(t_3136), .co(t_3137), .cout(t_3138));
compressor_4_2 u2_1074(.a(s_128_7), .b(s_128_6), .c(s_128_5), .d(s_128_4), .cin(t_3093), .o(t_3139), .co(t_3140), .cout(t_3141));
compressor_4_2 u2_1075(.a(s_128_11), .b(s_128_10), .c(s_128_9), .d(s_128_8), .cin(t_3096), .o(t_3142), .co(t_3143), .cout(t_3144));
compressor_4_2 u2_1076(.a(s_128_15), .b(s_128_14), .c(s_128_13), .d(s_128_12), .cin(t_3099), .o(t_3145), .co(t_3146), .cout(t_3147));
compressor_4_2 u2_1077(.a(s_128_19), .b(s_128_18), .c(s_128_17), .d(s_128_16), .cin(t_3102), .o(t_3148), .co(t_3149), .cout(t_3150));
compressor_4_2 u2_1078(.a(s_128_23), .b(s_128_22), .c(s_128_21), .d(s_128_20), .cin(t_3105), .o(t_3151), .co(t_3152), .cout(t_3153));
compressor_4_2 u2_1079(.a(s_128_27), .b(s_128_26), .c(s_128_25), .d(s_128_24), .cin(t_3108), .o(t_3154), .co(t_3155), .cout(t_3156));
compressor_4_2 u2_1080(.a(s_128_31), .b(s_128_30), .c(s_128_29), .d(s_128_28), .cin(t_3111), .o(t_3157), .co(t_3158), .cout(t_3159));
compressor_4_2 u2_1081(.a(s_128_35), .b(s_128_34), .c(s_128_33), .d(s_128_32), .cin(t_3114), .o(t_3160), .co(t_3161), .cout(t_3162));
compressor_4_2 u2_1082(.a(s_128_39), .b(s_128_38), .c(s_128_37), .d(s_128_36), .cin(t_3117), .o(t_3163), .co(t_3164), .cout(t_3165));
compressor_4_2 u2_1083(.a(s_128_43), .b(s_128_42), .c(s_128_41), .d(s_128_40), .cin(t_3120), .o(t_3166), .co(t_3167), .cout(t_3168));
compressor_4_2 u2_1084(.a(s_128_47), .b(s_128_46), .c(s_128_45), .d(s_128_44), .cin(t_3123), .o(t_3169), .co(t_3170), .cout(t_3171));
compressor_4_2 u2_1085(.a(s_128_51), .b(s_128_50), .c(s_128_49), .d(s_128_48), .cin(t_3126), .o(t_3172), .co(t_3173), .cout(t_3174));
compressor_4_2 u2_1086(.a(s_128_55), .b(s_128_54), .c(s_128_53), .d(s_128_52), .cin(t_3129), .o(t_3175), .co(t_3176), .cout(t_3177));
compressor_4_2 u2_1087(.a(s_128_59), .b(s_128_58), .c(s_128_57), .d(s_128_56), .cin(t_3132), .o(t_3178), .co(t_3179), .cout(t_3180));
compressor_4_2 u2_1088(.a(s_128_63), .b(s_128_62), .c(s_128_61), .d(s_128_60), .cin(t_3135), .o(t_3181), .co(t_3182), .cout(t_3183));
compressor_4_2 u2_1089(.a(s_129_3), .b(s_129_2), .c(s_129_1), .d(s_129_0), .cin(t_3138), .o(t_3184), .co(t_3185), .cout(t_3186));
compressor_4_2 u2_1090(.a(s_129_7), .b(s_129_6), .c(s_129_5), .d(s_129_4), .cin(t_3141), .o(t_3187), .co(t_3188), .cout(t_3189));
compressor_4_2 u2_1091(.a(s_129_11), .b(s_129_10), .c(s_129_9), .d(s_129_8), .cin(t_3144), .o(t_3190), .co(t_3191), .cout(t_3192));
compressor_4_2 u2_1092(.a(s_129_15), .b(s_129_14), .c(s_129_13), .d(s_129_12), .cin(t_3147), .o(t_3193), .co(t_3194), .cout(t_3195));
compressor_4_2 u2_1093(.a(s_129_19), .b(s_129_18), .c(s_129_17), .d(s_129_16), .cin(t_3150), .o(t_3196), .co(t_3197), .cout(t_3198));
compressor_4_2 u2_1094(.a(s_129_23), .b(s_129_22), .c(s_129_21), .d(s_129_20), .cin(t_3153), .o(t_3199), .co(t_3200), .cout(t_3201));
compressor_4_2 u2_1095(.a(s_129_27), .b(s_129_26), .c(s_129_25), .d(s_129_24), .cin(t_3156), .o(t_3202), .co(t_3203), .cout(t_3204));
compressor_4_2 u2_1096(.a(s_129_31), .b(s_129_30), .c(s_129_29), .d(s_129_28), .cin(t_3159), .o(t_3205), .co(t_3206), .cout(t_3207));
compressor_4_2 u2_1097(.a(s_129_35), .b(s_129_34), .c(s_129_33), .d(s_129_32), .cin(t_3162), .o(t_3208), .co(t_3209), .cout(t_3210));
compressor_4_2 u2_1098(.a(s_129_39), .b(s_129_38), .c(s_129_37), .d(s_129_36), .cin(t_3165), .o(t_3211), .co(t_3212), .cout(t_3213));
compressor_4_2 u2_1099(.a(s_129_43), .b(s_129_42), .c(s_129_41), .d(s_129_40), .cin(t_3168), .o(t_3214), .co(t_3215), .cout(t_3216));
compressor_4_2 u2_1100(.a(s_129_47), .b(s_129_46), .c(s_129_45), .d(s_129_44), .cin(t_3171), .o(t_3217), .co(t_3218), .cout(t_3219));
compressor_4_2 u2_1101(.a(s_129_51), .b(s_129_50), .c(s_129_49), .d(s_129_48), .cin(t_3174), .o(t_3220), .co(t_3221), .cout(t_3222));
compressor_4_2 u2_1102(.a(s_129_55), .b(s_129_54), .c(s_129_53), .d(s_129_52), .cin(t_3177), .o(t_3223), .co(t_3224), .cout(t_3225));
compressor_4_2 u2_1103(.a(s_129_59), .b(s_129_58), .c(s_129_57), .d(s_129_56), .cin(t_3180), .o(t_3226), .co(t_3227), .cout(t_3228));
compressor_4_2 u2_1104(.a(s_129_63), .b(s_129_62), .c(s_129_61), .d(s_129_60), .cin(t_3183), .o(t_3229), .co(t_3230), .cout(t_3231));
compressor_4_2 u2_1105(.a(s_130_3), .b(s_130_2), .c(s_130_1), .d(s_130_0), .cin(t_3186), .o(t_3232), .co(t_3233), .cout(t_3234));
compressor_4_2 u2_1106(.a(s_130_7), .b(s_130_6), .c(s_130_5), .d(s_130_4), .cin(t_3189), .o(t_3235), .co(t_3236), .cout(t_3237));
compressor_4_2 u2_1107(.a(s_130_11), .b(s_130_10), .c(s_130_9), .d(s_130_8), .cin(t_3192), .o(t_3238), .co(t_3239), .cout(t_3240));
compressor_4_2 u2_1108(.a(s_130_15), .b(s_130_14), .c(s_130_13), .d(s_130_12), .cin(t_3195), .o(t_3241), .co(t_3242), .cout(t_3243));
compressor_4_2 u2_1109(.a(s_130_19), .b(s_130_18), .c(s_130_17), .d(s_130_16), .cin(t_3198), .o(t_3244), .co(t_3245), .cout(t_3246));
compressor_4_2 u2_1110(.a(s_130_23), .b(s_130_22), .c(s_130_21), .d(s_130_20), .cin(t_3201), .o(t_3247), .co(t_3248), .cout(t_3249));
compressor_4_2 u2_1111(.a(s_130_27), .b(s_130_26), .c(s_130_25), .d(s_130_24), .cin(t_3204), .o(t_3250), .co(t_3251), .cout(t_3252));
compressor_4_2 u2_1112(.a(s_130_31), .b(s_130_30), .c(s_130_29), .d(s_130_28), .cin(t_3207), .o(t_3253), .co(t_3254), .cout(t_3255));
compressor_4_2 u2_1113(.a(s_130_35), .b(s_130_34), .c(s_130_33), .d(s_130_32), .cin(t_3210), .o(t_3256), .co(t_3257), .cout(t_3258));
compressor_4_2 u2_1114(.a(s_130_39), .b(s_130_38), .c(s_130_37), .d(s_130_36), .cin(t_3213), .o(t_3259), .co(t_3260), .cout(t_3261));
compressor_4_2 u2_1115(.a(s_130_43), .b(s_130_42), .c(s_130_41), .d(s_130_40), .cin(t_3216), .o(t_3262), .co(t_3263), .cout(t_3264));
compressor_4_2 u2_1116(.a(s_130_47), .b(s_130_46), .c(s_130_45), .d(s_130_44), .cin(t_3219), .o(t_3265), .co(t_3266), .cout(t_3267));
compressor_4_2 u2_1117(.a(s_130_51), .b(s_130_50), .c(s_130_49), .d(s_130_48), .cin(t_3222), .o(t_3268), .co(t_3269), .cout(t_3270));
compressor_4_2 u2_1118(.a(s_130_55), .b(s_130_54), .c(s_130_53), .d(s_130_52), .cin(t_3225), .o(t_3271), .co(t_3272), .cout(t_3273));
compressor_4_2 u2_1119(.a(s_130_59), .b(s_130_58), .c(s_130_57), .d(s_130_56), .cin(t_3228), .o(t_3274), .co(t_3275), .cout(t_3276));
compressor_4_2 u2_1120(.a(s_130_63), .b(s_130_62), .c(s_130_61), .d(s_130_60), .cin(t_3231), .o(t_3277), .co(t_3278), .cout(t_3279));
compressor_4_2 u2_1121(.a(s_131_3), .b(s_131_2), .c(s_131_1), .d(s_131_0), .cin(t_3234), .o(t_3280), .co(t_3281), .cout(t_3282));
compressor_4_2 u2_1122(.a(s_131_7), .b(s_131_6), .c(s_131_5), .d(s_131_4), .cin(t_3237), .o(t_3283), .co(t_3284), .cout(t_3285));
compressor_4_2 u2_1123(.a(s_131_11), .b(s_131_10), .c(s_131_9), .d(s_131_8), .cin(t_3240), .o(t_3286), .co(t_3287), .cout(t_3288));
compressor_4_2 u2_1124(.a(s_131_15), .b(s_131_14), .c(s_131_13), .d(s_131_12), .cin(t_3243), .o(t_3289), .co(t_3290), .cout(t_3291));
compressor_4_2 u2_1125(.a(s_131_19), .b(s_131_18), .c(s_131_17), .d(s_131_16), .cin(t_3246), .o(t_3292), .co(t_3293), .cout(t_3294));
compressor_4_2 u2_1126(.a(s_131_23), .b(s_131_22), .c(s_131_21), .d(s_131_20), .cin(t_3249), .o(t_3295), .co(t_3296), .cout(t_3297));
compressor_4_2 u2_1127(.a(s_131_27), .b(s_131_26), .c(s_131_25), .d(s_131_24), .cin(t_3252), .o(t_3298), .co(t_3299), .cout(t_3300));
compressor_4_2 u2_1128(.a(s_131_31), .b(s_131_30), .c(s_131_29), .d(s_131_28), .cin(t_3255), .o(t_3301), .co(t_3302), .cout(t_3303));
compressor_4_2 u2_1129(.a(s_131_35), .b(s_131_34), .c(s_131_33), .d(s_131_32), .cin(t_3258), .o(t_3304), .co(t_3305), .cout(t_3306));
compressor_4_2 u2_1130(.a(s_131_39), .b(s_131_38), .c(s_131_37), .d(s_131_36), .cin(t_3261), .o(t_3307), .co(t_3308), .cout(t_3309));
compressor_4_2 u2_1131(.a(s_131_43), .b(s_131_42), .c(s_131_41), .d(s_131_40), .cin(t_3264), .o(t_3310), .co(t_3311), .cout(t_3312));
compressor_4_2 u2_1132(.a(s_131_47), .b(s_131_46), .c(s_131_45), .d(s_131_44), .cin(t_3267), .o(t_3313), .co(t_3314), .cout(t_3315));
compressor_4_2 u2_1133(.a(s_131_51), .b(s_131_50), .c(s_131_49), .d(s_131_48), .cin(t_3270), .o(t_3316), .co(t_3317), .cout(t_3318));
compressor_4_2 u2_1134(.a(s_131_55), .b(s_131_54), .c(s_131_53), .d(s_131_52), .cin(t_3273), .o(t_3319), .co(t_3320), .cout(t_3321));
compressor_4_2 u2_1135(.a(s_131_59), .b(s_131_58), .c(s_131_57), .d(s_131_56), .cin(t_3276), .o(t_3322), .co(t_3323), .cout(t_3324));
compressor_4_2 u2_1136(.a(s_131_63), .b(s_131_62), .c(s_131_61), .d(s_131_60), .cin(t_3279), .o(t_3325), .co(t_3326), .cout(t_3327));
compressor_4_2 u2_1137(.a(s_132_3), .b(s_132_2), .c(s_132_1), .d(s_132_0), .cin(t_3282), .o(t_3328), .co(t_3329), .cout(t_3330));
compressor_4_2 u2_1138(.a(s_132_7), .b(s_132_6), .c(s_132_5), .d(s_132_4), .cin(t_3285), .o(t_3331), .co(t_3332), .cout(t_3333));
compressor_4_2 u2_1139(.a(s_132_11), .b(s_132_10), .c(s_132_9), .d(s_132_8), .cin(t_3288), .o(t_3334), .co(t_3335), .cout(t_3336));
compressor_4_2 u2_1140(.a(s_132_15), .b(s_132_14), .c(s_132_13), .d(s_132_12), .cin(t_3291), .o(t_3337), .co(t_3338), .cout(t_3339));
compressor_4_2 u2_1141(.a(s_132_19), .b(s_132_18), .c(s_132_17), .d(s_132_16), .cin(t_3294), .o(t_3340), .co(t_3341), .cout(t_3342));
compressor_4_2 u2_1142(.a(s_132_23), .b(s_132_22), .c(s_132_21), .d(s_132_20), .cin(t_3297), .o(t_3343), .co(t_3344), .cout(t_3345));
compressor_4_2 u2_1143(.a(s_132_27), .b(s_132_26), .c(s_132_25), .d(s_132_24), .cin(t_3300), .o(t_3346), .co(t_3347), .cout(t_3348));
compressor_4_2 u2_1144(.a(s_132_31), .b(s_132_30), .c(s_132_29), .d(s_132_28), .cin(t_3303), .o(t_3349), .co(t_3350), .cout(t_3351));
compressor_4_2 u2_1145(.a(s_132_35), .b(s_132_34), .c(s_132_33), .d(s_132_32), .cin(t_3306), .o(t_3352), .co(t_3353), .cout(t_3354));
compressor_4_2 u2_1146(.a(s_132_39), .b(s_132_38), .c(s_132_37), .d(s_132_36), .cin(t_3309), .o(t_3355), .co(t_3356), .cout(t_3357));
compressor_4_2 u2_1147(.a(s_132_43), .b(s_132_42), .c(s_132_41), .d(s_132_40), .cin(t_3312), .o(t_3358), .co(t_3359), .cout(t_3360));
compressor_4_2 u2_1148(.a(s_132_47), .b(s_132_46), .c(s_132_45), .d(s_132_44), .cin(t_3315), .o(t_3361), .co(t_3362), .cout(t_3363));
compressor_4_2 u2_1149(.a(s_132_51), .b(s_132_50), .c(s_132_49), .d(s_132_48), .cin(t_3318), .o(t_3364), .co(t_3365), .cout(t_3366));
compressor_4_2 u2_1150(.a(s_132_55), .b(s_132_54), .c(s_132_53), .d(s_132_52), .cin(t_3321), .o(t_3367), .co(t_3368), .cout(t_3369));
compressor_4_2 u2_1151(.a(s_132_59), .b(s_132_58), .c(s_132_57), .d(s_132_56), .cin(t_3324), .o(t_3370), .co(t_3371), .cout(t_3372));
compressor_3_2 u1_1152(.a(s_132_61), .b(s_132_60), .cin(t_3327), .o(t_3373), .cout(t_3374));
compressor_4_2 u2_1153(.a(s_133_3), .b(s_133_2), .c(s_133_1), .d(s_133_0), .cin(t_3330), .o(t_3375), .co(t_3376), .cout(t_3377));
compressor_4_2 u2_1154(.a(s_133_7), .b(s_133_6), .c(s_133_5), .d(s_133_4), .cin(t_3333), .o(t_3378), .co(t_3379), .cout(t_3380));
compressor_4_2 u2_1155(.a(s_133_11), .b(s_133_10), .c(s_133_9), .d(s_133_8), .cin(t_3336), .o(t_3381), .co(t_3382), .cout(t_3383));
compressor_4_2 u2_1156(.a(s_133_15), .b(s_133_14), .c(s_133_13), .d(s_133_12), .cin(t_3339), .o(t_3384), .co(t_3385), .cout(t_3386));
compressor_4_2 u2_1157(.a(s_133_19), .b(s_133_18), .c(s_133_17), .d(s_133_16), .cin(t_3342), .o(t_3387), .co(t_3388), .cout(t_3389));
compressor_4_2 u2_1158(.a(s_133_23), .b(s_133_22), .c(s_133_21), .d(s_133_20), .cin(t_3345), .o(t_3390), .co(t_3391), .cout(t_3392));
compressor_4_2 u2_1159(.a(s_133_27), .b(s_133_26), .c(s_133_25), .d(s_133_24), .cin(t_3348), .o(t_3393), .co(t_3394), .cout(t_3395));
compressor_4_2 u2_1160(.a(s_133_31), .b(s_133_30), .c(s_133_29), .d(s_133_28), .cin(t_3351), .o(t_3396), .co(t_3397), .cout(t_3398));
compressor_4_2 u2_1161(.a(s_133_35), .b(s_133_34), .c(s_133_33), .d(s_133_32), .cin(t_3354), .o(t_3399), .co(t_3400), .cout(t_3401));
compressor_4_2 u2_1162(.a(s_133_39), .b(s_133_38), .c(s_133_37), .d(s_133_36), .cin(t_3357), .o(t_3402), .co(t_3403), .cout(t_3404));
compressor_4_2 u2_1163(.a(s_133_43), .b(s_133_42), .c(s_133_41), .d(s_133_40), .cin(t_3360), .o(t_3405), .co(t_3406), .cout(t_3407));
compressor_4_2 u2_1164(.a(s_133_47), .b(s_133_46), .c(s_133_45), .d(s_133_44), .cin(t_3363), .o(t_3408), .co(t_3409), .cout(t_3410));
compressor_4_2 u2_1165(.a(s_133_51), .b(s_133_50), .c(s_133_49), .d(s_133_48), .cin(t_3366), .o(t_3411), .co(t_3412), .cout(t_3413));
compressor_4_2 u2_1166(.a(s_133_55), .b(s_133_54), .c(s_133_53), .d(s_133_52), .cin(t_3369), .o(t_3414), .co(t_3415), .cout(t_3416));
compressor_4_2 u2_1167(.a(s_133_59), .b(s_133_58), .c(s_133_57), .d(s_133_56), .cin(t_3372), .o(t_3417), .co(t_3418), .cout(t_3419));
compressor_3_2 u1_1168(.a(s_133_62), .b(s_133_61), .cin(s_133_60), .o(t_3420), .cout(t_3421));
compressor_4_2 u2_1169(.a(s_134_3), .b(s_134_2), .c(s_134_1), .d(s_134_0), .cin(t_3377), .o(t_3422), .co(t_3423), .cout(t_3424));
compressor_4_2 u2_1170(.a(s_134_7), .b(s_134_6), .c(s_134_5), .d(s_134_4), .cin(t_3380), .o(t_3425), .co(t_3426), .cout(t_3427));
compressor_4_2 u2_1171(.a(s_134_11), .b(s_134_10), .c(s_134_9), .d(s_134_8), .cin(t_3383), .o(t_3428), .co(t_3429), .cout(t_3430));
compressor_4_2 u2_1172(.a(s_134_15), .b(s_134_14), .c(s_134_13), .d(s_134_12), .cin(t_3386), .o(t_3431), .co(t_3432), .cout(t_3433));
compressor_4_2 u2_1173(.a(s_134_19), .b(s_134_18), .c(s_134_17), .d(s_134_16), .cin(t_3389), .o(t_3434), .co(t_3435), .cout(t_3436));
compressor_4_2 u2_1174(.a(s_134_23), .b(s_134_22), .c(s_134_21), .d(s_134_20), .cin(t_3392), .o(t_3437), .co(t_3438), .cout(t_3439));
compressor_4_2 u2_1175(.a(s_134_27), .b(s_134_26), .c(s_134_25), .d(s_134_24), .cin(t_3395), .o(t_3440), .co(t_3441), .cout(t_3442));
compressor_4_2 u2_1176(.a(s_134_31), .b(s_134_30), .c(s_134_29), .d(s_134_28), .cin(t_3398), .o(t_3443), .co(t_3444), .cout(t_3445));
compressor_4_2 u2_1177(.a(s_134_35), .b(s_134_34), .c(s_134_33), .d(s_134_32), .cin(t_3401), .o(t_3446), .co(t_3447), .cout(t_3448));
compressor_4_2 u2_1178(.a(s_134_39), .b(s_134_38), .c(s_134_37), .d(s_134_36), .cin(t_3404), .o(t_3449), .co(t_3450), .cout(t_3451));
compressor_4_2 u2_1179(.a(s_134_43), .b(s_134_42), .c(s_134_41), .d(s_134_40), .cin(t_3407), .o(t_3452), .co(t_3453), .cout(t_3454));
compressor_4_2 u2_1180(.a(s_134_47), .b(s_134_46), .c(s_134_45), .d(s_134_44), .cin(t_3410), .o(t_3455), .co(t_3456), .cout(t_3457));
compressor_4_2 u2_1181(.a(s_134_51), .b(s_134_50), .c(s_134_49), .d(s_134_48), .cin(t_3413), .o(t_3458), .co(t_3459), .cout(t_3460));
compressor_4_2 u2_1182(.a(s_134_55), .b(s_134_54), .c(s_134_53), .d(s_134_52), .cin(t_3416), .o(t_3461), .co(t_3462), .cout(t_3463));
compressor_4_2 u2_1183(.a(s_134_59), .b(s_134_58), .c(s_134_57), .d(s_134_56), .cin(t_3419), .o(t_3464), .co(t_3465), .cout(t_3466));
half_adder u0_1184(.a(s_134_61), .b(s_134_60), .o(t_3467), .cout(t_3468));
compressor_4_2 u2_1185(.a(s_135_3), .b(s_135_2), .c(s_135_1), .d(s_135_0), .cin(t_3424), .o(t_3469), .co(t_3470), .cout(t_3471));
compressor_4_2 u2_1186(.a(s_135_7), .b(s_135_6), .c(s_135_5), .d(s_135_4), .cin(t_3427), .o(t_3472), .co(t_3473), .cout(t_3474));
compressor_4_2 u2_1187(.a(s_135_11), .b(s_135_10), .c(s_135_9), .d(s_135_8), .cin(t_3430), .o(t_3475), .co(t_3476), .cout(t_3477));
compressor_4_2 u2_1188(.a(s_135_15), .b(s_135_14), .c(s_135_13), .d(s_135_12), .cin(t_3433), .o(t_3478), .co(t_3479), .cout(t_3480));
compressor_4_2 u2_1189(.a(s_135_19), .b(s_135_18), .c(s_135_17), .d(s_135_16), .cin(t_3436), .o(t_3481), .co(t_3482), .cout(t_3483));
compressor_4_2 u2_1190(.a(s_135_23), .b(s_135_22), .c(s_135_21), .d(s_135_20), .cin(t_3439), .o(t_3484), .co(t_3485), .cout(t_3486));
compressor_4_2 u2_1191(.a(s_135_27), .b(s_135_26), .c(s_135_25), .d(s_135_24), .cin(t_3442), .o(t_3487), .co(t_3488), .cout(t_3489));
compressor_4_2 u2_1192(.a(s_135_31), .b(s_135_30), .c(s_135_29), .d(s_135_28), .cin(t_3445), .o(t_3490), .co(t_3491), .cout(t_3492));
compressor_4_2 u2_1193(.a(s_135_35), .b(s_135_34), .c(s_135_33), .d(s_135_32), .cin(t_3448), .o(t_3493), .co(t_3494), .cout(t_3495));
compressor_4_2 u2_1194(.a(s_135_39), .b(s_135_38), .c(s_135_37), .d(s_135_36), .cin(t_3451), .o(t_3496), .co(t_3497), .cout(t_3498));
compressor_4_2 u2_1195(.a(s_135_43), .b(s_135_42), .c(s_135_41), .d(s_135_40), .cin(t_3454), .o(t_3499), .co(t_3500), .cout(t_3501));
compressor_4_2 u2_1196(.a(s_135_47), .b(s_135_46), .c(s_135_45), .d(s_135_44), .cin(t_3457), .o(t_3502), .co(t_3503), .cout(t_3504));
compressor_4_2 u2_1197(.a(s_135_51), .b(s_135_50), .c(s_135_49), .d(s_135_48), .cin(t_3460), .o(t_3505), .co(t_3506), .cout(t_3507));
compressor_4_2 u2_1198(.a(s_135_55), .b(s_135_54), .c(s_135_53), .d(s_135_52), .cin(t_3463), .o(t_3508), .co(t_3509), .cout(t_3510));
compressor_4_2 u2_1199(.a(s_135_59), .b(s_135_58), .c(s_135_57), .d(s_135_56), .cin(t_3466), .o(t_3511), .co(t_3512), .cout(t_3513));
half_adder u0_1200(.a(s_135_61), .b(s_135_60), .o(t_3514), .cout(t_3515));
compressor_4_2 u2_1201(.a(s_136_3), .b(s_136_2), .c(s_136_1), .d(s_136_0), .cin(t_3471), .o(t_3516), .co(t_3517), .cout(t_3518));
compressor_4_2 u2_1202(.a(s_136_7), .b(s_136_6), .c(s_136_5), .d(s_136_4), .cin(t_3474), .o(t_3519), .co(t_3520), .cout(t_3521));
compressor_4_2 u2_1203(.a(s_136_11), .b(s_136_10), .c(s_136_9), .d(s_136_8), .cin(t_3477), .o(t_3522), .co(t_3523), .cout(t_3524));
compressor_4_2 u2_1204(.a(s_136_15), .b(s_136_14), .c(s_136_13), .d(s_136_12), .cin(t_3480), .o(t_3525), .co(t_3526), .cout(t_3527));
compressor_4_2 u2_1205(.a(s_136_19), .b(s_136_18), .c(s_136_17), .d(s_136_16), .cin(t_3483), .o(t_3528), .co(t_3529), .cout(t_3530));
compressor_4_2 u2_1206(.a(s_136_23), .b(s_136_22), .c(s_136_21), .d(s_136_20), .cin(t_3486), .o(t_3531), .co(t_3532), .cout(t_3533));
compressor_4_2 u2_1207(.a(s_136_27), .b(s_136_26), .c(s_136_25), .d(s_136_24), .cin(t_3489), .o(t_3534), .co(t_3535), .cout(t_3536));
compressor_4_2 u2_1208(.a(s_136_31), .b(s_136_30), .c(s_136_29), .d(s_136_28), .cin(t_3492), .o(t_3537), .co(t_3538), .cout(t_3539));
compressor_4_2 u2_1209(.a(s_136_35), .b(s_136_34), .c(s_136_33), .d(s_136_32), .cin(t_3495), .o(t_3540), .co(t_3541), .cout(t_3542));
compressor_4_2 u2_1210(.a(s_136_39), .b(s_136_38), .c(s_136_37), .d(s_136_36), .cin(t_3498), .o(t_3543), .co(t_3544), .cout(t_3545));
compressor_4_2 u2_1211(.a(s_136_43), .b(s_136_42), .c(s_136_41), .d(s_136_40), .cin(t_3501), .o(t_3546), .co(t_3547), .cout(t_3548));
compressor_4_2 u2_1212(.a(s_136_47), .b(s_136_46), .c(s_136_45), .d(s_136_44), .cin(t_3504), .o(t_3549), .co(t_3550), .cout(t_3551));
compressor_4_2 u2_1213(.a(s_136_51), .b(s_136_50), .c(s_136_49), .d(s_136_48), .cin(t_3507), .o(t_3552), .co(t_3553), .cout(t_3554));
compressor_4_2 u2_1214(.a(s_136_55), .b(s_136_54), .c(s_136_53), .d(s_136_52), .cin(t_3510), .o(t_3555), .co(t_3556), .cout(t_3557));
compressor_4_2 u2_1215(.a(s_136_59), .b(s_136_58), .c(s_136_57), .d(s_136_56), .cin(t_3513), .o(t_3558), .co(t_3559), .cout(t_3560));
compressor_4_2 u2_1216(.a(s_137_3), .b(s_137_2), .c(s_137_1), .d(s_137_0), .cin(t_3518), .o(t_3561), .co(t_3562), .cout(t_3563));
compressor_4_2 u2_1217(.a(s_137_7), .b(s_137_6), .c(s_137_5), .d(s_137_4), .cin(t_3521), .o(t_3564), .co(t_3565), .cout(t_3566));
compressor_4_2 u2_1218(.a(s_137_11), .b(s_137_10), .c(s_137_9), .d(s_137_8), .cin(t_3524), .o(t_3567), .co(t_3568), .cout(t_3569));
compressor_4_2 u2_1219(.a(s_137_15), .b(s_137_14), .c(s_137_13), .d(s_137_12), .cin(t_3527), .o(t_3570), .co(t_3571), .cout(t_3572));
compressor_4_2 u2_1220(.a(s_137_19), .b(s_137_18), .c(s_137_17), .d(s_137_16), .cin(t_3530), .o(t_3573), .co(t_3574), .cout(t_3575));
compressor_4_2 u2_1221(.a(s_137_23), .b(s_137_22), .c(s_137_21), .d(s_137_20), .cin(t_3533), .o(t_3576), .co(t_3577), .cout(t_3578));
compressor_4_2 u2_1222(.a(s_137_27), .b(s_137_26), .c(s_137_25), .d(s_137_24), .cin(t_3536), .o(t_3579), .co(t_3580), .cout(t_3581));
compressor_4_2 u2_1223(.a(s_137_31), .b(s_137_30), .c(s_137_29), .d(s_137_28), .cin(t_3539), .o(t_3582), .co(t_3583), .cout(t_3584));
compressor_4_2 u2_1224(.a(s_137_35), .b(s_137_34), .c(s_137_33), .d(s_137_32), .cin(t_3542), .o(t_3585), .co(t_3586), .cout(t_3587));
compressor_4_2 u2_1225(.a(s_137_39), .b(s_137_38), .c(s_137_37), .d(s_137_36), .cin(t_3545), .o(t_3588), .co(t_3589), .cout(t_3590));
compressor_4_2 u2_1226(.a(s_137_43), .b(s_137_42), .c(s_137_41), .d(s_137_40), .cin(t_3548), .o(t_3591), .co(t_3592), .cout(t_3593));
compressor_4_2 u2_1227(.a(s_137_47), .b(s_137_46), .c(s_137_45), .d(s_137_44), .cin(t_3551), .o(t_3594), .co(t_3595), .cout(t_3596));
compressor_4_2 u2_1228(.a(s_137_51), .b(s_137_50), .c(s_137_49), .d(s_137_48), .cin(t_3554), .o(t_3597), .co(t_3598), .cout(t_3599));
compressor_4_2 u2_1229(.a(s_137_55), .b(s_137_54), .c(s_137_53), .d(s_137_52), .cin(t_3557), .o(t_3600), .co(t_3601), .cout(t_3602));
compressor_4_2 u2_1230(.a(s_137_59), .b(s_137_58), .c(s_137_57), .d(s_137_56), .cin(t_3560), .o(t_3603), .co(t_3604), .cout(t_3605));
compressor_4_2 u2_1231(.a(s_138_3), .b(s_138_2), .c(s_138_1), .d(s_138_0), .cin(t_3563), .o(t_3606), .co(t_3607), .cout(t_3608));
compressor_4_2 u2_1232(.a(s_138_7), .b(s_138_6), .c(s_138_5), .d(s_138_4), .cin(t_3566), .o(t_3609), .co(t_3610), .cout(t_3611));
compressor_4_2 u2_1233(.a(s_138_11), .b(s_138_10), .c(s_138_9), .d(s_138_8), .cin(t_3569), .o(t_3612), .co(t_3613), .cout(t_3614));
compressor_4_2 u2_1234(.a(s_138_15), .b(s_138_14), .c(s_138_13), .d(s_138_12), .cin(t_3572), .o(t_3615), .co(t_3616), .cout(t_3617));
compressor_4_2 u2_1235(.a(s_138_19), .b(s_138_18), .c(s_138_17), .d(s_138_16), .cin(t_3575), .o(t_3618), .co(t_3619), .cout(t_3620));
compressor_4_2 u2_1236(.a(s_138_23), .b(s_138_22), .c(s_138_21), .d(s_138_20), .cin(t_3578), .o(t_3621), .co(t_3622), .cout(t_3623));
compressor_4_2 u2_1237(.a(s_138_27), .b(s_138_26), .c(s_138_25), .d(s_138_24), .cin(t_3581), .o(t_3624), .co(t_3625), .cout(t_3626));
compressor_4_2 u2_1238(.a(s_138_31), .b(s_138_30), .c(s_138_29), .d(s_138_28), .cin(t_3584), .o(t_3627), .co(t_3628), .cout(t_3629));
compressor_4_2 u2_1239(.a(s_138_35), .b(s_138_34), .c(s_138_33), .d(s_138_32), .cin(t_3587), .o(t_3630), .co(t_3631), .cout(t_3632));
compressor_4_2 u2_1240(.a(s_138_39), .b(s_138_38), .c(s_138_37), .d(s_138_36), .cin(t_3590), .o(t_3633), .co(t_3634), .cout(t_3635));
compressor_4_2 u2_1241(.a(s_138_43), .b(s_138_42), .c(s_138_41), .d(s_138_40), .cin(t_3593), .o(t_3636), .co(t_3637), .cout(t_3638));
compressor_4_2 u2_1242(.a(s_138_47), .b(s_138_46), .c(s_138_45), .d(s_138_44), .cin(t_3596), .o(t_3639), .co(t_3640), .cout(t_3641));
compressor_4_2 u2_1243(.a(s_138_51), .b(s_138_50), .c(s_138_49), .d(s_138_48), .cin(t_3599), .o(t_3642), .co(t_3643), .cout(t_3644));
compressor_4_2 u2_1244(.a(s_138_55), .b(s_138_54), .c(s_138_53), .d(s_138_52), .cin(t_3602), .o(t_3645), .co(t_3646), .cout(t_3647));
compressor_4_2 u2_1245(.a(s_138_59), .b(s_138_58), .c(s_138_57), .d(s_138_56), .cin(t_3605), .o(t_3648), .co(t_3649), .cout(t_3650));
compressor_4_2 u2_1246(.a(s_139_3), .b(s_139_2), .c(s_139_1), .d(s_139_0), .cin(t_3608), .o(t_3651), .co(t_3652), .cout(t_3653));
compressor_4_2 u2_1247(.a(s_139_7), .b(s_139_6), .c(s_139_5), .d(s_139_4), .cin(t_3611), .o(t_3654), .co(t_3655), .cout(t_3656));
compressor_4_2 u2_1248(.a(s_139_11), .b(s_139_10), .c(s_139_9), .d(s_139_8), .cin(t_3614), .o(t_3657), .co(t_3658), .cout(t_3659));
compressor_4_2 u2_1249(.a(s_139_15), .b(s_139_14), .c(s_139_13), .d(s_139_12), .cin(t_3617), .o(t_3660), .co(t_3661), .cout(t_3662));
compressor_4_2 u2_1250(.a(s_139_19), .b(s_139_18), .c(s_139_17), .d(s_139_16), .cin(t_3620), .o(t_3663), .co(t_3664), .cout(t_3665));
compressor_4_2 u2_1251(.a(s_139_23), .b(s_139_22), .c(s_139_21), .d(s_139_20), .cin(t_3623), .o(t_3666), .co(t_3667), .cout(t_3668));
compressor_4_2 u2_1252(.a(s_139_27), .b(s_139_26), .c(s_139_25), .d(s_139_24), .cin(t_3626), .o(t_3669), .co(t_3670), .cout(t_3671));
compressor_4_2 u2_1253(.a(s_139_31), .b(s_139_30), .c(s_139_29), .d(s_139_28), .cin(t_3629), .o(t_3672), .co(t_3673), .cout(t_3674));
compressor_4_2 u2_1254(.a(s_139_35), .b(s_139_34), .c(s_139_33), .d(s_139_32), .cin(t_3632), .o(t_3675), .co(t_3676), .cout(t_3677));
compressor_4_2 u2_1255(.a(s_139_39), .b(s_139_38), .c(s_139_37), .d(s_139_36), .cin(t_3635), .o(t_3678), .co(t_3679), .cout(t_3680));
compressor_4_2 u2_1256(.a(s_139_43), .b(s_139_42), .c(s_139_41), .d(s_139_40), .cin(t_3638), .o(t_3681), .co(t_3682), .cout(t_3683));
compressor_4_2 u2_1257(.a(s_139_47), .b(s_139_46), .c(s_139_45), .d(s_139_44), .cin(t_3641), .o(t_3684), .co(t_3685), .cout(t_3686));
compressor_4_2 u2_1258(.a(s_139_51), .b(s_139_50), .c(s_139_49), .d(s_139_48), .cin(t_3644), .o(t_3687), .co(t_3688), .cout(t_3689));
compressor_4_2 u2_1259(.a(s_139_55), .b(s_139_54), .c(s_139_53), .d(s_139_52), .cin(t_3647), .o(t_3690), .co(t_3691), .cout(t_3692));
compressor_4_2 u2_1260(.a(s_139_59), .b(s_139_58), .c(s_139_57), .d(s_139_56), .cin(t_3650), .o(t_3693), .co(t_3694), .cout(t_3695));
compressor_4_2 u2_1261(.a(s_140_3), .b(s_140_2), .c(s_140_1), .d(s_140_0), .cin(t_3653), .o(t_3696), .co(t_3697), .cout(t_3698));
compressor_4_2 u2_1262(.a(s_140_7), .b(s_140_6), .c(s_140_5), .d(s_140_4), .cin(t_3656), .o(t_3699), .co(t_3700), .cout(t_3701));
compressor_4_2 u2_1263(.a(s_140_11), .b(s_140_10), .c(s_140_9), .d(s_140_8), .cin(t_3659), .o(t_3702), .co(t_3703), .cout(t_3704));
compressor_4_2 u2_1264(.a(s_140_15), .b(s_140_14), .c(s_140_13), .d(s_140_12), .cin(t_3662), .o(t_3705), .co(t_3706), .cout(t_3707));
compressor_4_2 u2_1265(.a(s_140_19), .b(s_140_18), .c(s_140_17), .d(s_140_16), .cin(t_3665), .o(t_3708), .co(t_3709), .cout(t_3710));
compressor_4_2 u2_1266(.a(s_140_23), .b(s_140_22), .c(s_140_21), .d(s_140_20), .cin(t_3668), .o(t_3711), .co(t_3712), .cout(t_3713));
compressor_4_2 u2_1267(.a(s_140_27), .b(s_140_26), .c(s_140_25), .d(s_140_24), .cin(t_3671), .o(t_3714), .co(t_3715), .cout(t_3716));
compressor_4_2 u2_1268(.a(s_140_31), .b(s_140_30), .c(s_140_29), .d(s_140_28), .cin(t_3674), .o(t_3717), .co(t_3718), .cout(t_3719));
compressor_4_2 u2_1269(.a(s_140_35), .b(s_140_34), .c(s_140_33), .d(s_140_32), .cin(t_3677), .o(t_3720), .co(t_3721), .cout(t_3722));
compressor_4_2 u2_1270(.a(s_140_39), .b(s_140_38), .c(s_140_37), .d(s_140_36), .cin(t_3680), .o(t_3723), .co(t_3724), .cout(t_3725));
compressor_4_2 u2_1271(.a(s_140_43), .b(s_140_42), .c(s_140_41), .d(s_140_40), .cin(t_3683), .o(t_3726), .co(t_3727), .cout(t_3728));
compressor_4_2 u2_1272(.a(s_140_47), .b(s_140_46), .c(s_140_45), .d(s_140_44), .cin(t_3686), .o(t_3729), .co(t_3730), .cout(t_3731));
compressor_4_2 u2_1273(.a(s_140_51), .b(s_140_50), .c(s_140_49), .d(s_140_48), .cin(t_3689), .o(t_3732), .co(t_3733), .cout(t_3734));
compressor_4_2 u2_1274(.a(s_140_55), .b(s_140_54), .c(s_140_53), .d(s_140_52), .cin(t_3692), .o(t_3735), .co(t_3736), .cout(t_3737));
compressor_3_2 u1_1275(.a(s_140_57), .b(s_140_56), .cin(t_3695), .o(t_3738), .cout(t_3739));
compressor_4_2 u2_1276(.a(s_141_3), .b(s_141_2), .c(s_141_1), .d(s_141_0), .cin(t_3698), .o(t_3740), .co(t_3741), .cout(t_3742));
compressor_4_2 u2_1277(.a(s_141_7), .b(s_141_6), .c(s_141_5), .d(s_141_4), .cin(t_3701), .o(t_3743), .co(t_3744), .cout(t_3745));
compressor_4_2 u2_1278(.a(s_141_11), .b(s_141_10), .c(s_141_9), .d(s_141_8), .cin(t_3704), .o(t_3746), .co(t_3747), .cout(t_3748));
compressor_4_2 u2_1279(.a(s_141_15), .b(s_141_14), .c(s_141_13), .d(s_141_12), .cin(t_3707), .o(t_3749), .co(t_3750), .cout(t_3751));
compressor_4_2 u2_1280(.a(s_141_19), .b(s_141_18), .c(s_141_17), .d(s_141_16), .cin(t_3710), .o(t_3752), .co(t_3753), .cout(t_3754));
compressor_4_2 u2_1281(.a(s_141_23), .b(s_141_22), .c(s_141_21), .d(s_141_20), .cin(t_3713), .o(t_3755), .co(t_3756), .cout(t_3757));
compressor_4_2 u2_1282(.a(s_141_27), .b(s_141_26), .c(s_141_25), .d(s_141_24), .cin(t_3716), .o(t_3758), .co(t_3759), .cout(t_3760));
compressor_4_2 u2_1283(.a(s_141_31), .b(s_141_30), .c(s_141_29), .d(s_141_28), .cin(t_3719), .o(t_3761), .co(t_3762), .cout(t_3763));
compressor_4_2 u2_1284(.a(s_141_35), .b(s_141_34), .c(s_141_33), .d(s_141_32), .cin(t_3722), .o(t_3764), .co(t_3765), .cout(t_3766));
compressor_4_2 u2_1285(.a(s_141_39), .b(s_141_38), .c(s_141_37), .d(s_141_36), .cin(t_3725), .o(t_3767), .co(t_3768), .cout(t_3769));
compressor_4_2 u2_1286(.a(s_141_43), .b(s_141_42), .c(s_141_41), .d(s_141_40), .cin(t_3728), .o(t_3770), .co(t_3771), .cout(t_3772));
compressor_4_2 u2_1287(.a(s_141_47), .b(s_141_46), .c(s_141_45), .d(s_141_44), .cin(t_3731), .o(t_3773), .co(t_3774), .cout(t_3775));
compressor_4_2 u2_1288(.a(s_141_51), .b(s_141_50), .c(s_141_49), .d(s_141_48), .cin(t_3734), .o(t_3776), .co(t_3777), .cout(t_3778));
compressor_4_2 u2_1289(.a(s_141_55), .b(s_141_54), .c(s_141_53), .d(s_141_52), .cin(t_3737), .o(t_3779), .co(t_3780), .cout(t_3781));
compressor_3_2 u1_1290(.a(s_141_58), .b(s_141_57), .cin(s_141_56), .o(t_3782), .cout(t_3783));
compressor_4_2 u2_1291(.a(s_142_3), .b(s_142_2), .c(s_142_1), .d(s_142_0), .cin(t_3742), .o(t_3784), .co(t_3785), .cout(t_3786));
compressor_4_2 u2_1292(.a(s_142_7), .b(s_142_6), .c(s_142_5), .d(s_142_4), .cin(t_3745), .o(t_3787), .co(t_3788), .cout(t_3789));
compressor_4_2 u2_1293(.a(s_142_11), .b(s_142_10), .c(s_142_9), .d(s_142_8), .cin(t_3748), .o(t_3790), .co(t_3791), .cout(t_3792));
compressor_4_2 u2_1294(.a(s_142_15), .b(s_142_14), .c(s_142_13), .d(s_142_12), .cin(t_3751), .o(t_3793), .co(t_3794), .cout(t_3795));
compressor_4_2 u2_1295(.a(s_142_19), .b(s_142_18), .c(s_142_17), .d(s_142_16), .cin(t_3754), .o(t_3796), .co(t_3797), .cout(t_3798));
compressor_4_2 u2_1296(.a(s_142_23), .b(s_142_22), .c(s_142_21), .d(s_142_20), .cin(t_3757), .o(t_3799), .co(t_3800), .cout(t_3801));
compressor_4_2 u2_1297(.a(s_142_27), .b(s_142_26), .c(s_142_25), .d(s_142_24), .cin(t_3760), .o(t_3802), .co(t_3803), .cout(t_3804));
compressor_4_2 u2_1298(.a(s_142_31), .b(s_142_30), .c(s_142_29), .d(s_142_28), .cin(t_3763), .o(t_3805), .co(t_3806), .cout(t_3807));
compressor_4_2 u2_1299(.a(s_142_35), .b(s_142_34), .c(s_142_33), .d(s_142_32), .cin(t_3766), .o(t_3808), .co(t_3809), .cout(t_3810));
compressor_4_2 u2_1300(.a(s_142_39), .b(s_142_38), .c(s_142_37), .d(s_142_36), .cin(t_3769), .o(t_3811), .co(t_3812), .cout(t_3813));
compressor_4_2 u2_1301(.a(s_142_43), .b(s_142_42), .c(s_142_41), .d(s_142_40), .cin(t_3772), .o(t_3814), .co(t_3815), .cout(t_3816));
compressor_4_2 u2_1302(.a(s_142_47), .b(s_142_46), .c(s_142_45), .d(s_142_44), .cin(t_3775), .o(t_3817), .co(t_3818), .cout(t_3819));
compressor_4_2 u2_1303(.a(s_142_51), .b(s_142_50), .c(s_142_49), .d(s_142_48), .cin(t_3778), .o(t_3820), .co(t_3821), .cout(t_3822));
compressor_4_2 u2_1304(.a(s_142_55), .b(s_142_54), .c(s_142_53), .d(s_142_52), .cin(t_3781), .o(t_3823), .co(t_3824), .cout(t_3825));
half_adder u0_1305(.a(s_142_57), .b(s_142_56), .o(t_3826), .cout(t_3827));
compressor_4_2 u2_1306(.a(s_143_3), .b(s_143_2), .c(s_143_1), .d(s_143_0), .cin(t_3786), .o(t_3828), .co(t_3829), .cout(t_3830));
compressor_4_2 u2_1307(.a(s_143_7), .b(s_143_6), .c(s_143_5), .d(s_143_4), .cin(t_3789), .o(t_3831), .co(t_3832), .cout(t_3833));
compressor_4_2 u2_1308(.a(s_143_11), .b(s_143_10), .c(s_143_9), .d(s_143_8), .cin(t_3792), .o(t_3834), .co(t_3835), .cout(t_3836));
compressor_4_2 u2_1309(.a(s_143_15), .b(s_143_14), .c(s_143_13), .d(s_143_12), .cin(t_3795), .o(t_3837), .co(t_3838), .cout(t_3839));
compressor_4_2 u2_1310(.a(s_143_19), .b(s_143_18), .c(s_143_17), .d(s_143_16), .cin(t_3798), .o(t_3840), .co(t_3841), .cout(t_3842));
compressor_4_2 u2_1311(.a(s_143_23), .b(s_143_22), .c(s_143_21), .d(s_143_20), .cin(t_3801), .o(t_3843), .co(t_3844), .cout(t_3845));
compressor_4_2 u2_1312(.a(s_143_27), .b(s_143_26), .c(s_143_25), .d(s_143_24), .cin(t_3804), .o(t_3846), .co(t_3847), .cout(t_3848));
compressor_4_2 u2_1313(.a(s_143_31), .b(s_143_30), .c(s_143_29), .d(s_143_28), .cin(t_3807), .o(t_3849), .co(t_3850), .cout(t_3851));
compressor_4_2 u2_1314(.a(s_143_35), .b(s_143_34), .c(s_143_33), .d(s_143_32), .cin(t_3810), .o(t_3852), .co(t_3853), .cout(t_3854));
compressor_4_2 u2_1315(.a(s_143_39), .b(s_143_38), .c(s_143_37), .d(s_143_36), .cin(t_3813), .o(t_3855), .co(t_3856), .cout(t_3857));
compressor_4_2 u2_1316(.a(s_143_43), .b(s_143_42), .c(s_143_41), .d(s_143_40), .cin(t_3816), .o(t_3858), .co(t_3859), .cout(t_3860));
compressor_4_2 u2_1317(.a(s_143_47), .b(s_143_46), .c(s_143_45), .d(s_143_44), .cin(t_3819), .o(t_3861), .co(t_3862), .cout(t_3863));
compressor_4_2 u2_1318(.a(s_143_51), .b(s_143_50), .c(s_143_49), .d(s_143_48), .cin(t_3822), .o(t_3864), .co(t_3865), .cout(t_3866));
compressor_4_2 u2_1319(.a(s_143_55), .b(s_143_54), .c(s_143_53), .d(s_143_52), .cin(t_3825), .o(t_3867), .co(t_3868), .cout(t_3869));
half_adder u0_1320(.a(s_143_57), .b(s_143_56), .o(t_3870), .cout(t_3871));
compressor_4_2 u2_1321(.a(s_144_3), .b(s_144_2), .c(s_144_1), .d(s_144_0), .cin(t_3830), .o(t_3872), .co(t_3873), .cout(t_3874));
compressor_4_2 u2_1322(.a(s_144_7), .b(s_144_6), .c(s_144_5), .d(s_144_4), .cin(t_3833), .o(t_3875), .co(t_3876), .cout(t_3877));
compressor_4_2 u2_1323(.a(s_144_11), .b(s_144_10), .c(s_144_9), .d(s_144_8), .cin(t_3836), .o(t_3878), .co(t_3879), .cout(t_3880));
compressor_4_2 u2_1324(.a(s_144_15), .b(s_144_14), .c(s_144_13), .d(s_144_12), .cin(t_3839), .o(t_3881), .co(t_3882), .cout(t_3883));
compressor_4_2 u2_1325(.a(s_144_19), .b(s_144_18), .c(s_144_17), .d(s_144_16), .cin(t_3842), .o(t_3884), .co(t_3885), .cout(t_3886));
compressor_4_2 u2_1326(.a(s_144_23), .b(s_144_22), .c(s_144_21), .d(s_144_20), .cin(t_3845), .o(t_3887), .co(t_3888), .cout(t_3889));
compressor_4_2 u2_1327(.a(s_144_27), .b(s_144_26), .c(s_144_25), .d(s_144_24), .cin(t_3848), .o(t_3890), .co(t_3891), .cout(t_3892));
compressor_4_2 u2_1328(.a(s_144_31), .b(s_144_30), .c(s_144_29), .d(s_144_28), .cin(t_3851), .o(t_3893), .co(t_3894), .cout(t_3895));
compressor_4_2 u2_1329(.a(s_144_35), .b(s_144_34), .c(s_144_33), .d(s_144_32), .cin(t_3854), .o(t_3896), .co(t_3897), .cout(t_3898));
compressor_4_2 u2_1330(.a(s_144_39), .b(s_144_38), .c(s_144_37), .d(s_144_36), .cin(t_3857), .o(t_3899), .co(t_3900), .cout(t_3901));
compressor_4_2 u2_1331(.a(s_144_43), .b(s_144_42), .c(s_144_41), .d(s_144_40), .cin(t_3860), .o(t_3902), .co(t_3903), .cout(t_3904));
compressor_4_2 u2_1332(.a(s_144_47), .b(s_144_46), .c(s_144_45), .d(s_144_44), .cin(t_3863), .o(t_3905), .co(t_3906), .cout(t_3907));
compressor_4_2 u2_1333(.a(s_144_51), .b(s_144_50), .c(s_144_49), .d(s_144_48), .cin(t_3866), .o(t_3908), .co(t_3909), .cout(t_3910));
compressor_4_2 u2_1334(.a(s_144_55), .b(s_144_54), .c(s_144_53), .d(s_144_52), .cin(t_3869), .o(t_3911), .co(t_3912), .cout(t_3913));
compressor_4_2 u2_1335(.a(s_145_3), .b(s_145_2), .c(s_145_1), .d(s_145_0), .cin(t_3874), .o(t_3914), .co(t_3915), .cout(t_3916));
compressor_4_2 u2_1336(.a(s_145_7), .b(s_145_6), .c(s_145_5), .d(s_145_4), .cin(t_3877), .o(t_3917), .co(t_3918), .cout(t_3919));
compressor_4_2 u2_1337(.a(s_145_11), .b(s_145_10), .c(s_145_9), .d(s_145_8), .cin(t_3880), .o(t_3920), .co(t_3921), .cout(t_3922));
compressor_4_2 u2_1338(.a(s_145_15), .b(s_145_14), .c(s_145_13), .d(s_145_12), .cin(t_3883), .o(t_3923), .co(t_3924), .cout(t_3925));
compressor_4_2 u2_1339(.a(s_145_19), .b(s_145_18), .c(s_145_17), .d(s_145_16), .cin(t_3886), .o(t_3926), .co(t_3927), .cout(t_3928));
compressor_4_2 u2_1340(.a(s_145_23), .b(s_145_22), .c(s_145_21), .d(s_145_20), .cin(t_3889), .o(t_3929), .co(t_3930), .cout(t_3931));
compressor_4_2 u2_1341(.a(s_145_27), .b(s_145_26), .c(s_145_25), .d(s_145_24), .cin(t_3892), .o(t_3932), .co(t_3933), .cout(t_3934));
compressor_4_2 u2_1342(.a(s_145_31), .b(s_145_30), .c(s_145_29), .d(s_145_28), .cin(t_3895), .o(t_3935), .co(t_3936), .cout(t_3937));
compressor_4_2 u2_1343(.a(s_145_35), .b(s_145_34), .c(s_145_33), .d(s_145_32), .cin(t_3898), .o(t_3938), .co(t_3939), .cout(t_3940));
compressor_4_2 u2_1344(.a(s_145_39), .b(s_145_38), .c(s_145_37), .d(s_145_36), .cin(t_3901), .o(t_3941), .co(t_3942), .cout(t_3943));
compressor_4_2 u2_1345(.a(s_145_43), .b(s_145_42), .c(s_145_41), .d(s_145_40), .cin(t_3904), .o(t_3944), .co(t_3945), .cout(t_3946));
compressor_4_2 u2_1346(.a(s_145_47), .b(s_145_46), .c(s_145_45), .d(s_145_44), .cin(t_3907), .o(t_3947), .co(t_3948), .cout(t_3949));
compressor_4_2 u2_1347(.a(s_145_51), .b(s_145_50), .c(s_145_49), .d(s_145_48), .cin(t_3910), .o(t_3950), .co(t_3951), .cout(t_3952));
compressor_4_2 u2_1348(.a(s_145_55), .b(s_145_54), .c(s_145_53), .d(s_145_52), .cin(t_3913), .o(t_3953), .co(t_3954), .cout(t_3955));
compressor_4_2 u2_1349(.a(s_146_3), .b(s_146_2), .c(s_146_1), .d(s_146_0), .cin(t_3916), .o(t_3956), .co(t_3957), .cout(t_3958));
compressor_4_2 u2_1350(.a(s_146_7), .b(s_146_6), .c(s_146_5), .d(s_146_4), .cin(t_3919), .o(t_3959), .co(t_3960), .cout(t_3961));
compressor_4_2 u2_1351(.a(s_146_11), .b(s_146_10), .c(s_146_9), .d(s_146_8), .cin(t_3922), .o(t_3962), .co(t_3963), .cout(t_3964));
compressor_4_2 u2_1352(.a(s_146_15), .b(s_146_14), .c(s_146_13), .d(s_146_12), .cin(t_3925), .o(t_3965), .co(t_3966), .cout(t_3967));
compressor_4_2 u2_1353(.a(s_146_19), .b(s_146_18), .c(s_146_17), .d(s_146_16), .cin(t_3928), .o(t_3968), .co(t_3969), .cout(t_3970));
compressor_4_2 u2_1354(.a(s_146_23), .b(s_146_22), .c(s_146_21), .d(s_146_20), .cin(t_3931), .o(t_3971), .co(t_3972), .cout(t_3973));
compressor_4_2 u2_1355(.a(s_146_27), .b(s_146_26), .c(s_146_25), .d(s_146_24), .cin(t_3934), .o(t_3974), .co(t_3975), .cout(t_3976));
compressor_4_2 u2_1356(.a(s_146_31), .b(s_146_30), .c(s_146_29), .d(s_146_28), .cin(t_3937), .o(t_3977), .co(t_3978), .cout(t_3979));
compressor_4_2 u2_1357(.a(s_146_35), .b(s_146_34), .c(s_146_33), .d(s_146_32), .cin(t_3940), .o(t_3980), .co(t_3981), .cout(t_3982));
compressor_4_2 u2_1358(.a(s_146_39), .b(s_146_38), .c(s_146_37), .d(s_146_36), .cin(t_3943), .o(t_3983), .co(t_3984), .cout(t_3985));
compressor_4_2 u2_1359(.a(s_146_43), .b(s_146_42), .c(s_146_41), .d(s_146_40), .cin(t_3946), .o(t_3986), .co(t_3987), .cout(t_3988));
compressor_4_2 u2_1360(.a(s_146_47), .b(s_146_46), .c(s_146_45), .d(s_146_44), .cin(t_3949), .o(t_3989), .co(t_3990), .cout(t_3991));
compressor_4_2 u2_1361(.a(s_146_51), .b(s_146_50), .c(s_146_49), .d(s_146_48), .cin(t_3952), .o(t_3992), .co(t_3993), .cout(t_3994));
compressor_4_2 u2_1362(.a(s_146_55), .b(s_146_54), .c(s_146_53), .d(s_146_52), .cin(t_3955), .o(t_3995), .co(t_3996), .cout(t_3997));
compressor_4_2 u2_1363(.a(s_147_3), .b(s_147_2), .c(s_147_1), .d(s_147_0), .cin(t_3958), .o(t_3998), .co(t_3999), .cout(t_4000));
compressor_4_2 u2_1364(.a(s_147_7), .b(s_147_6), .c(s_147_5), .d(s_147_4), .cin(t_3961), .o(t_4001), .co(t_4002), .cout(t_4003));
compressor_4_2 u2_1365(.a(s_147_11), .b(s_147_10), .c(s_147_9), .d(s_147_8), .cin(t_3964), .o(t_4004), .co(t_4005), .cout(t_4006));
compressor_4_2 u2_1366(.a(s_147_15), .b(s_147_14), .c(s_147_13), .d(s_147_12), .cin(t_3967), .o(t_4007), .co(t_4008), .cout(t_4009));
compressor_4_2 u2_1367(.a(s_147_19), .b(s_147_18), .c(s_147_17), .d(s_147_16), .cin(t_3970), .o(t_4010), .co(t_4011), .cout(t_4012));
compressor_4_2 u2_1368(.a(s_147_23), .b(s_147_22), .c(s_147_21), .d(s_147_20), .cin(t_3973), .o(t_4013), .co(t_4014), .cout(t_4015));
compressor_4_2 u2_1369(.a(s_147_27), .b(s_147_26), .c(s_147_25), .d(s_147_24), .cin(t_3976), .o(t_4016), .co(t_4017), .cout(t_4018));
compressor_4_2 u2_1370(.a(s_147_31), .b(s_147_30), .c(s_147_29), .d(s_147_28), .cin(t_3979), .o(t_4019), .co(t_4020), .cout(t_4021));
compressor_4_2 u2_1371(.a(s_147_35), .b(s_147_34), .c(s_147_33), .d(s_147_32), .cin(t_3982), .o(t_4022), .co(t_4023), .cout(t_4024));
compressor_4_2 u2_1372(.a(s_147_39), .b(s_147_38), .c(s_147_37), .d(s_147_36), .cin(t_3985), .o(t_4025), .co(t_4026), .cout(t_4027));
compressor_4_2 u2_1373(.a(s_147_43), .b(s_147_42), .c(s_147_41), .d(s_147_40), .cin(t_3988), .o(t_4028), .co(t_4029), .cout(t_4030));
compressor_4_2 u2_1374(.a(s_147_47), .b(s_147_46), .c(s_147_45), .d(s_147_44), .cin(t_3991), .o(t_4031), .co(t_4032), .cout(t_4033));
compressor_4_2 u2_1375(.a(s_147_51), .b(s_147_50), .c(s_147_49), .d(s_147_48), .cin(t_3994), .o(t_4034), .co(t_4035), .cout(t_4036));
compressor_4_2 u2_1376(.a(s_147_55), .b(s_147_54), .c(s_147_53), .d(s_147_52), .cin(t_3997), .o(t_4037), .co(t_4038), .cout(t_4039));
compressor_4_2 u2_1377(.a(s_148_3), .b(s_148_2), .c(s_148_1), .d(s_148_0), .cin(t_4000), .o(t_4040), .co(t_4041), .cout(t_4042));
compressor_4_2 u2_1378(.a(s_148_7), .b(s_148_6), .c(s_148_5), .d(s_148_4), .cin(t_4003), .o(t_4043), .co(t_4044), .cout(t_4045));
compressor_4_2 u2_1379(.a(s_148_11), .b(s_148_10), .c(s_148_9), .d(s_148_8), .cin(t_4006), .o(t_4046), .co(t_4047), .cout(t_4048));
compressor_4_2 u2_1380(.a(s_148_15), .b(s_148_14), .c(s_148_13), .d(s_148_12), .cin(t_4009), .o(t_4049), .co(t_4050), .cout(t_4051));
compressor_4_2 u2_1381(.a(s_148_19), .b(s_148_18), .c(s_148_17), .d(s_148_16), .cin(t_4012), .o(t_4052), .co(t_4053), .cout(t_4054));
compressor_4_2 u2_1382(.a(s_148_23), .b(s_148_22), .c(s_148_21), .d(s_148_20), .cin(t_4015), .o(t_4055), .co(t_4056), .cout(t_4057));
compressor_4_2 u2_1383(.a(s_148_27), .b(s_148_26), .c(s_148_25), .d(s_148_24), .cin(t_4018), .o(t_4058), .co(t_4059), .cout(t_4060));
compressor_4_2 u2_1384(.a(s_148_31), .b(s_148_30), .c(s_148_29), .d(s_148_28), .cin(t_4021), .o(t_4061), .co(t_4062), .cout(t_4063));
compressor_4_2 u2_1385(.a(s_148_35), .b(s_148_34), .c(s_148_33), .d(s_148_32), .cin(t_4024), .o(t_4064), .co(t_4065), .cout(t_4066));
compressor_4_2 u2_1386(.a(s_148_39), .b(s_148_38), .c(s_148_37), .d(s_148_36), .cin(t_4027), .o(t_4067), .co(t_4068), .cout(t_4069));
compressor_4_2 u2_1387(.a(s_148_43), .b(s_148_42), .c(s_148_41), .d(s_148_40), .cin(t_4030), .o(t_4070), .co(t_4071), .cout(t_4072));
compressor_4_2 u2_1388(.a(s_148_47), .b(s_148_46), .c(s_148_45), .d(s_148_44), .cin(t_4033), .o(t_4073), .co(t_4074), .cout(t_4075));
compressor_4_2 u2_1389(.a(s_148_51), .b(s_148_50), .c(s_148_49), .d(s_148_48), .cin(t_4036), .o(t_4076), .co(t_4077), .cout(t_4078));
compressor_3_2 u1_1390(.a(s_148_53), .b(s_148_52), .cin(t_4039), .o(t_4079), .cout(t_4080));
compressor_4_2 u2_1391(.a(s_149_3), .b(s_149_2), .c(s_149_1), .d(s_149_0), .cin(t_4042), .o(t_4081), .co(t_4082), .cout(t_4083));
compressor_4_2 u2_1392(.a(s_149_7), .b(s_149_6), .c(s_149_5), .d(s_149_4), .cin(t_4045), .o(t_4084), .co(t_4085), .cout(t_4086));
compressor_4_2 u2_1393(.a(s_149_11), .b(s_149_10), .c(s_149_9), .d(s_149_8), .cin(t_4048), .o(t_4087), .co(t_4088), .cout(t_4089));
compressor_4_2 u2_1394(.a(s_149_15), .b(s_149_14), .c(s_149_13), .d(s_149_12), .cin(t_4051), .o(t_4090), .co(t_4091), .cout(t_4092));
compressor_4_2 u2_1395(.a(s_149_19), .b(s_149_18), .c(s_149_17), .d(s_149_16), .cin(t_4054), .o(t_4093), .co(t_4094), .cout(t_4095));
compressor_4_2 u2_1396(.a(s_149_23), .b(s_149_22), .c(s_149_21), .d(s_149_20), .cin(t_4057), .o(t_4096), .co(t_4097), .cout(t_4098));
compressor_4_2 u2_1397(.a(s_149_27), .b(s_149_26), .c(s_149_25), .d(s_149_24), .cin(t_4060), .o(t_4099), .co(t_4100), .cout(t_4101));
compressor_4_2 u2_1398(.a(s_149_31), .b(s_149_30), .c(s_149_29), .d(s_149_28), .cin(t_4063), .o(t_4102), .co(t_4103), .cout(t_4104));
compressor_4_2 u2_1399(.a(s_149_35), .b(s_149_34), .c(s_149_33), .d(s_149_32), .cin(t_4066), .o(t_4105), .co(t_4106), .cout(t_4107));
compressor_4_2 u2_1400(.a(s_149_39), .b(s_149_38), .c(s_149_37), .d(s_149_36), .cin(t_4069), .o(t_4108), .co(t_4109), .cout(t_4110));
compressor_4_2 u2_1401(.a(s_149_43), .b(s_149_42), .c(s_149_41), .d(s_149_40), .cin(t_4072), .o(t_4111), .co(t_4112), .cout(t_4113));
compressor_4_2 u2_1402(.a(s_149_47), .b(s_149_46), .c(s_149_45), .d(s_149_44), .cin(t_4075), .o(t_4114), .co(t_4115), .cout(t_4116));
compressor_4_2 u2_1403(.a(s_149_51), .b(s_149_50), .c(s_149_49), .d(s_149_48), .cin(t_4078), .o(t_4117), .co(t_4118), .cout(t_4119));
compressor_3_2 u1_1404(.a(s_149_54), .b(s_149_53), .cin(s_149_52), .o(t_4120), .cout(t_4121));
compressor_4_2 u2_1405(.a(s_150_3), .b(s_150_2), .c(s_150_1), .d(s_150_0), .cin(t_4083), .o(t_4122), .co(t_4123), .cout(t_4124));
compressor_4_2 u2_1406(.a(s_150_7), .b(s_150_6), .c(s_150_5), .d(s_150_4), .cin(t_4086), .o(t_4125), .co(t_4126), .cout(t_4127));
compressor_4_2 u2_1407(.a(s_150_11), .b(s_150_10), .c(s_150_9), .d(s_150_8), .cin(t_4089), .o(t_4128), .co(t_4129), .cout(t_4130));
compressor_4_2 u2_1408(.a(s_150_15), .b(s_150_14), .c(s_150_13), .d(s_150_12), .cin(t_4092), .o(t_4131), .co(t_4132), .cout(t_4133));
compressor_4_2 u2_1409(.a(s_150_19), .b(s_150_18), .c(s_150_17), .d(s_150_16), .cin(t_4095), .o(t_4134), .co(t_4135), .cout(t_4136));
compressor_4_2 u2_1410(.a(s_150_23), .b(s_150_22), .c(s_150_21), .d(s_150_20), .cin(t_4098), .o(t_4137), .co(t_4138), .cout(t_4139));
compressor_4_2 u2_1411(.a(s_150_27), .b(s_150_26), .c(s_150_25), .d(s_150_24), .cin(t_4101), .o(t_4140), .co(t_4141), .cout(t_4142));
compressor_4_2 u2_1412(.a(s_150_31), .b(s_150_30), .c(s_150_29), .d(s_150_28), .cin(t_4104), .o(t_4143), .co(t_4144), .cout(t_4145));
compressor_4_2 u2_1413(.a(s_150_35), .b(s_150_34), .c(s_150_33), .d(s_150_32), .cin(t_4107), .o(t_4146), .co(t_4147), .cout(t_4148));
compressor_4_2 u2_1414(.a(s_150_39), .b(s_150_38), .c(s_150_37), .d(s_150_36), .cin(t_4110), .o(t_4149), .co(t_4150), .cout(t_4151));
compressor_4_2 u2_1415(.a(s_150_43), .b(s_150_42), .c(s_150_41), .d(s_150_40), .cin(t_4113), .o(t_4152), .co(t_4153), .cout(t_4154));
compressor_4_2 u2_1416(.a(s_150_47), .b(s_150_46), .c(s_150_45), .d(s_150_44), .cin(t_4116), .o(t_4155), .co(t_4156), .cout(t_4157));
compressor_4_2 u2_1417(.a(s_150_51), .b(s_150_50), .c(s_150_49), .d(s_150_48), .cin(t_4119), .o(t_4158), .co(t_4159), .cout(t_4160));
half_adder u0_1418(.a(s_150_53), .b(s_150_52), .o(t_4161), .cout(t_4162));
compressor_4_2 u2_1419(.a(s_151_3), .b(s_151_2), .c(s_151_1), .d(s_151_0), .cin(t_4124), .o(t_4163), .co(t_4164), .cout(t_4165));
compressor_4_2 u2_1420(.a(s_151_7), .b(s_151_6), .c(s_151_5), .d(s_151_4), .cin(t_4127), .o(t_4166), .co(t_4167), .cout(t_4168));
compressor_4_2 u2_1421(.a(s_151_11), .b(s_151_10), .c(s_151_9), .d(s_151_8), .cin(t_4130), .o(t_4169), .co(t_4170), .cout(t_4171));
compressor_4_2 u2_1422(.a(s_151_15), .b(s_151_14), .c(s_151_13), .d(s_151_12), .cin(t_4133), .o(t_4172), .co(t_4173), .cout(t_4174));
compressor_4_2 u2_1423(.a(s_151_19), .b(s_151_18), .c(s_151_17), .d(s_151_16), .cin(t_4136), .o(t_4175), .co(t_4176), .cout(t_4177));
compressor_4_2 u2_1424(.a(s_151_23), .b(s_151_22), .c(s_151_21), .d(s_151_20), .cin(t_4139), .o(t_4178), .co(t_4179), .cout(t_4180));
compressor_4_2 u2_1425(.a(s_151_27), .b(s_151_26), .c(s_151_25), .d(s_151_24), .cin(t_4142), .o(t_4181), .co(t_4182), .cout(t_4183));
compressor_4_2 u2_1426(.a(s_151_31), .b(s_151_30), .c(s_151_29), .d(s_151_28), .cin(t_4145), .o(t_4184), .co(t_4185), .cout(t_4186));
compressor_4_2 u2_1427(.a(s_151_35), .b(s_151_34), .c(s_151_33), .d(s_151_32), .cin(t_4148), .o(t_4187), .co(t_4188), .cout(t_4189));
compressor_4_2 u2_1428(.a(s_151_39), .b(s_151_38), .c(s_151_37), .d(s_151_36), .cin(t_4151), .o(t_4190), .co(t_4191), .cout(t_4192));
compressor_4_2 u2_1429(.a(s_151_43), .b(s_151_42), .c(s_151_41), .d(s_151_40), .cin(t_4154), .o(t_4193), .co(t_4194), .cout(t_4195));
compressor_4_2 u2_1430(.a(s_151_47), .b(s_151_46), .c(s_151_45), .d(s_151_44), .cin(t_4157), .o(t_4196), .co(t_4197), .cout(t_4198));
compressor_4_2 u2_1431(.a(s_151_51), .b(s_151_50), .c(s_151_49), .d(s_151_48), .cin(t_4160), .o(t_4199), .co(t_4200), .cout(t_4201));
half_adder u0_1432(.a(s_151_53), .b(s_151_52), .o(t_4202), .cout(t_4203));
compressor_4_2 u2_1433(.a(s_152_3), .b(s_152_2), .c(s_152_1), .d(s_152_0), .cin(t_4165), .o(t_4204), .co(t_4205), .cout(t_4206));
compressor_4_2 u2_1434(.a(s_152_7), .b(s_152_6), .c(s_152_5), .d(s_152_4), .cin(t_4168), .o(t_4207), .co(t_4208), .cout(t_4209));
compressor_4_2 u2_1435(.a(s_152_11), .b(s_152_10), .c(s_152_9), .d(s_152_8), .cin(t_4171), .o(t_4210), .co(t_4211), .cout(t_4212));
compressor_4_2 u2_1436(.a(s_152_15), .b(s_152_14), .c(s_152_13), .d(s_152_12), .cin(t_4174), .o(t_4213), .co(t_4214), .cout(t_4215));
compressor_4_2 u2_1437(.a(s_152_19), .b(s_152_18), .c(s_152_17), .d(s_152_16), .cin(t_4177), .o(t_4216), .co(t_4217), .cout(t_4218));
compressor_4_2 u2_1438(.a(s_152_23), .b(s_152_22), .c(s_152_21), .d(s_152_20), .cin(t_4180), .o(t_4219), .co(t_4220), .cout(t_4221));
compressor_4_2 u2_1439(.a(s_152_27), .b(s_152_26), .c(s_152_25), .d(s_152_24), .cin(t_4183), .o(t_4222), .co(t_4223), .cout(t_4224));
compressor_4_2 u2_1440(.a(s_152_31), .b(s_152_30), .c(s_152_29), .d(s_152_28), .cin(t_4186), .o(t_4225), .co(t_4226), .cout(t_4227));
compressor_4_2 u2_1441(.a(s_152_35), .b(s_152_34), .c(s_152_33), .d(s_152_32), .cin(t_4189), .o(t_4228), .co(t_4229), .cout(t_4230));
compressor_4_2 u2_1442(.a(s_152_39), .b(s_152_38), .c(s_152_37), .d(s_152_36), .cin(t_4192), .o(t_4231), .co(t_4232), .cout(t_4233));
compressor_4_2 u2_1443(.a(s_152_43), .b(s_152_42), .c(s_152_41), .d(s_152_40), .cin(t_4195), .o(t_4234), .co(t_4235), .cout(t_4236));
compressor_4_2 u2_1444(.a(s_152_47), .b(s_152_46), .c(s_152_45), .d(s_152_44), .cin(t_4198), .o(t_4237), .co(t_4238), .cout(t_4239));
compressor_4_2 u2_1445(.a(s_152_51), .b(s_152_50), .c(s_152_49), .d(s_152_48), .cin(t_4201), .o(t_4240), .co(t_4241), .cout(t_4242));
compressor_4_2 u2_1446(.a(s_153_3), .b(s_153_2), .c(s_153_1), .d(s_153_0), .cin(t_4206), .o(t_4243), .co(t_4244), .cout(t_4245));
compressor_4_2 u2_1447(.a(s_153_7), .b(s_153_6), .c(s_153_5), .d(s_153_4), .cin(t_4209), .o(t_4246), .co(t_4247), .cout(t_4248));
compressor_4_2 u2_1448(.a(s_153_11), .b(s_153_10), .c(s_153_9), .d(s_153_8), .cin(t_4212), .o(t_4249), .co(t_4250), .cout(t_4251));
compressor_4_2 u2_1449(.a(s_153_15), .b(s_153_14), .c(s_153_13), .d(s_153_12), .cin(t_4215), .o(t_4252), .co(t_4253), .cout(t_4254));
compressor_4_2 u2_1450(.a(s_153_19), .b(s_153_18), .c(s_153_17), .d(s_153_16), .cin(t_4218), .o(t_4255), .co(t_4256), .cout(t_4257));
compressor_4_2 u2_1451(.a(s_153_23), .b(s_153_22), .c(s_153_21), .d(s_153_20), .cin(t_4221), .o(t_4258), .co(t_4259), .cout(t_4260));
compressor_4_2 u2_1452(.a(s_153_27), .b(s_153_26), .c(s_153_25), .d(s_153_24), .cin(t_4224), .o(t_4261), .co(t_4262), .cout(t_4263));
compressor_4_2 u2_1453(.a(s_153_31), .b(s_153_30), .c(s_153_29), .d(s_153_28), .cin(t_4227), .o(t_4264), .co(t_4265), .cout(t_4266));
compressor_4_2 u2_1454(.a(s_153_35), .b(s_153_34), .c(s_153_33), .d(s_153_32), .cin(t_4230), .o(t_4267), .co(t_4268), .cout(t_4269));
compressor_4_2 u2_1455(.a(s_153_39), .b(s_153_38), .c(s_153_37), .d(s_153_36), .cin(t_4233), .o(t_4270), .co(t_4271), .cout(t_4272));
compressor_4_2 u2_1456(.a(s_153_43), .b(s_153_42), .c(s_153_41), .d(s_153_40), .cin(t_4236), .o(t_4273), .co(t_4274), .cout(t_4275));
compressor_4_2 u2_1457(.a(s_153_47), .b(s_153_46), .c(s_153_45), .d(s_153_44), .cin(t_4239), .o(t_4276), .co(t_4277), .cout(t_4278));
compressor_4_2 u2_1458(.a(s_153_51), .b(s_153_50), .c(s_153_49), .d(s_153_48), .cin(t_4242), .o(t_4279), .co(t_4280), .cout(t_4281));
compressor_4_2 u2_1459(.a(s_154_3), .b(s_154_2), .c(s_154_1), .d(s_154_0), .cin(t_4245), .o(t_4282), .co(t_4283), .cout(t_4284));
compressor_4_2 u2_1460(.a(s_154_7), .b(s_154_6), .c(s_154_5), .d(s_154_4), .cin(t_4248), .o(t_4285), .co(t_4286), .cout(t_4287));
compressor_4_2 u2_1461(.a(s_154_11), .b(s_154_10), .c(s_154_9), .d(s_154_8), .cin(t_4251), .o(t_4288), .co(t_4289), .cout(t_4290));
compressor_4_2 u2_1462(.a(s_154_15), .b(s_154_14), .c(s_154_13), .d(s_154_12), .cin(t_4254), .o(t_4291), .co(t_4292), .cout(t_4293));
compressor_4_2 u2_1463(.a(s_154_19), .b(s_154_18), .c(s_154_17), .d(s_154_16), .cin(t_4257), .o(t_4294), .co(t_4295), .cout(t_4296));
compressor_4_2 u2_1464(.a(s_154_23), .b(s_154_22), .c(s_154_21), .d(s_154_20), .cin(t_4260), .o(t_4297), .co(t_4298), .cout(t_4299));
compressor_4_2 u2_1465(.a(s_154_27), .b(s_154_26), .c(s_154_25), .d(s_154_24), .cin(t_4263), .o(t_4300), .co(t_4301), .cout(t_4302));
compressor_4_2 u2_1466(.a(s_154_31), .b(s_154_30), .c(s_154_29), .d(s_154_28), .cin(t_4266), .o(t_4303), .co(t_4304), .cout(t_4305));
compressor_4_2 u2_1467(.a(s_154_35), .b(s_154_34), .c(s_154_33), .d(s_154_32), .cin(t_4269), .o(t_4306), .co(t_4307), .cout(t_4308));
compressor_4_2 u2_1468(.a(s_154_39), .b(s_154_38), .c(s_154_37), .d(s_154_36), .cin(t_4272), .o(t_4309), .co(t_4310), .cout(t_4311));
compressor_4_2 u2_1469(.a(s_154_43), .b(s_154_42), .c(s_154_41), .d(s_154_40), .cin(t_4275), .o(t_4312), .co(t_4313), .cout(t_4314));
compressor_4_2 u2_1470(.a(s_154_47), .b(s_154_46), .c(s_154_45), .d(s_154_44), .cin(t_4278), .o(t_4315), .co(t_4316), .cout(t_4317));
compressor_4_2 u2_1471(.a(s_154_51), .b(s_154_50), .c(s_154_49), .d(s_154_48), .cin(t_4281), .o(t_4318), .co(t_4319), .cout(t_4320));
compressor_4_2 u2_1472(.a(s_155_3), .b(s_155_2), .c(s_155_1), .d(s_155_0), .cin(t_4284), .o(t_4321), .co(t_4322), .cout(t_4323));
compressor_4_2 u2_1473(.a(s_155_7), .b(s_155_6), .c(s_155_5), .d(s_155_4), .cin(t_4287), .o(t_4324), .co(t_4325), .cout(t_4326));
compressor_4_2 u2_1474(.a(s_155_11), .b(s_155_10), .c(s_155_9), .d(s_155_8), .cin(t_4290), .o(t_4327), .co(t_4328), .cout(t_4329));
compressor_4_2 u2_1475(.a(s_155_15), .b(s_155_14), .c(s_155_13), .d(s_155_12), .cin(t_4293), .o(t_4330), .co(t_4331), .cout(t_4332));
compressor_4_2 u2_1476(.a(s_155_19), .b(s_155_18), .c(s_155_17), .d(s_155_16), .cin(t_4296), .o(t_4333), .co(t_4334), .cout(t_4335));
compressor_4_2 u2_1477(.a(s_155_23), .b(s_155_22), .c(s_155_21), .d(s_155_20), .cin(t_4299), .o(t_4336), .co(t_4337), .cout(t_4338));
compressor_4_2 u2_1478(.a(s_155_27), .b(s_155_26), .c(s_155_25), .d(s_155_24), .cin(t_4302), .o(t_4339), .co(t_4340), .cout(t_4341));
compressor_4_2 u2_1479(.a(s_155_31), .b(s_155_30), .c(s_155_29), .d(s_155_28), .cin(t_4305), .o(t_4342), .co(t_4343), .cout(t_4344));
compressor_4_2 u2_1480(.a(s_155_35), .b(s_155_34), .c(s_155_33), .d(s_155_32), .cin(t_4308), .o(t_4345), .co(t_4346), .cout(t_4347));
compressor_4_2 u2_1481(.a(s_155_39), .b(s_155_38), .c(s_155_37), .d(s_155_36), .cin(t_4311), .o(t_4348), .co(t_4349), .cout(t_4350));
compressor_4_2 u2_1482(.a(s_155_43), .b(s_155_42), .c(s_155_41), .d(s_155_40), .cin(t_4314), .o(t_4351), .co(t_4352), .cout(t_4353));
compressor_4_2 u2_1483(.a(s_155_47), .b(s_155_46), .c(s_155_45), .d(s_155_44), .cin(t_4317), .o(t_4354), .co(t_4355), .cout(t_4356));
compressor_4_2 u2_1484(.a(s_155_51), .b(s_155_50), .c(s_155_49), .d(s_155_48), .cin(t_4320), .o(t_4357), .co(t_4358), .cout(t_4359));
compressor_4_2 u2_1485(.a(s_156_3), .b(s_156_2), .c(s_156_1), .d(s_156_0), .cin(t_4323), .o(t_4360), .co(t_4361), .cout(t_4362));
compressor_4_2 u2_1486(.a(s_156_7), .b(s_156_6), .c(s_156_5), .d(s_156_4), .cin(t_4326), .o(t_4363), .co(t_4364), .cout(t_4365));
compressor_4_2 u2_1487(.a(s_156_11), .b(s_156_10), .c(s_156_9), .d(s_156_8), .cin(t_4329), .o(t_4366), .co(t_4367), .cout(t_4368));
compressor_4_2 u2_1488(.a(s_156_15), .b(s_156_14), .c(s_156_13), .d(s_156_12), .cin(t_4332), .o(t_4369), .co(t_4370), .cout(t_4371));
compressor_4_2 u2_1489(.a(s_156_19), .b(s_156_18), .c(s_156_17), .d(s_156_16), .cin(t_4335), .o(t_4372), .co(t_4373), .cout(t_4374));
compressor_4_2 u2_1490(.a(s_156_23), .b(s_156_22), .c(s_156_21), .d(s_156_20), .cin(t_4338), .o(t_4375), .co(t_4376), .cout(t_4377));
compressor_4_2 u2_1491(.a(s_156_27), .b(s_156_26), .c(s_156_25), .d(s_156_24), .cin(t_4341), .o(t_4378), .co(t_4379), .cout(t_4380));
compressor_4_2 u2_1492(.a(s_156_31), .b(s_156_30), .c(s_156_29), .d(s_156_28), .cin(t_4344), .o(t_4381), .co(t_4382), .cout(t_4383));
compressor_4_2 u2_1493(.a(s_156_35), .b(s_156_34), .c(s_156_33), .d(s_156_32), .cin(t_4347), .o(t_4384), .co(t_4385), .cout(t_4386));
compressor_4_2 u2_1494(.a(s_156_39), .b(s_156_38), .c(s_156_37), .d(s_156_36), .cin(t_4350), .o(t_4387), .co(t_4388), .cout(t_4389));
compressor_4_2 u2_1495(.a(s_156_43), .b(s_156_42), .c(s_156_41), .d(s_156_40), .cin(t_4353), .o(t_4390), .co(t_4391), .cout(t_4392));
compressor_4_2 u2_1496(.a(s_156_47), .b(s_156_46), .c(s_156_45), .d(s_156_44), .cin(t_4356), .o(t_4393), .co(t_4394), .cout(t_4395));
compressor_3_2 u1_1497(.a(s_156_49), .b(s_156_48), .cin(t_4359), .o(t_4396), .cout(t_4397));
compressor_4_2 u2_1498(.a(s_157_3), .b(s_157_2), .c(s_157_1), .d(s_157_0), .cin(t_4362), .o(t_4398), .co(t_4399), .cout(t_4400));
compressor_4_2 u2_1499(.a(s_157_7), .b(s_157_6), .c(s_157_5), .d(s_157_4), .cin(t_4365), .o(t_4401), .co(t_4402), .cout(t_4403));
compressor_4_2 u2_1500(.a(s_157_11), .b(s_157_10), .c(s_157_9), .d(s_157_8), .cin(t_4368), .o(t_4404), .co(t_4405), .cout(t_4406));
compressor_4_2 u2_1501(.a(s_157_15), .b(s_157_14), .c(s_157_13), .d(s_157_12), .cin(t_4371), .o(t_4407), .co(t_4408), .cout(t_4409));
compressor_4_2 u2_1502(.a(s_157_19), .b(s_157_18), .c(s_157_17), .d(s_157_16), .cin(t_4374), .o(t_4410), .co(t_4411), .cout(t_4412));
compressor_4_2 u2_1503(.a(s_157_23), .b(s_157_22), .c(s_157_21), .d(s_157_20), .cin(t_4377), .o(t_4413), .co(t_4414), .cout(t_4415));
compressor_4_2 u2_1504(.a(s_157_27), .b(s_157_26), .c(s_157_25), .d(s_157_24), .cin(t_4380), .o(t_4416), .co(t_4417), .cout(t_4418));
compressor_4_2 u2_1505(.a(s_157_31), .b(s_157_30), .c(s_157_29), .d(s_157_28), .cin(t_4383), .o(t_4419), .co(t_4420), .cout(t_4421));
compressor_4_2 u2_1506(.a(s_157_35), .b(s_157_34), .c(s_157_33), .d(s_157_32), .cin(t_4386), .o(t_4422), .co(t_4423), .cout(t_4424));
compressor_4_2 u2_1507(.a(s_157_39), .b(s_157_38), .c(s_157_37), .d(s_157_36), .cin(t_4389), .o(t_4425), .co(t_4426), .cout(t_4427));
compressor_4_2 u2_1508(.a(s_157_43), .b(s_157_42), .c(s_157_41), .d(s_157_40), .cin(t_4392), .o(t_4428), .co(t_4429), .cout(t_4430));
compressor_4_2 u2_1509(.a(s_157_47), .b(s_157_46), .c(s_157_45), .d(s_157_44), .cin(t_4395), .o(t_4431), .co(t_4432), .cout(t_4433));
compressor_3_2 u1_1510(.a(s_157_50), .b(s_157_49), .cin(s_157_48), .o(t_4434), .cout(t_4435));
compressor_4_2 u2_1511(.a(s_158_3), .b(s_158_2), .c(s_158_1), .d(s_158_0), .cin(t_4400), .o(t_4436), .co(t_4437), .cout(t_4438));
compressor_4_2 u2_1512(.a(s_158_7), .b(s_158_6), .c(s_158_5), .d(s_158_4), .cin(t_4403), .o(t_4439), .co(t_4440), .cout(t_4441));
compressor_4_2 u2_1513(.a(s_158_11), .b(s_158_10), .c(s_158_9), .d(s_158_8), .cin(t_4406), .o(t_4442), .co(t_4443), .cout(t_4444));
compressor_4_2 u2_1514(.a(s_158_15), .b(s_158_14), .c(s_158_13), .d(s_158_12), .cin(t_4409), .o(t_4445), .co(t_4446), .cout(t_4447));
compressor_4_2 u2_1515(.a(s_158_19), .b(s_158_18), .c(s_158_17), .d(s_158_16), .cin(t_4412), .o(t_4448), .co(t_4449), .cout(t_4450));
compressor_4_2 u2_1516(.a(s_158_23), .b(s_158_22), .c(s_158_21), .d(s_158_20), .cin(t_4415), .o(t_4451), .co(t_4452), .cout(t_4453));
compressor_4_2 u2_1517(.a(s_158_27), .b(s_158_26), .c(s_158_25), .d(s_158_24), .cin(t_4418), .o(t_4454), .co(t_4455), .cout(t_4456));
compressor_4_2 u2_1518(.a(s_158_31), .b(s_158_30), .c(s_158_29), .d(s_158_28), .cin(t_4421), .o(t_4457), .co(t_4458), .cout(t_4459));
compressor_4_2 u2_1519(.a(s_158_35), .b(s_158_34), .c(s_158_33), .d(s_158_32), .cin(t_4424), .o(t_4460), .co(t_4461), .cout(t_4462));
compressor_4_2 u2_1520(.a(s_158_39), .b(s_158_38), .c(s_158_37), .d(s_158_36), .cin(t_4427), .o(t_4463), .co(t_4464), .cout(t_4465));
compressor_4_2 u2_1521(.a(s_158_43), .b(s_158_42), .c(s_158_41), .d(s_158_40), .cin(t_4430), .o(t_4466), .co(t_4467), .cout(t_4468));
compressor_4_2 u2_1522(.a(s_158_47), .b(s_158_46), .c(s_158_45), .d(s_158_44), .cin(t_4433), .o(t_4469), .co(t_4470), .cout(t_4471));
half_adder u0_1523(.a(s_158_49), .b(s_158_48), .o(t_4472), .cout(t_4473));
compressor_4_2 u2_1524(.a(s_159_3), .b(s_159_2), .c(s_159_1), .d(s_159_0), .cin(t_4438), .o(t_4474), .co(t_4475), .cout(t_4476));
compressor_4_2 u2_1525(.a(s_159_7), .b(s_159_6), .c(s_159_5), .d(s_159_4), .cin(t_4441), .o(t_4477), .co(t_4478), .cout(t_4479));
compressor_4_2 u2_1526(.a(s_159_11), .b(s_159_10), .c(s_159_9), .d(s_159_8), .cin(t_4444), .o(t_4480), .co(t_4481), .cout(t_4482));
compressor_4_2 u2_1527(.a(s_159_15), .b(s_159_14), .c(s_159_13), .d(s_159_12), .cin(t_4447), .o(t_4483), .co(t_4484), .cout(t_4485));
compressor_4_2 u2_1528(.a(s_159_19), .b(s_159_18), .c(s_159_17), .d(s_159_16), .cin(t_4450), .o(t_4486), .co(t_4487), .cout(t_4488));
compressor_4_2 u2_1529(.a(s_159_23), .b(s_159_22), .c(s_159_21), .d(s_159_20), .cin(t_4453), .o(t_4489), .co(t_4490), .cout(t_4491));
compressor_4_2 u2_1530(.a(s_159_27), .b(s_159_26), .c(s_159_25), .d(s_159_24), .cin(t_4456), .o(t_4492), .co(t_4493), .cout(t_4494));
compressor_4_2 u2_1531(.a(s_159_31), .b(s_159_30), .c(s_159_29), .d(s_159_28), .cin(t_4459), .o(t_4495), .co(t_4496), .cout(t_4497));
compressor_4_2 u2_1532(.a(s_159_35), .b(s_159_34), .c(s_159_33), .d(s_159_32), .cin(t_4462), .o(t_4498), .co(t_4499), .cout(t_4500));
compressor_4_2 u2_1533(.a(s_159_39), .b(s_159_38), .c(s_159_37), .d(s_159_36), .cin(t_4465), .o(t_4501), .co(t_4502), .cout(t_4503));
compressor_4_2 u2_1534(.a(s_159_43), .b(s_159_42), .c(s_159_41), .d(s_159_40), .cin(t_4468), .o(t_4504), .co(t_4505), .cout(t_4506));
compressor_4_2 u2_1535(.a(s_159_47), .b(s_159_46), .c(s_159_45), .d(s_159_44), .cin(t_4471), .o(t_4507), .co(t_4508), .cout(t_4509));
half_adder u0_1536(.a(s_159_49), .b(s_159_48), .o(t_4510), .cout(t_4511));
compressor_4_2 u2_1537(.a(s_160_3), .b(s_160_2), .c(s_160_1), .d(s_160_0), .cin(t_4476), .o(t_4512), .co(t_4513), .cout(t_4514));
compressor_4_2 u2_1538(.a(s_160_7), .b(s_160_6), .c(s_160_5), .d(s_160_4), .cin(t_4479), .o(t_4515), .co(t_4516), .cout(t_4517));
compressor_4_2 u2_1539(.a(s_160_11), .b(s_160_10), .c(s_160_9), .d(s_160_8), .cin(t_4482), .o(t_4518), .co(t_4519), .cout(t_4520));
compressor_4_2 u2_1540(.a(s_160_15), .b(s_160_14), .c(s_160_13), .d(s_160_12), .cin(t_4485), .o(t_4521), .co(t_4522), .cout(t_4523));
compressor_4_2 u2_1541(.a(s_160_19), .b(s_160_18), .c(s_160_17), .d(s_160_16), .cin(t_4488), .o(t_4524), .co(t_4525), .cout(t_4526));
compressor_4_2 u2_1542(.a(s_160_23), .b(s_160_22), .c(s_160_21), .d(s_160_20), .cin(t_4491), .o(t_4527), .co(t_4528), .cout(t_4529));
compressor_4_2 u2_1543(.a(s_160_27), .b(s_160_26), .c(s_160_25), .d(s_160_24), .cin(t_4494), .o(t_4530), .co(t_4531), .cout(t_4532));
compressor_4_2 u2_1544(.a(s_160_31), .b(s_160_30), .c(s_160_29), .d(s_160_28), .cin(t_4497), .o(t_4533), .co(t_4534), .cout(t_4535));
compressor_4_2 u2_1545(.a(s_160_35), .b(s_160_34), .c(s_160_33), .d(s_160_32), .cin(t_4500), .o(t_4536), .co(t_4537), .cout(t_4538));
compressor_4_2 u2_1546(.a(s_160_39), .b(s_160_38), .c(s_160_37), .d(s_160_36), .cin(t_4503), .o(t_4539), .co(t_4540), .cout(t_4541));
compressor_4_2 u2_1547(.a(s_160_43), .b(s_160_42), .c(s_160_41), .d(s_160_40), .cin(t_4506), .o(t_4542), .co(t_4543), .cout(t_4544));
compressor_4_2 u2_1548(.a(s_160_47), .b(s_160_46), .c(s_160_45), .d(s_160_44), .cin(t_4509), .o(t_4545), .co(t_4546), .cout(t_4547));
compressor_4_2 u2_1549(.a(s_161_3), .b(s_161_2), .c(s_161_1), .d(s_161_0), .cin(t_4514), .o(t_4548), .co(t_4549), .cout(t_4550));
compressor_4_2 u2_1550(.a(s_161_7), .b(s_161_6), .c(s_161_5), .d(s_161_4), .cin(t_4517), .o(t_4551), .co(t_4552), .cout(t_4553));
compressor_4_2 u2_1551(.a(s_161_11), .b(s_161_10), .c(s_161_9), .d(s_161_8), .cin(t_4520), .o(t_4554), .co(t_4555), .cout(t_4556));
compressor_4_2 u2_1552(.a(s_161_15), .b(s_161_14), .c(s_161_13), .d(s_161_12), .cin(t_4523), .o(t_4557), .co(t_4558), .cout(t_4559));
compressor_4_2 u2_1553(.a(s_161_19), .b(s_161_18), .c(s_161_17), .d(s_161_16), .cin(t_4526), .o(t_4560), .co(t_4561), .cout(t_4562));
compressor_4_2 u2_1554(.a(s_161_23), .b(s_161_22), .c(s_161_21), .d(s_161_20), .cin(t_4529), .o(t_4563), .co(t_4564), .cout(t_4565));
compressor_4_2 u2_1555(.a(s_161_27), .b(s_161_26), .c(s_161_25), .d(s_161_24), .cin(t_4532), .o(t_4566), .co(t_4567), .cout(t_4568));
compressor_4_2 u2_1556(.a(s_161_31), .b(s_161_30), .c(s_161_29), .d(s_161_28), .cin(t_4535), .o(t_4569), .co(t_4570), .cout(t_4571));
compressor_4_2 u2_1557(.a(s_161_35), .b(s_161_34), .c(s_161_33), .d(s_161_32), .cin(t_4538), .o(t_4572), .co(t_4573), .cout(t_4574));
compressor_4_2 u2_1558(.a(s_161_39), .b(s_161_38), .c(s_161_37), .d(s_161_36), .cin(t_4541), .o(t_4575), .co(t_4576), .cout(t_4577));
compressor_4_2 u2_1559(.a(s_161_43), .b(s_161_42), .c(s_161_41), .d(s_161_40), .cin(t_4544), .o(t_4578), .co(t_4579), .cout(t_4580));
compressor_4_2 u2_1560(.a(s_161_47), .b(s_161_46), .c(s_161_45), .d(s_161_44), .cin(t_4547), .o(t_4581), .co(t_4582), .cout(t_4583));
compressor_4_2 u2_1561(.a(s_162_3), .b(s_162_2), .c(s_162_1), .d(s_162_0), .cin(t_4550), .o(t_4584), .co(t_4585), .cout(t_4586));
compressor_4_2 u2_1562(.a(s_162_7), .b(s_162_6), .c(s_162_5), .d(s_162_4), .cin(t_4553), .o(t_4587), .co(t_4588), .cout(t_4589));
compressor_4_2 u2_1563(.a(s_162_11), .b(s_162_10), .c(s_162_9), .d(s_162_8), .cin(t_4556), .o(t_4590), .co(t_4591), .cout(t_4592));
compressor_4_2 u2_1564(.a(s_162_15), .b(s_162_14), .c(s_162_13), .d(s_162_12), .cin(t_4559), .o(t_4593), .co(t_4594), .cout(t_4595));
compressor_4_2 u2_1565(.a(s_162_19), .b(s_162_18), .c(s_162_17), .d(s_162_16), .cin(t_4562), .o(t_4596), .co(t_4597), .cout(t_4598));
compressor_4_2 u2_1566(.a(s_162_23), .b(s_162_22), .c(s_162_21), .d(s_162_20), .cin(t_4565), .o(t_4599), .co(t_4600), .cout(t_4601));
compressor_4_2 u2_1567(.a(s_162_27), .b(s_162_26), .c(s_162_25), .d(s_162_24), .cin(t_4568), .o(t_4602), .co(t_4603), .cout(t_4604));
compressor_4_2 u2_1568(.a(s_162_31), .b(s_162_30), .c(s_162_29), .d(s_162_28), .cin(t_4571), .o(t_4605), .co(t_4606), .cout(t_4607));
compressor_4_2 u2_1569(.a(s_162_35), .b(s_162_34), .c(s_162_33), .d(s_162_32), .cin(t_4574), .o(t_4608), .co(t_4609), .cout(t_4610));
compressor_4_2 u2_1570(.a(s_162_39), .b(s_162_38), .c(s_162_37), .d(s_162_36), .cin(t_4577), .o(t_4611), .co(t_4612), .cout(t_4613));
compressor_4_2 u2_1571(.a(s_162_43), .b(s_162_42), .c(s_162_41), .d(s_162_40), .cin(t_4580), .o(t_4614), .co(t_4615), .cout(t_4616));
compressor_4_2 u2_1572(.a(s_162_47), .b(s_162_46), .c(s_162_45), .d(s_162_44), .cin(t_4583), .o(t_4617), .co(t_4618), .cout(t_4619));
compressor_4_2 u2_1573(.a(s_163_3), .b(s_163_2), .c(s_163_1), .d(s_163_0), .cin(t_4586), .o(t_4620), .co(t_4621), .cout(t_4622));
compressor_4_2 u2_1574(.a(s_163_7), .b(s_163_6), .c(s_163_5), .d(s_163_4), .cin(t_4589), .o(t_4623), .co(t_4624), .cout(t_4625));
compressor_4_2 u2_1575(.a(s_163_11), .b(s_163_10), .c(s_163_9), .d(s_163_8), .cin(t_4592), .o(t_4626), .co(t_4627), .cout(t_4628));
compressor_4_2 u2_1576(.a(s_163_15), .b(s_163_14), .c(s_163_13), .d(s_163_12), .cin(t_4595), .o(t_4629), .co(t_4630), .cout(t_4631));
compressor_4_2 u2_1577(.a(s_163_19), .b(s_163_18), .c(s_163_17), .d(s_163_16), .cin(t_4598), .o(t_4632), .co(t_4633), .cout(t_4634));
compressor_4_2 u2_1578(.a(s_163_23), .b(s_163_22), .c(s_163_21), .d(s_163_20), .cin(t_4601), .o(t_4635), .co(t_4636), .cout(t_4637));
compressor_4_2 u2_1579(.a(s_163_27), .b(s_163_26), .c(s_163_25), .d(s_163_24), .cin(t_4604), .o(t_4638), .co(t_4639), .cout(t_4640));
compressor_4_2 u2_1580(.a(s_163_31), .b(s_163_30), .c(s_163_29), .d(s_163_28), .cin(t_4607), .o(t_4641), .co(t_4642), .cout(t_4643));
compressor_4_2 u2_1581(.a(s_163_35), .b(s_163_34), .c(s_163_33), .d(s_163_32), .cin(t_4610), .o(t_4644), .co(t_4645), .cout(t_4646));
compressor_4_2 u2_1582(.a(s_163_39), .b(s_163_38), .c(s_163_37), .d(s_163_36), .cin(t_4613), .o(t_4647), .co(t_4648), .cout(t_4649));
compressor_4_2 u2_1583(.a(s_163_43), .b(s_163_42), .c(s_163_41), .d(s_163_40), .cin(t_4616), .o(t_4650), .co(t_4651), .cout(t_4652));
compressor_4_2 u2_1584(.a(s_163_47), .b(s_163_46), .c(s_163_45), .d(s_163_44), .cin(t_4619), .o(t_4653), .co(t_4654), .cout(t_4655));
compressor_4_2 u2_1585(.a(s_164_3), .b(s_164_2), .c(s_164_1), .d(s_164_0), .cin(t_4622), .o(t_4656), .co(t_4657), .cout(t_4658));
compressor_4_2 u2_1586(.a(s_164_7), .b(s_164_6), .c(s_164_5), .d(s_164_4), .cin(t_4625), .o(t_4659), .co(t_4660), .cout(t_4661));
compressor_4_2 u2_1587(.a(s_164_11), .b(s_164_10), .c(s_164_9), .d(s_164_8), .cin(t_4628), .o(t_4662), .co(t_4663), .cout(t_4664));
compressor_4_2 u2_1588(.a(s_164_15), .b(s_164_14), .c(s_164_13), .d(s_164_12), .cin(t_4631), .o(t_4665), .co(t_4666), .cout(t_4667));
compressor_4_2 u2_1589(.a(s_164_19), .b(s_164_18), .c(s_164_17), .d(s_164_16), .cin(t_4634), .o(t_4668), .co(t_4669), .cout(t_4670));
compressor_4_2 u2_1590(.a(s_164_23), .b(s_164_22), .c(s_164_21), .d(s_164_20), .cin(t_4637), .o(t_4671), .co(t_4672), .cout(t_4673));
compressor_4_2 u2_1591(.a(s_164_27), .b(s_164_26), .c(s_164_25), .d(s_164_24), .cin(t_4640), .o(t_4674), .co(t_4675), .cout(t_4676));
compressor_4_2 u2_1592(.a(s_164_31), .b(s_164_30), .c(s_164_29), .d(s_164_28), .cin(t_4643), .o(t_4677), .co(t_4678), .cout(t_4679));
compressor_4_2 u2_1593(.a(s_164_35), .b(s_164_34), .c(s_164_33), .d(s_164_32), .cin(t_4646), .o(t_4680), .co(t_4681), .cout(t_4682));
compressor_4_2 u2_1594(.a(s_164_39), .b(s_164_38), .c(s_164_37), .d(s_164_36), .cin(t_4649), .o(t_4683), .co(t_4684), .cout(t_4685));
compressor_4_2 u2_1595(.a(s_164_43), .b(s_164_42), .c(s_164_41), .d(s_164_40), .cin(t_4652), .o(t_4686), .co(t_4687), .cout(t_4688));
compressor_3_2 u1_1596(.a(s_164_45), .b(s_164_44), .cin(t_4655), .o(t_4689), .cout(t_4690));
compressor_4_2 u2_1597(.a(s_165_3), .b(s_165_2), .c(s_165_1), .d(s_165_0), .cin(t_4658), .o(t_4691), .co(t_4692), .cout(t_4693));
compressor_4_2 u2_1598(.a(s_165_7), .b(s_165_6), .c(s_165_5), .d(s_165_4), .cin(t_4661), .o(t_4694), .co(t_4695), .cout(t_4696));
compressor_4_2 u2_1599(.a(s_165_11), .b(s_165_10), .c(s_165_9), .d(s_165_8), .cin(t_4664), .o(t_4697), .co(t_4698), .cout(t_4699));
compressor_4_2 u2_1600(.a(s_165_15), .b(s_165_14), .c(s_165_13), .d(s_165_12), .cin(t_4667), .o(t_4700), .co(t_4701), .cout(t_4702));
compressor_4_2 u2_1601(.a(s_165_19), .b(s_165_18), .c(s_165_17), .d(s_165_16), .cin(t_4670), .o(t_4703), .co(t_4704), .cout(t_4705));
compressor_4_2 u2_1602(.a(s_165_23), .b(s_165_22), .c(s_165_21), .d(s_165_20), .cin(t_4673), .o(t_4706), .co(t_4707), .cout(t_4708));
compressor_4_2 u2_1603(.a(s_165_27), .b(s_165_26), .c(s_165_25), .d(s_165_24), .cin(t_4676), .o(t_4709), .co(t_4710), .cout(t_4711));
compressor_4_2 u2_1604(.a(s_165_31), .b(s_165_30), .c(s_165_29), .d(s_165_28), .cin(t_4679), .o(t_4712), .co(t_4713), .cout(t_4714));
compressor_4_2 u2_1605(.a(s_165_35), .b(s_165_34), .c(s_165_33), .d(s_165_32), .cin(t_4682), .o(t_4715), .co(t_4716), .cout(t_4717));
compressor_4_2 u2_1606(.a(s_165_39), .b(s_165_38), .c(s_165_37), .d(s_165_36), .cin(t_4685), .o(t_4718), .co(t_4719), .cout(t_4720));
compressor_4_2 u2_1607(.a(s_165_43), .b(s_165_42), .c(s_165_41), .d(s_165_40), .cin(t_4688), .o(t_4721), .co(t_4722), .cout(t_4723));
compressor_3_2 u1_1608(.a(s_165_46), .b(s_165_45), .cin(s_165_44), .o(t_4724), .cout(t_4725));
compressor_4_2 u2_1609(.a(s_166_3), .b(s_166_2), .c(s_166_1), .d(s_166_0), .cin(t_4693), .o(t_4726), .co(t_4727), .cout(t_4728));
compressor_4_2 u2_1610(.a(s_166_7), .b(s_166_6), .c(s_166_5), .d(s_166_4), .cin(t_4696), .o(t_4729), .co(t_4730), .cout(t_4731));
compressor_4_2 u2_1611(.a(s_166_11), .b(s_166_10), .c(s_166_9), .d(s_166_8), .cin(t_4699), .o(t_4732), .co(t_4733), .cout(t_4734));
compressor_4_2 u2_1612(.a(s_166_15), .b(s_166_14), .c(s_166_13), .d(s_166_12), .cin(t_4702), .o(t_4735), .co(t_4736), .cout(t_4737));
compressor_4_2 u2_1613(.a(s_166_19), .b(s_166_18), .c(s_166_17), .d(s_166_16), .cin(t_4705), .o(t_4738), .co(t_4739), .cout(t_4740));
compressor_4_2 u2_1614(.a(s_166_23), .b(s_166_22), .c(s_166_21), .d(s_166_20), .cin(t_4708), .o(t_4741), .co(t_4742), .cout(t_4743));
compressor_4_2 u2_1615(.a(s_166_27), .b(s_166_26), .c(s_166_25), .d(s_166_24), .cin(t_4711), .o(t_4744), .co(t_4745), .cout(t_4746));
compressor_4_2 u2_1616(.a(s_166_31), .b(s_166_30), .c(s_166_29), .d(s_166_28), .cin(t_4714), .o(t_4747), .co(t_4748), .cout(t_4749));
compressor_4_2 u2_1617(.a(s_166_35), .b(s_166_34), .c(s_166_33), .d(s_166_32), .cin(t_4717), .o(t_4750), .co(t_4751), .cout(t_4752));
compressor_4_2 u2_1618(.a(s_166_39), .b(s_166_38), .c(s_166_37), .d(s_166_36), .cin(t_4720), .o(t_4753), .co(t_4754), .cout(t_4755));
compressor_4_2 u2_1619(.a(s_166_43), .b(s_166_42), .c(s_166_41), .d(s_166_40), .cin(t_4723), .o(t_4756), .co(t_4757), .cout(t_4758));
half_adder u0_1620(.a(s_166_45), .b(s_166_44), .o(t_4759), .cout(t_4760));
compressor_4_2 u2_1621(.a(s_167_3), .b(s_167_2), .c(s_167_1), .d(s_167_0), .cin(t_4728), .o(t_4761), .co(t_4762), .cout(t_4763));
compressor_4_2 u2_1622(.a(s_167_7), .b(s_167_6), .c(s_167_5), .d(s_167_4), .cin(t_4731), .o(t_4764), .co(t_4765), .cout(t_4766));
compressor_4_2 u2_1623(.a(s_167_11), .b(s_167_10), .c(s_167_9), .d(s_167_8), .cin(t_4734), .o(t_4767), .co(t_4768), .cout(t_4769));
compressor_4_2 u2_1624(.a(s_167_15), .b(s_167_14), .c(s_167_13), .d(s_167_12), .cin(t_4737), .o(t_4770), .co(t_4771), .cout(t_4772));
compressor_4_2 u2_1625(.a(s_167_19), .b(s_167_18), .c(s_167_17), .d(s_167_16), .cin(t_4740), .o(t_4773), .co(t_4774), .cout(t_4775));
compressor_4_2 u2_1626(.a(s_167_23), .b(s_167_22), .c(s_167_21), .d(s_167_20), .cin(t_4743), .o(t_4776), .co(t_4777), .cout(t_4778));
compressor_4_2 u2_1627(.a(s_167_27), .b(s_167_26), .c(s_167_25), .d(s_167_24), .cin(t_4746), .o(t_4779), .co(t_4780), .cout(t_4781));
compressor_4_2 u2_1628(.a(s_167_31), .b(s_167_30), .c(s_167_29), .d(s_167_28), .cin(t_4749), .o(t_4782), .co(t_4783), .cout(t_4784));
compressor_4_2 u2_1629(.a(s_167_35), .b(s_167_34), .c(s_167_33), .d(s_167_32), .cin(t_4752), .o(t_4785), .co(t_4786), .cout(t_4787));
compressor_4_2 u2_1630(.a(s_167_39), .b(s_167_38), .c(s_167_37), .d(s_167_36), .cin(t_4755), .o(t_4788), .co(t_4789), .cout(t_4790));
compressor_4_2 u2_1631(.a(s_167_43), .b(s_167_42), .c(s_167_41), .d(s_167_40), .cin(t_4758), .o(t_4791), .co(t_4792), .cout(t_4793));
half_adder u0_1632(.a(s_167_45), .b(s_167_44), .o(t_4794), .cout(t_4795));
compressor_4_2 u2_1633(.a(s_168_3), .b(s_168_2), .c(s_168_1), .d(s_168_0), .cin(t_4763), .o(t_4796), .co(t_4797), .cout(t_4798));
compressor_4_2 u2_1634(.a(s_168_7), .b(s_168_6), .c(s_168_5), .d(s_168_4), .cin(t_4766), .o(t_4799), .co(t_4800), .cout(t_4801));
compressor_4_2 u2_1635(.a(s_168_11), .b(s_168_10), .c(s_168_9), .d(s_168_8), .cin(t_4769), .o(t_4802), .co(t_4803), .cout(t_4804));
compressor_4_2 u2_1636(.a(s_168_15), .b(s_168_14), .c(s_168_13), .d(s_168_12), .cin(t_4772), .o(t_4805), .co(t_4806), .cout(t_4807));
compressor_4_2 u2_1637(.a(s_168_19), .b(s_168_18), .c(s_168_17), .d(s_168_16), .cin(t_4775), .o(t_4808), .co(t_4809), .cout(t_4810));
compressor_4_2 u2_1638(.a(s_168_23), .b(s_168_22), .c(s_168_21), .d(s_168_20), .cin(t_4778), .o(t_4811), .co(t_4812), .cout(t_4813));
compressor_4_2 u2_1639(.a(s_168_27), .b(s_168_26), .c(s_168_25), .d(s_168_24), .cin(t_4781), .o(t_4814), .co(t_4815), .cout(t_4816));
compressor_4_2 u2_1640(.a(s_168_31), .b(s_168_30), .c(s_168_29), .d(s_168_28), .cin(t_4784), .o(t_4817), .co(t_4818), .cout(t_4819));
compressor_4_2 u2_1641(.a(s_168_35), .b(s_168_34), .c(s_168_33), .d(s_168_32), .cin(t_4787), .o(t_4820), .co(t_4821), .cout(t_4822));
compressor_4_2 u2_1642(.a(s_168_39), .b(s_168_38), .c(s_168_37), .d(s_168_36), .cin(t_4790), .o(t_4823), .co(t_4824), .cout(t_4825));
compressor_4_2 u2_1643(.a(s_168_43), .b(s_168_42), .c(s_168_41), .d(s_168_40), .cin(t_4793), .o(t_4826), .co(t_4827), .cout(t_4828));
compressor_4_2 u2_1644(.a(s_169_3), .b(s_169_2), .c(s_169_1), .d(s_169_0), .cin(t_4798), .o(t_4829), .co(t_4830), .cout(t_4831));
compressor_4_2 u2_1645(.a(s_169_7), .b(s_169_6), .c(s_169_5), .d(s_169_4), .cin(t_4801), .o(t_4832), .co(t_4833), .cout(t_4834));
compressor_4_2 u2_1646(.a(s_169_11), .b(s_169_10), .c(s_169_9), .d(s_169_8), .cin(t_4804), .o(t_4835), .co(t_4836), .cout(t_4837));
compressor_4_2 u2_1647(.a(s_169_15), .b(s_169_14), .c(s_169_13), .d(s_169_12), .cin(t_4807), .o(t_4838), .co(t_4839), .cout(t_4840));
compressor_4_2 u2_1648(.a(s_169_19), .b(s_169_18), .c(s_169_17), .d(s_169_16), .cin(t_4810), .o(t_4841), .co(t_4842), .cout(t_4843));
compressor_4_2 u2_1649(.a(s_169_23), .b(s_169_22), .c(s_169_21), .d(s_169_20), .cin(t_4813), .o(t_4844), .co(t_4845), .cout(t_4846));
compressor_4_2 u2_1650(.a(s_169_27), .b(s_169_26), .c(s_169_25), .d(s_169_24), .cin(t_4816), .o(t_4847), .co(t_4848), .cout(t_4849));
compressor_4_2 u2_1651(.a(s_169_31), .b(s_169_30), .c(s_169_29), .d(s_169_28), .cin(t_4819), .o(t_4850), .co(t_4851), .cout(t_4852));
compressor_4_2 u2_1652(.a(s_169_35), .b(s_169_34), .c(s_169_33), .d(s_169_32), .cin(t_4822), .o(t_4853), .co(t_4854), .cout(t_4855));
compressor_4_2 u2_1653(.a(s_169_39), .b(s_169_38), .c(s_169_37), .d(s_169_36), .cin(t_4825), .o(t_4856), .co(t_4857), .cout(t_4858));
compressor_4_2 u2_1654(.a(s_169_43), .b(s_169_42), .c(s_169_41), .d(s_169_40), .cin(t_4828), .o(t_4859), .co(t_4860), .cout(t_4861));
compressor_4_2 u2_1655(.a(s_170_3), .b(s_170_2), .c(s_170_1), .d(s_170_0), .cin(t_4831), .o(t_4862), .co(t_4863), .cout(t_4864));
compressor_4_2 u2_1656(.a(s_170_7), .b(s_170_6), .c(s_170_5), .d(s_170_4), .cin(t_4834), .o(t_4865), .co(t_4866), .cout(t_4867));
compressor_4_2 u2_1657(.a(s_170_11), .b(s_170_10), .c(s_170_9), .d(s_170_8), .cin(t_4837), .o(t_4868), .co(t_4869), .cout(t_4870));
compressor_4_2 u2_1658(.a(s_170_15), .b(s_170_14), .c(s_170_13), .d(s_170_12), .cin(t_4840), .o(t_4871), .co(t_4872), .cout(t_4873));
compressor_4_2 u2_1659(.a(s_170_19), .b(s_170_18), .c(s_170_17), .d(s_170_16), .cin(t_4843), .o(t_4874), .co(t_4875), .cout(t_4876));
compressor_4_2 u2_1660(.a(s_170_23), .b(s_170_22), .c(s_170_21), .d(s_170_20), .cin(t_4846), .o(t_4877), .co(t_4878), .cout(t_4879));
compressor_4_2 u2_1661(.a(s_170_27), .b(s_170_26), .c(s_170_25), .d(s_170_24), .cin(t_4849), .o(t_4880), .co(t_4881), .cout(t_4882));
compressor_4_2 u2_1662(.a(s_170_31), .b(s_170_30), .c(s_170_29), .d(s_170_28), .cin(t_4852), .o(t_4883), .co(t_4884), .cout(t_4885));
compressor_4_2 u2_1663(.a(s_170_35), .b(s_170_34), .c(s_170_33), .d(s_170_32), .cin(t_4855), .o(t_4886), .co(t_4887), .cout(t_4888));
compressor_4_2 u2_1664(.a(s_170_39), .b(s_170_38), .c(s_170_37), .d(s_170_36), .cin(t_4858), .o(t_4889), .co(t_4890), .cout(t_4891));
compressor_4_2 u2_1665(.a(s_170_43), .b(s_170_42), .c(s_170_41), .d(s_170_40), .cin(t_4861), .o(t_4892), .co(t_4893), .cout(t_4894));
compressor_4_2 u2_1666(.a(s_171_3), .b(s_171_2), .c(s_171_1), .d(s_171_0), .cin(t_4864), .o(t_4895), .co(t_4896), .cout(t_4897));
compressor_4_2 u2_1667(.a(s_171_7), .b(s_171_6), .c(s_171_5), .d(s_171_4), .cin(t_4867), .o(t_4898), .co(t_4899), .cout(t_4900));
compressor_4_2 u2_1668(.a(s_171_11), .b(s_171_10), .c(s_171_9), .d(s_171_8), .cin(t_4870), .o(t_4901), .co(t_4902), .cout(t_4903));
compressor_4_2 u2_1669(.a(s_171_15), .b(s_171_14), .c(s_171_13), .d(s_171_12), .cin(t_4873), .o(t_4904), .co(t_4905), .cout(t_4906));
compressor_4_2 u2_1670(.a(s_171_19), .b(s_171_18), .c(s_171_17), .d(s_171_16), .cin(t_4876), .o(t_4907), .co(t_4908), .cout(t_4909));
compressor_4_2 u2_1671(.a(s_171_23), .b(s_171_22), .c(s_171_21), .d(s_171_20), .cin(t_4879), .o(t_4910), .co(t_4911), .cout(t_4912));
compressor_4_2 u2_1672(.a(s_171_27), .b(s_171_26), .c(s_171_25), .d(s_171_24), .cin(t_4882), .o(t_4913), .co(t_4914), .cout(t_4915));
compressor_4_2 u2_1673(.a(s_171_31), .b(s_171_30), .c(s_171_29), .d(s_171_28), .cin(t_4885), .o(t_4916), .co(t_4917), .cout(t_4918));
compressor_4_2 u2_1674(.a(s_171_35), .b(s_171_34), .c(s_171_33), .d(s_171_32), .cin(t_4888), .o(t_4919), .co(t_4920), .cout(t_4921));
compressor_4_2 u2_1675(.a(s_171_39), .b(s_171_38), .c(s_171_37), .d(s_171_36), .cin(t_4891), .o(t_4922), .co(t_4923), .cout(t_4924));
compressor_4_2 u2_1676(.a(s_171_43), .b(s_171_42), .c(s_171_41), .d(s_171_40), .cin(t_4894), .o(t_4925), .co(t_4926), .cout(t_4927));
compressor_4_2 u2_1677(.a(s_172_3), .b(s_172_2), .c(s_172_1), .d(s_172_0), .cin(t_4897), .o(t_4928), .co(t_4929), .cout(t_4930));
compressor_4_2 u2_1678(.a(s_172_7), .b(s_172_6), .c(s_172_5), .d(s_172_4), .cin(t_4900), .o(t_4931), .co(t_4932), .cout(t_4933));
compressor_4_2 u2_1679(.a(s_172_11), .b(s_172_10), .c(s_172_9), .d(s_172_8), .cin(t_4903), .o(t_4934), .co(t_4935), .cout(t_4936));
compressor_4_2 u2_1680(.a(s_172_15), .b(s_172_14), .c(s_172_13), .d(s_172_12), .cin(t_4906), .o(t_4937), .co(t_4938), .cout(t_4939));
compressor_4_2 u2_1681(.a(s_172_19), .b(s_172_18), .c(s_172_17), .d(s_172_16), .cin(t_4909), .o(t_4940), .co(t_4941), .cout(t_4942));
compressor_4_2 u2_1682(.a(s_172_23), .b(s_172_22), .c(s_172_21), .d(s_172_20), .cin(t_4912), .o(t_4943), .co(t_4944), .cout(t_4945));
compressor_4_2 u2_1683(.a(s_172_27), .b(s_172_26), .c(s_172_25), .d(s_172_24), .cin(t_4915), .o(t_4946), .co(t_4947), .cout(t_4948));
compressor_4_2 u2_1684(.a(s_172_31), .b(s_172_30), .c(s_172_29), .d(s_172_28), .cin(t_4918), .o(t_4949), .co(t_4950), .cout(t_4951));
compressor_4_2 u2_1685(.a(s_172_35), .b(s_172_34), .c(s_172_33), .d(s_172_32), .cin(t_4921), .o(t_4952), .co(t_4953), .cout(t_4954));
compressor_4_2 u2_1686(.a(s_172_39), .b(s_172_38), .c(s_172_37), .d(s_172_36), .cin(t_4924), .o(t_4955), .co(t_4956), .cout(t_4957));
compressor_3_2 u1_1687(.a(s_172_41), .b(s_172_40), .cin(t_4927), .o(t_4958), .cout(t_4959));
compressor_4_2 u2_1688(.a(s_173_3), .b(s_173_2), .c(s_173_1), .d(s_173_0), .cin(t_4930), .o(t_4960), .co(t_4961), .cout(t_4962));
compressor_4_2 u2_1689(.a(s_173_7), .b(s_173_6), .c(s_173_5), .d(s_173_4), .cin(t_4933), .o(t_4963), .co(t_4964), .cout(t_4965));
compressor_4_2 u2_1690(.a(s_173_11), .b(s_173_10), .c(s_173_9), .d(s_173_8), .cin(t_4936), .o(t_4966), .co(t_4967), .cout(t_4968));
compressor_4_2 u2_1691(.a(s_173_15), .b(s_173_14), .c(s_173_13), .d(s_173_12), .cin(t_4939), .o(t_4969), .co(t_4970), .cout(t_4971));
compressor_4_2 u2_1692(.a(s_173_19), .b(s_173_18), .c(s_173_17), .d(s_173_16), .cin(t_4942), .o(t_4972), .co(t_4973), .cout(t_4974));
compressor_4_2 u2_1693(.a(s_173_23), .b(s_173_22), .c(s_173_21), .d(s_173_20), .cin(t_4945), .o(t_4975), .co(t_4976), .cout(t_4977));
compressor_4_2 u2_1694(.a(s_173_27), .b(s_173_26), .c(s_173_25), .d(s_173_24), .cin(t_4948), .o(t_4978), .co(t_4979), .cout(t_4980));
compressor_4_2 u2_1695(.a(s_173_31), .b(s_173_30), .c(s_173_29), .d(s_173_28), .cin(t_4951), .o(t_4981), .co(t_4982), .cout(t_4983));
compressor_4_2 u2_1696(.a(s_173_35), .b(s_173_34), .c(s_173_33), .d(s_173_32), .cin(t_4954), .o(t_4984), .co(t_4985), .cout(t_4986));
compressor_4_2 u2_1697(.a(s_173_39), .b(s_173_38), .c(s_173_37), .d(s_173_36), .cin(t_4957), .o(t_4987), .co(t_4988), .cout(t_4989));
compressor_3_2 u1_1698(.a(s_173_42), .b(s_173_41), .cin(s_173_40), .o(t_4990), .cout(t_4991));
compressor_4_2 u2_1699(.a(s_174_3), .b(s_174_2), .c(s_174_1), .d(s_174_0), .cin(t_4962), .o(t_4992), .co(t_4993), .cout(t_4994));
compressor_4_2 u2_1700(.a(s_174_7), .b(s_174_6), .c(s_174_5), .d(s_174_4), .cin(t_4965), .o(t_4995), .co(t_4996), .cout(t_4997));
compressor_4_2 u2_1701(.a(s_174_11), .b(s_174_10), .c(s_174_9), .d(s_174_8), .cin(t_4968), .o(t_4998), .co(t_4999), .cout(t_5000));
compressor_4_2 u2_1702(.a(s_174_15), .b(s_174_14), .c(s_174_13), .d(s_174_12), .cin(t_4971), .o(t_5001), .co(t_5002), .cout(t_5003));
compressor_4_2 u2_1703(.a(s_174_19), .b(s_174_18), .c(s_174_17), .d(s_174_16), .cin(t_4974), .o(t_5004), .co(t_5005), .cout(t_5006));
compressor_4_2 u2_1704(.a(s_174_23), .b(s_174_22), .c(s_174_21), .d(s_174_20), .cin(t_4977), .o(t_5007), .co(t_5008), .cout(t_5009));
compressor_4_2 u2_1705(.a(s_174_27), .b(s_174_26), .c(s_174_25), .d(s_174_24), .cin(t_4980), .o(t_5010), .co(t_5011), .cout(t_5012));
compressor_4_2 u2_1706(.a(s_174_31), .b(s_174_30), .c(s_174_29), .d(s_174_28), .cin(t_4983), .o(t_5013), .co(t_5014), .cout(t_5015));
compressor_4_2 u2_1707(.a(s_174_35), .b(s_174_34), .c(s_174_33), .d(s_174_32), .cin(t_4986), .o(t_5016), .co(t_5017), .cout(t_5018));
compressor_4_2 u2_1708(.a(s_174_39), .b(s_174_38), .c(s_174_37), .d(s_174_36), .cin(t_4989), .o(t_5019), .co(t_5020), .cout(t_5021));
half_adder u0_1709(.a(s_174_41), .b(s_174_40), .o(t_5022), .cout(t_5023));
compressor_4_2 u2_1710(.a(s_175_3), .b(s_175_2), .c(s_175_1), .d(s_175_0), .cin(t_4994), .o(t_5024), .co(t_5025), .cout(t_5026));
compressor_4_2 u2_1711(.a(s_175_7), .b(s_175_6), .c(s_175_5), .d(s_175_4), .cin(t_4997), .o(t_5027), .co(t_5028), .cout(t_5029));
compressor_4_2 u2_1712(.a(s_175_11), .b(s_175_10), .c(s_175_9), .d(s_175_8), .cin(t_5000), .o(t_5030), .co(t_5031), .cout(t_5032));
compressor_4_2 u2_1713(.a(s_175_15), .b(s_175_14), .c(s_175_13), .d(s_175_12), .cin(t_5003), .o(t_5033), .co(t_5034), .cout(t_5035));
compressor_4_2 u2_1714(.a(s_175_19), .b(s_175_18), .c(s_175_17), .d(s_175_16), .cin(t_5006), .o(t_5036), .co(t_5037), .cout(t_5038));
compressor_4_2 u2_1715(.a(s_175_23), .b(s_175_22), .c(s_175_21), .d(s_175_20), .cin(t_5009), .o(t_5039), .co(t_5040), .cout(t_5041));
compressor_4_2 u2_1716(.a(s_175_27), .b(s_175_26), .c(s_175_25), .d(s_175_24), .cin(t_5012), .o(t_5042), .co(t_5043), .cout(t_5044));
compressor_4_2 u2_1717(.a(s_175_31), .b(s_175_30), .c(s_175_29), .d(s_175_28), .cin(t_5015), .o(t_5045), .co(t_5046), .cout(t_5047));
compressor_4_2 u2_1718(.a(s_175_35), .b(s_175_34), .c(s_175_33), .d(s_175_32), .cin(t_5018), .o(t_5048), .co(t_5049), .cout(t_5050));
compressor_4_2 u2_1719(.a(s_175_39), .b(s_175_38), .c(s_175_37), .d(s_175_36), .cin(t_5021), .o(t_5051), .co(t_5052), .cout(t_5053));
half_adder u0_1720(.a(s_175_41), .b(s_175_40), .o(t_5054), .cout(t_5055));
compressor_4_2 u2_1721(.a(s_176_3), .b(s_176_2), .c(s_176_1), .d(s_176_0), .cin(t_5026), .o(t_5056), .co(t_5057), .cout(t_5058));
compressor_4_2 u2_1722(.a(s_176_7), .b(s_176_6), .c(s_176_5), .d(s_176_4), .cin(t_5029), .o(t_5059), .co(t_5060), .cout(t_5061));
compressor_4_2 u2_1723(.a(s_176_11), .b(s_176_10), .c(s_176_9), .d(s_176_8), .cin(t_5032), .o(t_5062), .co(t_5063), .cout(t_5064));
compressor_4_2 u2_1724(.a(s_176_15), .b(s_176_14), .c(s_176_13), .d(s_176_12), .cin(t_5035), .o(t_5065), .co(t_5066), .cout(t_5067));
compressor_4_2 u2_1725(.a(s_176_19), .b(s_176_18), .c(s_176_17), .d(s_176_16), .cin(t_5038), .o(t_5068), .co(t_5069), .cout(t_5070));
compressor_4_2 u2_1726(.a(s_176_23), .b(s_176_22), .c(s_176_21), .d(s_176_20), .cin(t_5041), .o(t_5071), .co(t_5072), .cout(t_5073));
compressor_4_2 u2_1727(.a(s_176_27), .b(s_176_26), .c(s_176_25), .d(s_176_24), .cin(t_5044), .o(t_5074), .co(t_5075), .cout(t_5076));
compressor_4_2 u2_1728(.a(s_176_31), .b(s_176_30), .c(s_176_29), .d(s_176_28), .cin(t_5047), .o(t_5077), .co(t_5078), .cout(t_5079));
compressor_4_2 u2_1729(.a(s_176_35), .b(s_176_34), .c(s_176_33), .d(s_176_32), .cin(t_5050), .o(t_5080), .co(t_5081), .cout(t_5082));
compressor_4_2 u2_1730(.a(s_176_39), .b(s_176_38), .c(s_176_37), .d(s_176_36), .cin(t_5053), .o(t_5083), .co(t_5084), .cout(t_5085));
compressor_4_2 u2_1731(.a(s_177_3), .b(s_177_2), .c(s_177_1), .d(s_177_0), .cin(t_5058), .o(t_5086), .co(t_5087), .cout(t_5088));
compressor_4_2 u2_1732(.a(s_177_7), .b(s_177_6), .c(s_177_5), .d(s_177_4), .cin(t_5061), .o(t_5089), .co(t_5090), .cout(t_5091));
compressor_4_2 u2_1733(.a(s_177_11), .b(s_177_10), .c(s_177_9), .d(s_177_8), .cin(t_5064), .o(t_5092), .co(t_5093), .cout(t_5094));
compressor_4_2 u2_1734(.a(s_177_15), .b(s_177_14), .c(s_177_13), .d(s_177_12), .cin(t_5067), .o(t_5095), .co(t_5096), .cout(t_5097));
compressor_4_2 u2_1735(.a(s_177_19), .b(s_177_18), .c(s_177_17), .d(s_177_16), .cin(t_5070), .o(t_5098), .co(t_5099), .cout(t_5100));
compressor_4_2 u2_1736(.a(s_177_23), .b(s_177_22), .c(s_177_21), .d(s_177_20), .cin(t_5073), .o(t_5101), .co(t_5102), .cout(t_5103));
compressor_4_2 u2_1737(.a(s_177_27), .b(s_177_26), .c(s_177_25), .d(s_177_24), .cin(t_5076), .o(t_5104), .co(t_5105), .cout(t_5106));
compressor_4_2 u2_1738(.a(s_177_31), .b(s_177_30), .c(s_177_29), .d(s_177_28), .cin(t_5079), .o(t_5107), .co(t_5108), .cout(t_5109));
compressor_4_2 u2_1739(.a(s_177_35), .b(s_177_34), .c(s_177_33), .d(s_177_32), .cin(t_5082), .o(t_5110), .co(t_5111), .cout(t_5112));
compressor_4_2 u2_1740(.a(s_177_39), .b(s_177_38), .c(s_177_37), .d(s_177_36), .cin(t_5085), .o(t_5113), .co(t_5114), .cout(t_5115));
compressor_4_2 u2_1741(.a(s_178_3), .b(s_178_2), .c(s_178_1), .d(s_178_0), .cin(t_5088), .o(t_5116), .co(t_5117), .cout(t_5118));
compressor_4_2 u2_1742(.a(s_178_7), .b(s_178_6), .c(s_178_5), .d(s_178_4), .cin(t_5091), .o(t_5119), .co(t_5120), .cout(t_5121));
compressor_4_2 u2_1743(.a(s_178_11), .b(s_178_10), .c(s_178_9), .d(s_178_8), .cin(t_5094), .o(t_5122), .co(t_5123), .cout(t_5124));
compressor_4_2 u2_1744(.a(s_178_15), .b(s_178_14), .c(s_178_13), .d(s_178_12), .cin(t_5097), .o(t_5125), .co(t_5126), .cout(t_5127));
compressor_4_2 u2_1745(.a(s_178_19), .b(s_178_18), .c(s_178_17), .d(s_178_16), .cin(t_5100), .o(t_5128), .co(t_5129), .cout(t_5130));
compressor_4_2 u2_1746(.a(s_178_23), .b(s_178_22), .c(s_178_21), .d(s_178_20), .cin(t_5103), .o(t_5131), .co(t_5132), .cout(t_5133));
compressor_4_2 u2_1747(.a(s_178_27), .b(s_178_26), .c(s_178_25), .d(s_178_24), .cin(t_5106), .o(t_5134), .co(t_5135), .cout(t_5136));
compressor_4_2 u2_1748(.a(s_178_31), .b(s_178_30), .c(s_178_29), .d(s_178_28), .cin(t_5109), .o(t_5137), .co(t_5138), .cout(t_5139));
compressor_4_2 u2_1749(.a(s_178_35), .b(s_178_34), .c(s_178_33), .d(s_178_32), .cin(t_5112), .o(t_5140), .co(t_5141), .cout(t_5142));
compressor_4_2 u2_1750(.a(s_178_39), .b(s_178_38), .c(s_178_37), .d(s_178_36), .cin(t_5115), .o(t_5143), .co(t_5144), .cout(t_5145));
compressor_4_2 u2_1751(.a(s_179_3), .b(s_179_2), .c(s_179_1), .d(s_179_0), .cin(t_5118), .o(t_5146), .co(t_5147), .cout(t_5148));
compressor_4_2 u2_1752(.a(s_179_7), .b(s_179_6), .c(s_179_5), .d(s_179_4), .cin(t_5121), .o(t_5149), .co(t_5150), .cout(t_5151));
compressor_4_2 u2_1753(.a(s_179_11), .b(s_179_10), .c(s_179_9), .d(s_179_8), .cin(t_5124), .o(t_5152), .co(t_5153), .cout(t_5154));
compressor_4_2 u2_1754(.a(s_179_15), .b(s_179_14), .c(s_179_13), .d(s_179_12), .cin(t_5127), .o(t_5155), .co(t_5156), .cout(t_5157));
compressor_4_2 u2_1755(.a(s_179_19), .b(s_179_18), .c(s_179_17), .d(s_179_16), .cin(t_5130), .o(t_5158), .co(t_5159), .cout(t_5160));
compressor_4_2 u2_1756(.a(s_179_23), .b(s_179_22), .c(s_179_21), .d(s_179_20), .cin(t_5133), .o(t_5161), .co(t_5162), .cout(t_5163));
compressor_4_2 u2_1757(.a(s_179_27), .b(s_179_26), .c(s_179_25), .d(s_179_24), .cin(t_5136), .o(t_5164), .co(t_5165), .cout(t_5166));
compressor_4_2 u2_1758(.a(s_179_31), .b(s_179_30), .c(s_179_29), .d(s_179_28), .cin(t_5139), .o(t_5167), .co(t_5168), .cout(t_5169));
compressor_4_2 u2_1759(.a(s_179_35), .b(s_179_34), .c(s_179_33), .d(s_179_32), .cin(t_5142), .o(t_5170), .co(t_5171), .cout(t_5172));
compressor_4_2 u2_1760(.a(s_179_39), .b(s_179_38), .c(s_179_37), .d(s_179_36), .cin(t_5145), .o(t_5173), .co(t_5174), .cout(t_5175));
compressor_4_2 u2_1761(.a(s_180_3), .b(s_180_2), .c(s_180_1), .d(s_180_0), .cin(t_5148), .o(t_5176), .co(t_5177), .cout(t_5178));
compressor_4_2 u2_1762(.a(s_180_7), .b(s_180_6), .c(s_180_5), .d(s_180_4), .cin(t_5151), .o(t_5179), .co(t_5180), .cout(t_5181));
compressor_4_2 u2_1763(.a(s_180_11), .b(s_180_10), .c(s_180_9), .d(s_180_8), .cin(t_5154), .o(t_5182), .co(t_5183), .cout(t_5184));
compressor_4_2 u2_1764(.a(s_180_15), .b(s_180_14), .c(s_180_13), .d(s_180_12), .cin(t_5157), .o(t_5185), .co(t_5186), .cout(t_5187));
compressor_4_2 u2_1765(.a(s_180_19), .b(s_180_18), .c(s_180_17), .d(s_180_16), .cin(t_5160), .o(t_5188), .co(t_5189), .cout(t_5190));
compressor_4_2 u2_1766(.a(s_180_23), .b(s_180_22), .c(s_180_21), .d(s_180_20), .cin(t_5163), .o(t_5191), .co(t_5192), .cout(t_5193));
compressor_4_2 u2_1767(.a(s_180_27), .b(s_180_26), .c(s_180_25), .d(s_180_24), .cin(t_5166), .o(t_5194), .co(t_5195), .cout(t_5196));
compressor_4_2 u2_1768(.a(s_180_31), .b(s_180_30), .c(s_180_29), .d(s_180_28), .cin(t_5169), .o(t_5197), .co(t_5198), .cout(t_5199));
compressor_4_2 u2_1769(.a(s_180_35), .b(s_180_34), .c(s_180_33), .d(s_180_32), .cin(t_5172), .o(t_5200), .co(t_5201), .cout(t_5202));
compressor_3_2 u1_1770(.a(s_180_37), .b(s_180_36), .cin(t_5175), .o(t_5203), .cout(t_5204));
compressor_4_2 u2_1771(.a(s_181_3), .b(s_181_2), .c(s_181_1), .d(s_181_0), .cin(t_5178), .o(t_5205), .co(t_5206), .cout(t_5207));
compressor_4_2 u2_1772(.a(s_181_7), .b(s_181_6), .c(s_181_5), .d(s_181_4), .cin(t_5181), .o(t_5208), .co(t_5209), .cout(t_5210));
compressor_4_2 u2_1773(.a(s_181_11), .b(s_181_10), .c(s_181_9), .d(s_181_8), .cin(t_5184), .o(t_5211), .co(t_5212), .cout(t_5213));
compressor_4_2 u2_1774(.a(s_181_15), .b(s_181_14), .c(s_181_13), .d(s_181_12), .cin(t_5187), .o(t_5214), .co(t_5215), .cout(t_5216));
compressor_4_2 u2_1775(.a(s_181_19), .b(s_181_18), .c(s_181_17), .d(s_181_16), .cin(t_5190), .o(t_5217), .co(t_5218), .cout(t_5219));
compressor_4_2 u2_1776(.a(s_181_23), .b(s_181_22), .c(s_181_21), .d(s_181_20), .cin(t_5193), .o(t_5220), .co(t_5221), .cout(t_5222));
compressor_4_2 u2_1777(.a(s_181_27), .b(s_181_26), .c(s_181_25), .d(s_181_24), .cin(t_5196), .o(t_5223), .co(t_5224), .cout(t_5225));
compressor_4_2 u2_1778(.a(s_181_31), .b(s_181_30), .c(s_181_29), .d(s_181_28), .cin(t_5199), .o(t_5226), .co(t_5227), .cout(t_5228));
compressor_4_2 u2_1779(.a(s_181_35), .b(s_181_34), .c(s_181_33), .d(s_181_32), .cin(t_5202), .o(t_5229), .co(t_5230), .cout(t_5231));
compressor_3_2 u1_1780(.a(s_181_38), .b(s_181_37), .cin(s_181_36), .o(t_5232), .cout(t_5233));
compressor_4_2 u2_1781(.a(s_182_3), .b(s_182_2), .c(s_182_1), .d(s_182_0), .cin(t_5207), .o(t_5234), .co(t_5235), .cout(t_5236));
compressor_4_2 u2_1782(.a(s_182_7), .b(s_182_6), .c(s_182_5), .d(s_182_4), .cin(t_5210), .o(t_5237), .co(t_5238), .cout(t_5239));
compressor_4_2 u2_1783(.a(s_182_11), .b(s_182_10), .c(s_182_9), .d(s_182_8), .cin(t_5213), .o(t_5240), .co(t_5241), .cout(t_5242));
compressor_4_2 u2_1784(.a(s_182_15), .b(s_182_14), .c(s_182_13), .d(s_182_12), .cin(t_5216), .o(t_5243), .co(t_5244), .cout(t_5245));
compressor_4_2 u2_1785(.a(s_182_19), .b(s_182_18), .c(s_182_17), .d(s_182_16), .cin(t_5219), .o(t_5246), .co(t_5247), .cout(t_5248));
compressor_4_2 u2_1786(.a(s_182_23), .b(s_182_22), .c(s_182_21), .d(s_182_20), .cin(t_5222), .o(t_5249), .co(t_5250), .cout(t_5251));
compressor_4_2 u2_1787(.a(s_182_27), .b(s_182_26), .c(s_182_25), .d(s_182_24), .cin(t_5225), .o(t_5252), .co(t_5253), .cout(t_5254));
compressor_4_2 u2_1788(.a(s_182_31), .b(s_182_30), .c(s_182_29), .d(s_182_28), .cin(t_5228), .o(t_5255), .co(t_5256), .cout(t_5257));
compressor_4_2 u2_1789(.a(s_182_35), .b(s_182_34), .c(s_182_33), .d(s_182_32), .cin(t_5231), .o(t_5258), .co(t_5259), .cout(t_5260));
half_adder u0_1790(.a(s_182_37), .b(s_182_36), .o(t_5261), .cout(t_5262));
compressor_4_2 u2_1791(.a(s_183_3), .b(s_183_2), .c(s_183_1), .d(s_183_0), .cin(t_5236), .o(t_5263), .co(t_5264), .cout(t_5265));
compressor_4_2 u2_1792(.a(s_183_7), .b(s_183_6), .c(s_183_5), .d(s_183_4), .cin(t_5239), .o(t_5266), .co(t_5267), .cout(t_5268));
compressor_4_2 u2_1793(.a(s_183_11), .b(s_183_10), .c(s_183_9), .d(s_183_8), .cin(t_5242), .o(t_5269), .co(t_5270), .cout(t_5271));
compressor_4_2 u2_1794(.a(s_183_15), .b(s_183_14), .c(s_183_13), .d(s_183_12), .cin(t_5245), .o(t_5272), .co(t_5273), .cout(t_5274));
compressor_4_2 u2_1795(.a(s_183_19), .b(s_183_18), .c(s_183_17), .d(s_183_16), .cin(t_5248), .o(t_5275), .co(t_5276), .cout(t_5277));
compressor_4_2 u2_1796(.a(s_183_23), .b(s_183_22), .c(s_183_21), .d(s_183_20), .cin(t_5251), .o(t_5278), .co(t_5279), .cout(t_5280));
compressor_4_2 u2_1797(.a(s_183_27), .b(s_183_26), .c(s_183_25), .d(s_183_24), .cin(t_5254), .o(t_5281), .co(t_5282), .cout(t_5283));
compressor_4_2 u2_1798(.a(s_183_31), .b(s_183_30), .c(s_183_29), .d(s_183_28), .cin(t_5257), .o(t_5284), .co(t_5285), .cout(t_5286));
compressor_4_2 u2_1799(.a(s_183_35), .b(s_183_34), .c(s_183_33), .d(s_183_32), .cin(t_5260), .o(t_5287), .co(t_5288), .cout(t_5289));
half_adder u0_1800(.a(s_183_37), .b(s_183_36), .o(t_5290), .cout(t_5291));
compressor_4_2 u2_1801(.a(s_184_3), .b(s_184_2), .c(s_184_1), .d(s_184_0), .cin(t_5265), .o(t_5292), .co(t_5293), .cout(t_5294));
compressor_4_2 u2_1802(.a(s_184_7), .b(s_184_6), .c(s_184_5), .d(s_184_4), .cin(t_5268), .o(t_5295), .co(t_5296), .cout(t_5297));
compressor_4_2 u2_1803(.a(s_184_11), .b(s_184_10), .c(s_184_9), .d(s_184_8), .cin(t_5271), .o(t_5298), .co(t_5299), .cout(t_5300));
compressor_4_2 u2_1804(.a(s_184_15), .b(s_184_14), .c(s_184_13), .d(s_184_12), .cin(t_5274), .o(t_5301), .co(t_5302), .cout(t_5303));
compressor_4_2 u2_1805(.a(s_184_19), .b(s_184_18), .c(s_184_17), .d(s_184_16), .cin(t_5277), .o(t_5304), .co(t_5305), .cout(t_5306));
compressor_4_2 u2_1806(.a(s_184_23), .b(s_184_22), .c(s_184_21), .d(s_184_20), .cin(t_5280), .o(t_5307), .co(t_5308), .cout(t_5309));
compressor_4_2 u2_1807(.a(s_184_27), .b(s_184_26), .c(s_184_25), .d(s_184_24), .cin(t_5283), .o(t_5310), .co(t_5311), .cout(t_5312));
compressor_4_2 u2_1808(.a(s_184_31), .b(s_184_30), .c(s_184_29), .d(s_184_28), .cin(t_5286), .o(t_5313), .co(t_5314), .cout(t_5315));
compressor_4_2 u2_1809(.a(s_184_35), .b(s_184_34), .c(s_184_33), .d(s_184_32), .cin(t_5289), .o(t_5316), .co(t_5317), .cout(t_5318));
compressor_4_2 u2_1810(.a(s_185_3), .b(s_185_2), .c(s_185_1), .d(s_185_0), .cin(t_5294), .o(t_5319), .co(t_5320), .cout(t_5321));
compressor_4_2 u2_1811(.a(s_185_7), .b(s_185_6), .c(s_185_5), .d(s_185_4), .cin(t_5297), .o(t_5322), .co(t_5323), .cout(t_5324));
compressor_4_2 u2_1812(.a(s_185_11), .b(s_185_10), .c(s_185_9), .d(s_185_8), .cin(t_5300), .o(t_5325), .co(t_5326), .cout(t_5327));
compressor_4_2 u2_1813(.a(s_185_15), .b(s_185_14), .c(s_185_13), .d(s_185_12), .cin(t_5303), .o(t_5328), .co(t_5329), .cout(t_5330));
compressor_4_2 u2_1814(.a(s_185_19), .b(s_185_18), .c(s_185_17), .d(s_185_16), .cin(t_5306), .o(t_5331), .co(t_5332), .cout(t_5333));
compressor_4_2 u2_1815(.a(s_185_23), .b(s_185_22), .c(s_185_21), .d(s_185_20), .cin(t_5309), .o(t_5334), .co(t_5335), .cout(t_5336));
compressor_4_2 u2_1816(.a(s_185_27), .b(s_185_26), .c(s_185_25), .d(s_185_24), .cin(t_5312), .o(t_5337), .co(t_5338), .cout(t_5339));
compressor_4_2 u2_1817(.a(s_185_31), .b(s_185_30), .c(s_185_29), .d(s_185_28), .cin(t_5315), .o(t_5340), .co(t_5341), .cout(t_5342));
compressor_4_2 u2_1818(.a(s_185_35), .b(s_185_34), .c(s_185_33), .d(s_185_32), .cin(t_5318), .o(t_5343), .co(t_5344), .cout(t_5345));
compressor_4_2 u2_1819(.a(s_186_3), .b(s_186_2), .c(s_186_1), .d(s_186_0), .cin(t_5321), .o(t_5346), .co(t_5347), .cout(t_5348));
compressor_4_2 u2_1820(.a(s_186_7), .b(s_186_6), .c(s_186_5), .d(s_186_4), .cin(t_5324), .o(t_5349), .co(t_5350), .cout(t_5351));
compressor_4_2 u2_1821(.a(s_186_11), .b(s_186_10), .c(s_186_9), .d(s_186_8), .cin(t_5327), .o(t_5352), .co(t_5353), .cout(t_5354));
compressor_4_2 u2_1822(.a(s_186_15), .b(s_186_14), .c(s_186_13), .d(s_186_12), .cin(t_5330), .o(t_5355), .co(t_5356), .cout(t_5357));
compressor_4_2 u2_1823(.a(s_186_19), .b(s_186_18), .c(s_186_17), .d(s_186_16), .cin(t_5333), .o(t_5358), .co(t_5359), .cout(t_5360));
compressor_4_2 u2_1824(.a(s_186_23), .b(s_186_22), .c(s_186_21), .d(s_186_20), .cin(t_5336), .o(t_5361), .co(t_5362), .cout(t_5363));
compressor_4_2 u2_1825(.a(s_186_27), .b(s_186_26), .c(s_186_25), .d(s_186_24), .cin(t_5339), .o(t_5364), .co(t_5365), .cout(t_5366));
compressor_4_2 u2_1826(.a(s_186_31), .b(s_186_30), .c(s_186_29), .d(s_186_28), .cin(t_5342), .o(t_5367), .co(t_5368), .cout(t_5369));
compressor_4_2 u2_1827(.a(s_186_35), .b(s_186_34), .c(s_186_33), .d(s_186_32), .cin(t_5345), .o(t_5370), .co(t_5371), .cout(t_5372));
compressor_4_2 u2_1828(.a(s_187_3), .b(s_187_2), .c(s_187_1), .d(s_187_0), .cin(t_5348), .o(t_5373), .co(t_5374), .cout(t_5375));
compressor_4_2 u2_1829(.a(s_187_7), .b(s_187_6), .c(s_187_5), .d(s_187_4), .cin(t_5351), .o(t_5376), .co(t_5377), .cout(t_5378));
compressor_4_2 u2_1830(.a(s_187_11), .b(s_187_10), .c(s_187_9), .d(s_187_8), .cin(t_5354), .o(t_5379), .co(t_5380), .cout(t_5381));
compressor_4_2 u2_1831(.a(s_187_15), .b(s_187_14), .c(s_187_13), .d(s_187_12), .cin(t_5357), .o(t_5382), .co(t_5383), .cout(t_5384));
compressor_4_2 u2_1832(.a(s_187_19), .b(s_187_18), .c(s_187_17), .d(s_187_16), .cin(t_5360), .o(t_5385), .co(t_5386), .cout(t_5387));
compressor_4_2 u2_1833(.a(s_187_23), .b(s_187_22), .c(s_187_21), .d(s_187_20), .cin(t_5363), .o(t_5388), .co(t_5389), .cout(t_5390));
compressor_4_2 u2_1834(.a(s_187_27), .b(s_187_26), .c(s_187_25), .d(s_187_24), .cin(t_5366), .o(t_5391), .co(t_5392), .cout(t_5393));
compressor_4_2 u2_1835(.a(s_187_31), .b(s_187_30), .c(s_187_29), .d(s_187_28), .cin(t_5369), .o(t_5394), .co(t_5395), .cout(t_5396));
compressor_4_2 u2_1836(.a(s_187_35), .b(s_187_34), .c(s_187_33), .d(s_187_32), .cin(t_5372), .o(t_5397), .co(t_5398), .cout(t_5399));
compressor_4_2 u2_1837(.a(s_188_3), .b(s_188_2), .c(s_188_1), .d(s_188_0), .cin(t_5375), .o(t_5400), .co(t_5401), .cout(t_5402));
compressor_4_2 u2_1838(.a(s_188_7), .b(s_188_6), .c(s_188_5), .d(s_188_4), .cin(t_5378), .o(t_5403), .co(t_5404), .cout(t_5405));
compressor_4_2 u2_1839(.a(s_188_11), .b(s_188_10), .c(s_188_9), .d(s_188_8), .cin(t_5381), .o(t_5406), .co(t_5407), .cout(t_5408));
compressor_4_2 u2_1840(.a(s_188_15), .b(s_188_14), .c(s_188_13), .d(s_188_12), .cin(t_5384), .o(t_5409), .co(t_5410), .cout(t_5411));
compressor_4_2 u2_1841(.a(s_188_19), .b(s_188_18), .c(s_188_17), .d(s_188_16), .cin(t_5387), .o(t_5412), .co(t_5413), .cout(t_5414));
compressor_4_2 u2_1842(.a(s_188_23), .b(s_188_22), .c(s_188_21), .d(s_188_20), .cin(t_5390), .o(t_5415), .co(t_5416), .cout(t_5417));
compressor_4_2 u2_1843(.a(s_188_27), .b(s_188_26), .c(s_188_25), .d(s_188_24), .cin(t_5393), .o(t_5418), .co(t_5419), .cout(t_5420));
compressor_4_2 u2_1844(.a(s_188_31), .b(s_188_30), .c(s_188_29), .d(s_188_28), .cin(t_5396), .o(t_5421), .co(t_5422), .cout(t_5423));
compressor_3_2 u1_1845(.a(s_188_33), .b(s_188_32), .cin(t_5399), .o(t_5424), .cout(t_5425));
compressor_4_2 u2_1846(.a(s_189_3), .b(s_189_2), .c(s_189_1), .d(s_189_0), .cin(t_5402), .o(t_5426), .co(t_5427), .cout(t_5428));
compressor_4_2 u2_1847(.a(s_189_7), .b(s_189_6), .c(s_189_5), .d(s_189_4), .cin(t_5405), .o(t_5429), .co(t_5430), .cout(t_5431));
compressor_4_2 u2_1848(.a(s_189_11), .b(s_189_10), .c(s_189_9), .d(s_189_8), .cin(t_5408), .o(t_5432), .co(t_5433), .cout(t_5434));
compressor_4_2 u2_1849(.a(s_189_15), .b(s_189_14), .c(s_189_13), .d(s_189_12), .cin(t_5411), .o(t_5435), .co(t_5436), .cout(t_5437));
compressor_4_2 u2_1850(.a(s_189_19), .b(s_189_18), .c(s_189_17), .d(s_189_16), .cin(t_5414), .o(t_5438), .co(t_5439), .cout(t_5440));
compressor_4_2 u2_1851(.a(s_189_23), .b(s_189_22), .c(s_189_21), .d(s_189_20), .cin(t_5417), .o(t_5441), .co(t_5442), .cout(t_5443));
compressor_4_2 u2_1852(.a(s_189_27), .b(s_189_26), .c(s_189_25), .d(s_189_24), .cin(t_5420), .o(t_5444), .co(t_5445), .cout(t_5446));
compressor_4_2 u2_1853(.a(s_189_31), .b(s_189_30), .c(s_189_29), .d(s_189_28), .cin(t_5423), .o(t_5447), .co(t_5448), .cout(t_5449));
compressor_3_2 u1_1854(.a(s_189_34), .b(s_189_33), .cin(s_189_32), .o(t_5450), .cout(t_5451));
compressor_4_2 u2_1855(.a(s_190_3), .b(s_190_2), .c(s_190_1), .d(s_190_0), .cin(t_5428), .o(t_5452), .co(t_5453), .cout(t_5454));
compressor_4_2 u2_1856(.a(s_190_7), .b(s_190_6), .c(s_190_5), .d(s_190_4), .cin(t_5431), .o(t_5455), .co(t_5456), .cout(t_5457));
compressor_4_2 u2_1857(.a(s_190_11), .b(s_190_10), .c(s_190_9), .d(s_190_8), .cin(t_5434), .o(t_5458), .co(t_5459), .cout(t_5460));
compressor_4_2 u2_1858(.a(s_190_15), .b(s_190_14), .c(s_190_13), .d(s_190_12), .cin(t_5437), .o(t_5461), .co(t_5462), .cout(t_5463));
compressor_4_2 u2_1859(.a(s_190_19), .b(s_190_18), .c(s_190_17), .d(s_190_16), .cin(t_5440), .o(t_5464), .co(t_5465), .cout(t_5466));
compressor_4_2 u2_1860(.a(s_190_23), .b(s_190_22), .c(s_190_21), .d(s_190_20), .cin(t_5443), .o(t_5467), .co(t_5468), .cout(t_5469));
compressor_4_2 u2_1861(.a(s_190_27), .b(s_190_26), .c(s_190_25), .d(s_190_24), .cin(t_5446), .o(t_5470), .co(t_5471), .cout(t_5472));
compressor_4_2 u2_1862(.a(s_190_31), .b(s_190_30), .c(s_190_29), .d(s_190_28), .cin(t_5449), .o(t_5473), .co(t_5474), .cout(t_5475));
half_adder u0_1863(.a(s_190_33), .b(s_190_32), .o(t_5476), .cout(t_5477));
compressor_4_2 u2_1864(.a(s_191_3), .b(s_191_2), .c(s_191_1), .d(s_191_0), .cin(t_5454), .o(t_5478), .co(t_5479), .cout(t_5480));
compressor_4_2 u2_1865(.a(s_191_7), .b(s_191_6), .c(s_191_5), .d(s_191_4), .cin(t_5457), .o(t_5481), .co(t_5482), .cout(t_5483));
compressor_4_2 u2_1866(.a(s_191_11), .b(s_191_10), .c(s_191_9), .d(s_191_8), .cin(t_5460), .o(t_5484), .co(t_5485), .cout(t_5486));
compressor_4_2 u2_1867(.a(s_191_15), .b(s_191_14), .c(s_191_13), .d(s_191_12), .cin(t_5463), .o(t_5487), .co(t_5488), .cout(t_5489));
compressor_4_2 u2_1868(.a(s_191_19), .b(s_191_18), .c(s_191_17), .d(s_191_16), .cin(t_5466), .o(t_5490), .co(t_5491), .cout(t_5492));
compressor_4_2 u2_1869(.a(s_191_23), .b(s_191_22), .c(s_191_21), .d(s_191_20), .cin(t_5469), .o(t_5493), .co(t_5494), .cout(t_5495));
compressor_4_2 u2_1870(.a(s_191_27), .b(s_191_26), .c(s_191_25), .d(s_191_24), .cin(t_5472), .o(t_5496), .co(t_5497), .cout(t_5498));
compressor_4_2 u2_1871(.a(s_191_31), .b(s_191_30), .c(s_191_29), .d(s_191_28), .cin(t_5475), .o(t_5499), .co(t_5500), .cout(t_5501));
half_adder u0_1872(.a(s_191_33), .b(s_191_32), .o(t_5502), .cout(t_5503));
compressor_4_2 u2_1873(.a(s_192_3), .b(s_192_2), .c(s_192_1), .d(s_192_0), .cin(t_5480), .o(t_5504), .co(t_5505), .cout(t_5506));
compressor_4_2 u2_1874(.a(s_192_7), .b(s_192_6), .c(s_192_5), .d(s_192_4), .cin(t_5483), .o(t_5507), .co(t_5508), .cout(t_5509));
compressor_4_2 u2_1875(.a(s_192_11), .b(s_192_10), .c(s_192_9), .d(s_192_8), .cin(t_5486), .o(t_5510), .co(t_5511), .cout(t_5512));
compressor_4_2 u2_1876(.a(s_192_15), .b(s_192_14), .c(s_192_13), .d(s_192_12), .cin(t_5489), .o(t_5513), .co(t_5514), .cout(t_5515));
compressor_4_2 u2_1877(.a(s_192_19), .b(s_192_18), .c(s_192_17), .d(s_192_16), .cin(t_5492), .o(t_5516), .co(t_5517), .cout(t_5518));
compressor_4_2 u2_1878(.a(s_192_23), .b(s_192_22), .c(s_192_21), .d(s_192_20), .cin(t_5495), .o(t_5519), .co(t_5520), .cout(t_5521));
compressor_4_2 u2_1879(.a(s_192_27), .b(s_192_26), .c(s_192_25), .d(s_192_24), .cin(t_5498), .o(t_5522), .co(t_5523), .cout(t_5524));
compressor_4_2 u2_1880(.a(s_192_31), .b(s_192_30), .c(s_192_29), .d(s_192_28), .cin(t_5501), .o(t_5525), .co(t_5526), .cout(t_5527));
compressor_4_2 u2_1881(.a(s_193_3), .b(s_193_2), .c(s_193_1), .d(s_193_0), .cin(t_5506), .o(t_5528), .co(t_5529), .cout(t_5530));
compressor_4_2 u2_1882(.a(s_193_7), .b(s_193_6), .c(s_193_5), .d(s_193_4), .cin(t_5509), .o(t_5531), .co(t_5532), .cout(t_5533));
compressor_4_2 u2_1883(.a(s_193_11), .b(s_193_10), .c(s_193_9), .d(s_193_8), .cin(t_5512), .o(t_5534), .co(t_5535), .cout(t_5536));
compressor_4_2 u2_1884(.a(s_193_15), .b(s_193_14), .c(s_193_13), .d(s_193_12), .cin(t_5515), .o(t_5537), .co(t_5538), .cout(t_5539));
compressor_4_2 u2_1885(.a(s_193_19), .b(s_193_18), .c(s_193_17), .d(s_193_16), .cin(t_5518), .o(t_5540), .co(t_5541), .cout(t_5542));
compressor_4_2 u2_1886(.a(s_193_23), .b(s_193_22), .c(s_193_21), .d(s_193_20), .cin(t_5521), .o(t_5543), .co(t_5544), .cout(t_5545));
compressor_4_2 u2_1887(.a(s_193_27), .b(s_193_26), .c(s_193_25), .d(s_193_24), .cin(t_5524), .o(t_5546), .co(t_5547), .cout(t_5548));
compressor_4_2 u2_1888(.a(s_193_31), .b(s_193_30), .c(s_193_29), .d(s_193_28), .cin(t_5527), .o(t_5549), .co(t_5550), .cout(t_5551));
compressor_4_2 u2_1889(.a(s_194_3), .b(s_194_2), .c(s_194_1), .d(s_194_0), .cin(t_5530), .o(t_5552), .co(t_5553), .cout(t_5554));
compressor_4_2 u2_1890(.a(s_194_7), .b(s_194_6), .c(s_194_5), .d(s_194_4), .cin(t_5533), .o(t_5555), .co(t_5556), .cout(t_5557));
compressor_4_2 u2_1891(.a(s_194_11), .b(s_194_10), .c(s_194_9), .d(s_194_8), .cin(t_5536), .o(t_5558), .co(t_5559), .cout(t_5560));
compressor_4_2 u2_1892(.a(s_194_15), .b(s_194_14), .c(s_194_13), .d(s_194_12), .cin(t_5539), .o(t_5561), .co(t_5562), .cout(t_5563));
compressor_4_2 u2_1893(.a(s_194_19), .b(s_194_18), .c(s_194_17), .d(s_194_16), .cin(t_5542), .o(t_5564), .co(t_5565), .cout(t_5566));
compressor_4_2 u2_1894(.a(s_194_23), .b(s_194_22), .c(s_194_21), .d(s_194_20), .cin(t_5545), .o(t_5567), .co(t_5568), .cout(t_5569));
compressor_4_2 u2_1895(.a(s_194_27), .b(s_194_26), .c(s_194_25), .d(s_194_24), .cin(t_5548), .o(t_5570), .co(t_5571), .cout(t_5572));
compressor_4_2 u2_1896(.a(s_194_31), .b(s_194_30), .c(s_194_29), .d(s_194_28), .cin(t_5551), .o(t_5573), .co(t_5574), .cout(t_5575));
compressor_4_2 u2_1897(.a(s_195_3), .b(s_195_2), .c(s_195_1), .d(s_195_0), .cin(t_5554), .o(t_5576), .co(t_5577), .cout(t_5578));
compressor_4_2 u2_1898(.a(s_195_7), .b(s_195_6), .c(s_195_5), .d(s_195_4), .cin(t_5557), .o(t_5579), .co(t_5580), .cout(t_5581));
compressor_4_2 u2_1899(.a(s_195_11), .b(s_195_10), .c(s_195_9), .d(s_195_8), .cin(t_5560), .o(t_5582), .co(t_5583), .cout(t_5584));
compressor_4_2 u2_1900(.a(s_195_15), .b(s_195_14), .c(s_195_13), .d(s_195_12), .cin(t_5563), .o(t_5585), .co(t_5586), .cout(t_5587));
compressor_4_2 u2_1901(.a(s_195_19), .b(s_195_18), .c(s_195_17), .d(s_195_16), .cin(t_5566), .o(t_5588), .co(t_5589), .cout(t_5590));
compressor_4_2 u2_1902(.a(s_195_23), .b(s_195_22), .c(s_195_21), .d(s_195_20), .cin(t_5569), .o(t_5591), .co(t_5592), .cout(t_5593));
compressor_4_2 u2_1903(.a(s_195_27), .b(s_195_26), .c(s_195_25), .d(s_195_24), .cin(t_5572), .o(t_5594), .co(t_5595), .cout(t_5596));
compressor_4_2 u2_1904(.a(s_195_31), .b(s_195_30), .c(s_195_29), .d(s_195_28), .cin(t_5575), .o(t_5597), .co(t_5598), .cout(t_5599));
compressor_4_2 u2_1905(.a(s_196_3), .b(s_196_2), .c(s_196_1), .d(s_196_0), .cin(t_5578), .o(t_5600), .co(t_5601), .cout(t_5602));
compressor_4_2 u2_1906(.a(s_196_7), .b(s_196_6), .c(s_196_5), .d(s_196_4), .cin(t_5581), .o(t_5603), .co(t_5604), .cout(t_5605));
compressor_4_2 u2_1907(.a(s_196_11), .b(s_196_10), .c(s_196_9), .d(s_196_8), .cin(t_5584), .o(t_5606), .co(t_5607), .cout(t_5608));
compressor_4_2 u2_1908(.a(s_196_15), .b(s_196_14), .c(s_196_13), .d(s_196_12), .cin(t_5587), .o(t_5609), .co(t_5610), .cout(t_5611));
compressor_4_2 u2_1909(.a(s_196_19), .b(s_196_18), .c(s_196_17), .d(s_196_16), .cin(t_5590), .o(t_5612), .co(t_5613), .cout(t_5614));
compressor_4_2 u2_1910(.a(s_196_23), .b(s_196_22), .c(s_196_21), .d(s_196_20), .cin(t_5593), .o(t_5615), .co(t_5616), .cout(t_5617));
compressor_4_2 u2_1911(.a(s_196_27), .b(s_196_26), .c(s_196_25), .d(s_196_24), .cin(t_5596), .o(t_5618), .co(t_5619), .cout(t_5620));
compressor_3_2 u1_1912(.a(s_196_29), .b(s_196_28), .cin(t_5599), .o(t_5621), .cout(t_5622));
compressor_4_2 u2_1913(.a(s_197_3), .b(s_197_2), .c(s_197_1), .d(s_197_0), .cin(t_5602), .o(t_5623), .co(t_5624), .cout(t_5625));
compressor_4_2 u2_1914(.a(s_197_7), .b(s_197_6), .c(s_197_5), .d(s_197_4), .cin(t_5605), .o(t_5626), .co(t_5627), .cout(t_5628));
compressor_4_2 u2_1915(.a(s_197_11), .b(s_197_10), .c(s_197_9), .d(s_197_8), .cin(t_5608), .o(t_5629), .co(t_5630), .cout(t_5631));
compressor_4_2 u2_1916(.a(s_197_15), .b(s_197_14), .c(s_197_13), .d(s_197_12), .cin(t_5611), .o(t_5632), .co(t_5633), .cout(t_5634));
compressor_4_2 u2_1917(.a(s_197_19), .b(s_197_18), .c(s_197_17), .d(s_197_16), .cin(t_5614), .o(t_5635), .co(t_5636), .cout(t_5637));
compressor_4_2 u2_1918(.a(s_197_23), .b(s_197_22), .c(s_197_21), .d(s_197_20), .cin(t_5617), .o(t_5638), .co(t_5639), .cout(t_5640));
compressor_4_2 u2_1919(.a(s_197_27), .b(s_197_26), .c(s_197_25), .d(s_197_24), .cin(t_5620), .o(t_5641), .co(t_5642), .cout(t_5643));
compressor_3_2 u1_1920(.a(s_197_30), .b(s_197_29), .cin(s_197_28), .o(t_5644), .cout(t_5645));
compressor_4_2 u2_1921(.a(s_198_3), .b(s_198_2), .c(s_198_1), .d(s_198_0), .cin(t_5625), .o(t_5646), .co(t_5647), .cout(t_5648));
compressor_4_2 u2_1922(.a(s_198_7), .b(s_198_6), .c(s_198_5), .d(s_198_4), .cin(t_5628), .o(t_5649), .co(t_5650), .cout(t_5651));
compressor_4_2 u2_1923(.a(s_198_11), .b(s_198_10), .c(s_198_9), .d(s_198_8), .cin(t_5631), .o(t_5652), .co(t_5653), .cout(t_5654));
compressor_4_2 u2_1924(.a(s_198_15), .b(s_198_14), .c(s_198_13), .d(s_198_12), .cin(t_5634), .o(t_5655), .co(t_5656), .cout(t_5657));
compressor_4_2 u2_1925(.a(s_198_19), .b(s_198_18), .c(s_198_17), .d(s_198_16), .cin(t_5637), .o(t_5658), .co(t_5659), .cout(t_5660));
compressor_4_2 u2_1926(.a(s_198_23), .b(s_198_22), .c(s_198_21), .d(s_198_20), .cin(t_5640), .o(t_5661), .co(t_5662), .cout(t_5663));
compressor_4_2 u2_1927(.a(s_198_27), .b(s_198_26), .c(s_198_25), .d(s_198_24), .cin(t_5643), .o(t_5664), .co(t_5665), .cout(t_5666));
half_adder u0_1928(.a(s_198_29), .b(s_198_28), .o(t_5667), .cout(t_5668));
compressor_4_2 u2_1929(.a(s_199_3), .b(s_199_2), .c(s_199_1), .d(s_199_0), .cin(t_5648), .o(t_5669), .co(t_5670), .cout(t_5671));
compressor_4_2 u2_1930(.a(s_199_7), .b(s_199_6), .c(s_199_5), .d(s_199_4), .cin(t_5651), .o(t_5672), .co(t_5673), .cout(t_5674));
compressor_4_2 u2_1931(.a(s_199_11), .b(s_199_10), .c(s_199_9), .d(s_199_8), .cin(t_5654), .o(t_5675), .co(t_5676), .cout(t_5677));
compressor_4_2 u2_1932(.a(s_199_15), .b(s_199_14), .c(s_199_13), .d(s_199_12), .cin(t_5657), .o(t_5678), .co(t_5679), .cout(t_5680));
compressor_4_2 u2_1933(.a(s_199_19), .b(s_199_18), .c(s_199_17), .d(s_199_16), .cin(t_5660), .o(t_5681), .co(t_5682), .cout(t_5683));
compressor_4_2 u2_1934(.a(s_199_23), .b(s_199_22), .c(s_199_21), .d(s_199_20), .cin(t_5663), .o(t_5684), .co(t_5685), .cout(t_5686));
compressor_4_2 u2_1935(.a(s_199_27), .b(s_199_26), .c(s_199_25), .d(s_199_24), .cin(t_5666), .o(t_5687), .co(t_5688), .cout(t_5689));
half_adder u0_1936(.a(s_199_29), .b(s_199_28), .o(t_5690), .cout(t_5691));
compressor_4_2 u2_1937(.a(s_200_3), .b(s_200_2), .c(s_200_1), .d(s_200_0), .cin(t_5671), .o(t_5692), .co(t_5693), .cout(t_5694));
compressor_4_2 u2_1938(.a(s_200_7), .b(s_200_6), .c(s_200_5), .d(s_200_4), .cin(t_5674), .o(t_5695), .co(t_5696), .cout(t_5697));
compressor_4_2 u2_1939(.a(s_200_11), .b(s_200_10), .c(s_200_9), .d(s_200_8), .cin(t_5677), .o(t_5698), .co(t_5699), .cout(t_5700));
compressor_4_2 u2_1940(.a(s_200_15), .b(s_200_14), .c(s_200_13), .d(s_200_12), .cin(t_5680), .o(t_5701), .co(t_5702), .cout(t_5703));
compressor_4_2 u2_1941(.a(s_200_19), .b(s_200_18), .c(s_200_17), .d(s_200_16), .cin(t_5683), .o(t_5704), .co(t_5705), .cout(t_5706));
compressor_4_2 u2_1942(.a(s_200_23), .b(s_200_22), .c(s_200_21), .d(s_200_20), .cin(t_5686), .o(t_5707), .co(t_5708), .cout(t_5709));
compressor_4_2 u2_1943(.a(s_200_27), .b(s_200_26), .c(s_200_25), .d(s_200_24), .cin(t_5689), .o(t_5710), .co(t_5711), .cout(t_5712));
compressor_4_2 u2_1944(.a(s_201_3), .b(s_201_2), .c(s_201_1), .d(s_201_0), .cin(t_5694), .o(t_5713), .co(t_5714), .cout(t_5715));
compressor_4_2 u2_1945(.a(s_201_7), .b(s_201_6), .c(s_201_5), .d(s_201_4), .cin(t_5697), .o(t_5716), .co(t_5717), .cout(t_5718));
compressor_4_2 u2_1946(.a(s_201_11), .b(s_201_10), .c(s_201_9), .d(s_201_8), .cin(t_5700), .o(t_5719), .co(t_5720), .cout(t_5721));
compressor_4_2 u2_1947(.a(s_201_15), .b(s_201_14), .c(s_201_13), .d(s_201_12), .cin(t_5703), .o(t_5722), .co(t_5723), .cout(t_5724));
compressor_4_2 u2_1948(.a(s_201_19), .b(s_201_18), .c(s_201_17), .d(s_201_16), .cin(t_5706), .o(t_5725), .co(t_5726), .cout(t_5727));
compressor_4_2 u2_1949(.a(s_201_23), .b(s_201_22), .c(s_201_21), .d(s_201_20), .cin(t_5709), .o(t_5728), .co(t_5729), .cout(t_5730));
compressor_4_2 u2_1950(.a(s_201_27), .b(s_201_26), .c(s_201_25), .d(s_201_24), .cin(t_5712), .o(t_5731), .co(t_5732), .cout(t_5733));
compressor_4_2 u2_1951(.a(s_202_3), .b(s_202_2), .c(s_202_1), .d(s_202_0), .cin(t_5715), .o(t_5734), .co(t_5735), .cout(t_5736));
compressor_4_2 u2_1952(.a(s_202_7), .b(s_202_6), .c(s_202_5), .d(s_202_4), .cin(t_5718), .o(t_5737), .co(t_5738), .cout(t_5739));
compressor_4_2 u2_1953(.a(s_202_11), .b(s_202_10), .c(s_202_9), .d(s_202_8), .cin(t_5721), .o(t_5740), .co(t_5741), .cout(t_5742));
compressor_4_2 u2_1954(.a(s_202_15), .b(s_202_14), .c(s_202_13), .d(s_202_12), .cin(t_5724), .o(t_5743), .co(t_5744), .cout(t_5745));
compressor_4_2 u2_1955(.a(s_202_19), .b(s_202_18), .c(s_202_17), .d(s_202_16), .cin(t_5727), .o(t_5746), .co(t_5747), .cout(t_5748));
compressor_4_2 u2_1956(.a(s_202_23), .b(s_202_22), .c(s_202_21), .d(s_202_20), .cin(t_5730), .o(t_5749), .co(t_5750), .cout(t_5751));
compressor_4_2 u2_1957(.a(s_202_27), .b(s_202_26), .c(s_202_25), .d(s_202_24), .cin(t_5733), .o(t_5752), .co(t_5753), .cout(t_5754));
compressor_4_2 u2_1958(.a(s_203_3), .b(s_203_2), .c(s_203_1), .d(s_203_0), .cin(t_5736), .o(t_5755), .co(t_5756), .cout(t_5757));
compressor_4_2 u2_1959(.a(s_203_7), .b(s_203_6), .c(s_203_5), .d(s_203_4), .cin(t_5739), .o(t_5758), .co(t_5759), .cout(t_5760));
compressor_4_2 u2_1960(.a(s_203_11), .b(s_203_10), .c(s_203_9), .d(s_203_8), .cin(t_5742), .o(t_5761), .co(t_5762), .cout(t_5763));
compressor_4_2 u2_1961(.a(s_203_15), .b(s_203_14), .c(s_203_13), .d(s_203_12), .cin(t_5745), .o(t_5764), .co(t_5765), .cout(t_5766));
compressor_4_2 u2_1962(.a(s_203_19), .b(s_203_18), .c(s_203_17), .d(s_203_16), .cin(t_5748), .o(t_5767), .co(t_5768), .cout(t_5769));
compressor_4_2 u2_1963(.a(s_203_23), .b(s_203_22), .c(s_203_21), .d(s_203_20), .cin(t_5751), .o(t_5770), .co(t_5771), .cout(t_5772));
compressor_4_2 u2_1964(.a(s_203_27), .b(s_203_26), .c(s_203_25), .d(s_203_24), .cin(t_5754), .o(t_5773), .co(t_5774), .cout(t_5775));
compressor_4_2 u2_1965(.a(s_204_3), .b(s_204_2), .c(s_204_1), .d(s_204_0), .cin(t_5757), .o(t_5776), .co(t_5777), .cout(t_5778));
compressor_4_2 u2_1966(.a(s_204_7), .b(s_204_6), .c(s_204_5), .d(s_204_4), .cin(t_5760), .o(t_5779), .co(t_5780), .cout(t_5781));
compressor_4_2 u2_1967(.a(s_204_11), .b(s_204_10), .c(s_204_9), .d(s_204_8), .cin(t_5763), .o(t_5782), .co(t_5783), .cout(t_5784));
compressor_4_2 u2_1968(.a(s_204_15), .b(s_204_14), .c(s_204_13), .d(s_204_12), .cin(t_5766), .o(t_5785), .co(t_5786), .cout(t_5787));
compressor_4_2 u2_1969(.a(s_204_19), .b(s_204_18), .c(s_204_17), .d(s_204_16), .cin(t_5769), .o(t_5788), .co(t_5789), .cout(t_5790));
compressor_4_2 u2_1970(.a(s_204_23), .b(s_204_22), .c(s_204_21), .d(s_204_20), .cin(t_5772), .o(t_5791), .co(t_5792), .cout(t_5793));
compressor_3_2 u1_1971(.a(s_204_25), .b(s_204_24), .cin(t_5775), .o(t_5794), .cout(t_5795));
compressor_4_2 u2_1972(.a(s_205_3), .b(s_205_2), .c(s_205_1), .d(s_205_0), .cin(t_5778), .o(t_5796), .co(t_5797), .cout(t_5798));
compressor_4_2 u2_1973(.a(s_205_7), .b(s_205_6), .c(s_205_5), .d(s_205_4), .cin(t_5781), .o(t_5799), .co(t_5800), .cout(t_5801));
compressor_4_2 u2_1974(.a(s_205_11), .b(s_205_10), .c(s_205_9), .d(s_205_8), .cin(t_5784), .o(t_5802), .co(t_5803), .cout(t_5804));
compressor_4_2 u2_1975(.a(s_205_15), .b(s_205_14), .c(s_205_13), .d(s_205_12), .cin(t_5787), .o(t_5805), .co(t_5806), .cout(t_5807));
compressor_4_2 u2_1976(.a(s_205_19), .b(s_205_18), .c(s_205_17), .d(s_205_16), .cin(t_5790), .o(t_5808), .co(t_5809), .cout(t_5810));
compressor_4_2 u2_1977(.a(s_205_23), .b(s_205_22), .c(s_205_21), .d(s_205_20), .cin(t_5793), .o(t_5811), .co(t_5812), .cout(t_5813));
compressor_3_2 u1_1978(.a(s_205_26), .b(s_205_25), .cin(s_205_24), .o(t_5814), .cout(t_5815));
compressor_4_2 u2_1979(.a(s_206_3), .b(s_206_2), .c(s_206_1), .d(s_206_0), .cin(t_5798), .o(t_5816), .co(t_5817), .cout(t_5818));
compressor_4_2 u2_1980(.a(s_206_7), .b(s_206_6), .c(s_206_5), .d(s_206_4), .cin(t_5801), .o(t_5819), .co(t_5820), .cout(t_5821));
compressor_4_2 u2_1981(.a(s_206_11), .b(s_206_10), .c(s_206_9), .d(s_206_8), .cin(t_5804), .o(t_5822), .co(t_5823), .cout(t_5824));
compressor_4_2 u2_1982(.a(s_206_15), .b(s_206_14), .c(s_206_13), .d(s_206_12), .cin(t_5807), .o(t_5825), .co(t_5826), .cout(t_5827));
compressor_4_2 u2_1983(.a(s_206_19), .b(s_206_18), .c(s_206_17), .d(s_206_16), .cin(t_5810), .o(t_5828), .co(t_5829), .cout(t_5830));
compressor_4_2 u2_1984(.a(s_206_23), .b(s_206_22), .c(s_206_21), .d(s_206_20), .cin(t_5813), .o(t_5831), .co(t_5832), .cout(t_5833));
half_adder u0_1985(.a(s_206_25), .b(s_206_24), .o(t_5834), .cout(t_5835));
compressor_4_2 u2_1986(.a(s_207_3), .b(s_207_2), .c(s_207_1), .d(s_207_0), .cin(t_5818), .o(t_5836), .co(t_5837), .cout(t_5838));
compressor_4_2 u2_1987(.a(s_207_7), .b(s_207_6), .c(s_207_5), .d(s_207_4), .cin(t_5821), .o(t_5839), .co(t_5840), .cout(t_5841));
compressor_4_2 u2_1988(.a(s_207_11), .b(s_207_10), .c(s_207_9), .d(s_207_8), .cin(t_5824), .o(t_5842), .co(t_5843), .cout(t_5844));
compressor_4_2 u2_1989(.a(s_207_15), .b(s_207_14), .c(s_207_13), .d(s_207_12), .cin(t_5827), .o(t_5845), .co(t_5846), .cout(t_5847));
compressor_4_2 u2_1990(.a(s_207_19), .b(s_207_18), .c(s_207_17), .d(s_207_16), .cin(t_5830), .o(t_5848), .co(t_5849), .cout(t_5850));
compressor_4_2 u2_1991(.a(s_207_23), .b(s_207_22), .c(s_207_21), .d(s_207_20), .cin(t_5833), .o(t_5851), .co(t_5852), .cout(t_5853));
half_adder u0_1992(.a(s_207_25), .b(s_207_24), .o(t_5854), .cout(t_5855));
compressor_4_2 u2_1993(.a(s_208_3), .b(s_208_2), .c(s_208_1), .d(s_208_0), .cin(t_5838), .o(t_5856), .co(t_5857), .cout(t_5858));
compressor_4_2 u2_1994(.a(s_208_7), .b(s_208_6), .c(s_208_5), .d(s_208_4), .cin(t_5841), .o(t_5859), .co(t_5860), .cout(t_5861));
compressor_4_2 u2_1995(.a(s_208_11), .b(s_208_10), .c(s_208_9), .d(s_208_8), .cin(t_5844), .o(t_5862), .co(t_5863), .cout(t_5864));
compressor_4_2 u2_1996(.a(s_208_15), .b(s_208_14), .c(s_208_13), .d(s_208_12), .cin(t_5847), .o(t_5865), .co(t_5866), .cout(t_5867));
compressor_4_2 u2_1997(.a(s_208_19), .b(s_208_18), .c(s_208_17), .d(s_208_16), .cin(t_5850), .o(t_5868), .co(t_5869), .cout(t_5870));
compressor_4_2 u2_1998(.a(s_208_23), .b(s_208_22), .c(s_208_21), .d(s_208_20), .cin(t_5853), .o(t_5871), .co(t_5872), .cout(t_5873));
compressor_4_2 u2_1999(.a(s_209_3), .b(s_209_2), .c(s_209_1), .d(s_209_0), .cin(t_5858), .o(t_5874), .co(t_5875), .cout(t_5876));
compressor_4_2 u2_2000(.a(s_209_7), .b(s_209_6), .c(s_209_5), .d(s_209_4), .cin(t_5861), .o(t_5877), .co(t_5878), .cout(t_5879));
compressor_4_2 u2_2001(.a(s_209_11), .b(s_209_10), .c(s_209_9), .d(s_209_8), .cin(t_5864), .o(t_5880), .co(t_5881), .cout(t_5882));
compressor_4_2 u2_2002(.a(s_209_15), .b(s_209_14), .c(s_209_13), .d(s_209_12), .cin(t_5867), .o(t_5883), .co(t_5884), .cout(t_5885));
compressor_4_2 u2_2003(.a(s_209_19), .b(s_209_18), .c(s_209_17), .d(s_209_16), .cin(t_5870), .o(t_5886), .co(t_5887), .cout(t_5888));
compressor_4_2 u2_2004(.a(s_209_23), .b(s_209_22), .c(s_209_21), .d(s_209_20), .cin(t_5873), .o(t_5889), .co(t_5890), .cout(t_5891));
compressor_4_2 u2_2005(.a(s_210_3), .b(s_210_2), .c(s_210_1), .d(s_210_0), .cin(t_5876), .o(t_5892), .co(t_5893), .cout(t_5894));
compressor_4_2 u2_2006(.a(s_210_7), .b(s_210_6), .c(s_210_5), .d(s_210_4), .cin(t_5879), .o(t_5895), .co(t_5896), .cout(t_5897));
compressor_4_2 u2_2007(.a(s_210_11), .b(s_210_10), .c(s_210_9), .d(s_210_8), .cin(t_5882), .o(t_5898), .co(t_5899), .cout(t_5900));
compressor_4_2 u2_2008(.a(s_210_15), .b(s_210_14), .c(s_210_13), .d(s_210_12), .cin(t_5885), .o(t_5901), .co(t_5902), .cout(t_5903));
compressor_4_2 u2_2009(.a(s_210_19), .b(s_210_18), .c(s_210_17), .d(s_210_16), .cin(t_5888), .o(t_5904), .co(t_5905), .cout(t_5906));
compressor_4_2 u2_2010(.a(s_210_23), .b(s_210_22), .c(s_210_21), .d(s_210_20), .cin(t_5891), .o(t_5907), .co(t_5908), .cout(t_5909));
compressor_4_2 u2_2011(.a(s_211_3), .b(s_211_2), .c(s_211_1), .d(s_211_0), .cin(t_5894), .o(t_5910), .co(t_5911), .cout(t_5912));
compressor_4_2 u2_2012(.a(s_211_7), .b(s_211_6), .c(s_211_5), .d(s_211_4), .cin(t_5897), .o(t_5913), .co(t_5914), .cout(t_5915));
compressor_4_2 u2_2013(.a(s_211_11), .b(s_211_10), .c(s_211_9), .d(s_211_8), .cin(t_5900), .o(t_5916), .co(t_5917), .cout(t_5918));
compressor_4_2 u2_2014(.a(s_211_15), .b(s_211_14), .c(s_211_13), .d(s_211_12), .cin(t_5903), .o(t_5919), .co(t_5920), .cout(t_5921));
compressor_4_2 u2_2015(.a(s_211_19), .b(s_211_18), .c(s_211_17), .d(s_211_16), .cin(t_5906), .o(t_5922), .co(t_5923), .cout(t_5924));
compressor_4_2 u2_2016(.a(s_211_23), .b(s_211_22), .c(s_211_21), .d(s_211_20), .cin(t_5909), .o(t_5925), .co(t_5926), .cout(t_5927));
compressor_4_2 u2_2017(.a(s_212_3), .b(s_212_2), .c(s_212_1), .d(s_212_0), .cin(t_5912), .o(t_5928), .co(t_5929), .cout(t_5930));
compressor_4_2 u2_2018(.a(s_212_7), .b(s_212_6), .c(s_212_5), .d(s_212_4), .cin(t_5915), .o(t_5931), .co(t_5932), .cout(t_5933));
compressor_4_2 u2_2019(.a(s_212_11), .b(s_212_10), .c(s_212_9), .d(s_212_8), .cin(t_5918), .o(t_5934), .co(t_5935), .cout(t_5936));
compressor_4_2 u2_2020(.a(s_212_15), .b(s_212_14), .c(s_212_13), .d(s_212_12), .cin(t_5921), .o(t_5937), .co(t_5938), .cout(t_5939));
compressor_4_2 u2_2021(.a(s_212_19), .b(s_212_18), .c(s_212_17), .d(s_212_16), .cin(t_5924), .o(t_5940), .co(t_5941), .cout(t_5942));
compressor_3_2 u1_2022(.a(s_212_21), .b(s_212_20), .cin(t_5927), .o(t_5943), .cout(t_5944));
compressor_4_2 u2_2023(.a(s_213_3), .b(s_213_2), .c(s_213_1), .d(s_213_0), .cin(t_5930), .o(t_5945), .co(t_5946), .cout(t_5947));
compressor_4_2 u2_2024(.a(s_213_7), .b(s_213_6), .c(s_213_5), .d(s_213_4), .cin(t_5933), .o(t_5948), .co(t_5949), .cout(t_5950));
compressor_4_2 u2_2025(.a(s_213_11), .b(s_213_10), .c(s_213_9), .d(s_213_8), .cin(t_5936), .o(t_5951), .co(t_5952), .cout(t_5953));
compressor_4_2 u2_2026(.a(s_213_15), .b(s_213_14), .c(s_213_13), .d(s_213_12), .cin(t_5939), .o(t_5954), .co(t_5955), .cout(t_5956));
compressor_4_2 u2_2027(.a(s_213_19), .b(s_213_18), .c(s_213_17), .d(s_213_16), .cin(t_5942), .o(t_5957), .co(t_5958), .cout(t_5959));
compressor_3_2 u1_2028(.a(s_213_22), .b(s_213_21), .cin(s_213_20), .o(t_5960), .cout(t_5961));
compressor_4_2 u2_2029(.a(s_214_3), .b(s_214_2), .c(s_214_1), .d(s_214_0), .cin(t_5947), .o(t_5962), .co(t_5963), .cout(t_5964));
compressor_4_2 u2_2030(.a(s_214_7), .b(s_214_6), .c(s_214_5), .d(s_214_4), .cin(t_5950), .o(t_5965), .co(t_5966), .cout(t_5967));
compressor_4_2 u2_2031(.a(s_214_11), .b(s_214_10), .c(s_214_9), .d(s_214_8), .cin(t_5953), .o(t_5968), .co(t_5969), .cout(t_5970));
compressor_4_2 u2_2032(.a(s_214_15), .b(s_214_14), .c(s_214_13), .d(s_214_12), .cin(t_5956), .o(t_5971), .co(t_5972), .cout(t_5973));
compressor_4_2 u2_2033(.a(s_214_19), .b(s_214_18), .c(s_214_17), .d(s_214_16), .cin(t_5959), .o(t_5974), .co(t_5975), .cout(t_5976));
half_adder u0_2034(.a(s_214_21), .b(s_214_20), .o(t_5977), .cout(t_5978));
compressor_4_2 u2_2035(.a(s_215_3), .b(s_215_2), .c(s_215_1), .d(s_215_0), .cin(t_5964), .o(t_5979), .co(t_5980), .cout(t_5981));
compressor_4_2 u2_2036(.a(s_215_7), .b(s_215_6), .c(s_215_5), .d(s_215_4), .cin(t_5967), .o(t_5982), .co(t_5983), .cout(t_5984));
compressor_4_2 u2_2037(.a(s_215_11), .b(s_215_10), .c(s_215_9), .d(s_215_8), .cin(t_5970), .o(t_5985), .co(t_5986), .cout(t_5987));
compressor_4_2 u2_2038(.a(s_215_15), .b(s_215_14), .c(s_215_13), .d(s_215_12), .cin(t_5973), .o(t_5988), .co(t_5989), .cout(t_5990));
compressor_4_2 u2_2039(.a(s_215_19), .b(s_215_18), .c(s_215_17), .d(s_215_16), .cin(t_5976), .o(t_5991), .co(t_5992), .cout(t_5993));
half_adder u0_2040(.a(s_215_21), .b(s_215_20), .o(t_5994), .cout(t_5995));
compressor_4_2 u2_2041(.a(s_216_3), .b(s_216_2), .c(s_216_1), .d(s_216_0), .cin(t_5981), .o(t_5996), .co(t_5997), .cout(t_5998));
compressor_4_2 u2_2042(.a(s_216_7), .b(s_216_6), .c(s_216_5), .d(s_216_4), .cin(t_5984), .o(t_5999), .co(t_6000), .cout(t_6001));
compressor_4_2 u2_2043(.a(s_216_11), .b(s_216_10), .c(s_216_9), .d(s_216_8), .cin(t_5987), .o(t_6002), .co(t_6003), .cout(t_6004));
compressor_4_2 u2_2044(.a(s_216_15), .b(s_216_14), .c(s_216_13), .d(s_216_12), .cin(t_5990), .o(t_6005), .co(t_6006), .cout(t_6007));
compressor_4_2 u2_2045(.a(s_216_19), .b(s_216_18), .c(s_216_17), .d(s_216_16), .cin(t_5993), .o(t_6008), .co(t_6009), .cout(t_6010));
compressor_4_2 u2_2046(.a(s_217_3), .b(s_217_2), .c(s_217_1), .d(s_217_0), .cin(t_5998), .o(t_6011), .co(t_6012), .cout(t_6013));
compressor_4_2 u2_2047(.a(s_217_7), .b(s_217_6), .c(s_217_5), .d(s_217_4), .cin(t_6001), .o(t_6014), .co(t_6015), .cout(t_6016));
compressor_4_2 u2_2048(.a(s_217_11), .b(s_217_10), .c(s_217_9), .d(s_217_8), .cin(t_6004), .o(t_6017), .co(t_6018), .cout(t_6019));
compressor_4_2 u2_2049(.a(s_217_15), .b(s_217_14), .c(s_217_13), .d(s_217_12), .cin(t_6007), .o(t_6020), .co(t_6021), .cout(t_6022));
compressor_4_2 u2_2050(.a(s_217_19), .b(s_217_18), .c(s_217_17), .d(s_217_16), .cin(t_6010), .o(t_6023), .co(t_6024), .cout(t_6025));
compressor_4_2 u2_2051(.a(s_218_3), .b(s_218_2), .c(s_218_1), .d(s_218_0), .cin(t_6013), .o(t_6026), .co(t_6027), .cout(t_6028));
compressor_4_2 u2_2052(.a(s_218_7), .b(s_218_6), .c(s_218_5), .d(s_218_4), .cin(t_6016), .o(t_6029), .co(t_6030), .cout(t_6031));
compressor_4_2 u2_2053(.a(s_218_11), .b(s_218_10), .c(s_218_9), .d(s_218_8), .cin(t_6019), .o(t_6032), .co(t_6033), .cout(t_6034));
compressor_4_2 u2_2054(.a(s_218_15), .b(s_218_14), .c(s_218_13), .d(s_218_12), .cin(t_6022), .o(t_6035), .co(t_6036), .cout(t_6037));
compressor_4_2 u2_2055(.a(s_218_19), .b(s_218_18), .c(s_218_17), .d(s_218_16), .cin(t_6025), .o(t_6038), .co(t_6039), .cout(t_6040));
compressor_4_2 u2_2056(.a(s_219_3), .b(s_219_2), .c(s_219_1), .d(s_219_0), .cin(t_6028), .o(t_6041), .co(t_6042), .cout(t_6043));
compressor_4_2 u2_2057(.a(s_219_7), .b(s_219_6), .c(s_219_5), .d(s_219_4), .cin(t_6031), .o(t_6044), .co(t_6045), .cout(t_6046));
compressor_4_2 u2_2058(.a(s_219_11), .b(s_219_10), .c(s_219_9), .d(s_219_8), .cin(t_6034), .o(t_6047), .co(t_6048), .cout(t_6049));
compressor_4_2 u2_2059(.a(s_219_15), .b(s_219_14), .c(s_219_13), .d(s_219_12), .cin(t_6037), .o(t_6050), .co(t_6051), .cout(t_6052));
compressor_4_2 u2_2060(.a(s_219_19), .b(s_219_18), .c(s_219_17), .d(s_219_16), .cin(t_6040), .o(t_6053), .co(t_6054), .cout(t_6055));
compressor_4_2 u2_2061(.a(s_220_3), .b(s_220_2), .c(s_220_1), .d(s_220_0), .cin(t_6043), .o(t_6056), .co(t_6057), .cout(t_6058));
compressor_4_2 u2_2062(.a(s_220_7), .b(s_220_6), .c(s_220_5), .d(s_220_4), .cin(t_6046), .o(t_6059), .co(t_6060), .cout(t_6061));
compressor_4_2 u2_2063(.a(s_220_11), .b(s_220_10), .c(s_220_9), .d(s_220_8), .cin(t_6049), .o(t_6062), .co(t_6063), .cout(t_6064));
compressor_4_2 u2_2064(.a(s_220_15), .b(s_220_14), .c(s_220_13), .d(s_220_12), .cin(t_6052), .o(t_6065), .co(t_6066), .cout(t_6067));
compressor_3_2 u1_2065(.a(s_220_17), .b(s_220_16), .cin(t_6055), .o(t_6068), .cout(t_6069));
compressor_4_2 u2_2066(.a(s_221_3), .b(s_221_2), .c(s_221_1), .d(s_221_0), .cin(t_6058), .o(t_6070), .co(t_6071), .cout(t_6072));
compressor_4_2 u2_2067(.a(s_221_7), .b(s_221_6), .c(s_221_5), .d(s_221_4), .cin(t_6061), .o(t_6073), .co(t_6074), .cout(t_6075));
compressor_4_2 u2_2068(.a(s_221_11), .b(s_221_10), .c(s_221_9), .d(s_221_8), .cin(t_6064), .o(t_6076), .co(t_6077), .cout(t_6078));
compressor_4_2 u2_2069(.a(s_221_15), .b(s_221_14), .c(s_221_13), .d(s_221_12), .cin(t_6067), .o(t_6079), .co(t_6080), .cout(t_6081));
compressor_3_2 u1_2070(.a(s_221_18), .b(s_221_17), .cin(s_221_16), .o(t_6082), .cout(t_6083));
compressor_4_2 u2_2071(.a(s_222_3), .b(s_222_2), .c(s_222_1), .d(s_222_0), .cin(t_6072), .o(t_6084), .co(t_6085), .cout(t_6086));
compressor_4_2 u2_2072(.a(s_222_7), .b(s_222_6), .c(s_222_5), .d(s_222_4), .cin(t_6075), .o(t_6087), .co(t_6088), .cout(t_6089));
compressor_4_2 u2_2073(.a(s_222_11), .b(s_222_10), .c(s_222_9), .d(s_222_8), .cin(t_6078), .o(t_6090), .co(t_6091), .cout(t_6092));
compressor_4_2 u2_2074(.a(s_222_15), .b(s_222_14), .c(s_222_13), .d(s_222_12), .cin(t_6081), .o(t_6093), .co(t_6094), .cout(t_6095));
half_adder u0_2075(.a(s_222_17), .b(s_222_16), .o(t_6096), .cout(t_6097));
compressor_4_2 u2_2076(.a(s_223_3), .b(s_223_2), .c(s_223_1), .d(s_223_0), .cin(t_6086), .o(t_6098), .co(t_6099), .cout(t_6100));
compressor_4_2 u2_2077(.a(s_223_7), .b(s_223_6), .c(s_223_5), .d(s_223_4), .cin(t_6089), .o(t_6101), .co(t_6102), .cout(t_6103));
compressor_4_2 u2_2078(.a(s_223_11), .b(s_223_10), .c(s_223_9), .d(s_223_8), .cin(t_6092), .o(t_6104), .co(t_6105), .cout(t_6106));
compressor_4_2 u2_2079(.a(s_223_15), .b(s_223_14), .c(s_223_13), .d(s_223_12), .cin(t_6095), .o(t_6107), .co(t_6108), .cout(t_6109));
half_adder u0_2080(.a(s_223_17), .b(s_223_16), .o(t_6110), .cout(t_6111));
compressor_4_2 u2_2081(.a(s_224_3), .b(s_224_2), .c(s_224_1), .d(s_224_0), .cin(t_6100), .o(t_6112), .co(t_6113), .cout(t_6114));
compressor_4_2 u2_2082(.a(s_224_7), .b(s_224_6), .c(s_224_5), .d(s_224_4), .cin(t_6103), .o(t_6115), .co(t_6116), .cout(t_6117));
compressor_4_2 u2_2083(.a(s_224_11), .b(s_224_10), .c(s_224_9), .d(s_224_8), .cin(t_6106), .o(t_6118), .co(t_6119), .cout(t_6120));
compressor_4_2 u2_2084(.a(s_224_15), .b(s_224_14), .c(s_224_13), .d(s_224_12), .cin(t_6109), .o(t_6121), .co(t_6122), .cout(t_6123));
compressor_4_2 u2_2085(.a(s_225_3), .b(s_225_2), .c(s_225_1), .d(s_225_0), .cin(t_6114), .o(t_6124), .co(t_6125), .cout(t_6126));
compressor_4_2 u2_2086(.a(s_225_7), .b(s_225_6), .c(s_225_5), .d(s_225_4), .cin(t_6117), .o(t_6127), .co(t_6128), .cout(t_6129));
compressor_4_2 u2_2087(.a(s_225_11), .b(s_225_10), .c(s_225_9), .d(s_225_8), .cin(t_6120), .o(t_6130), .co(t_6131), .cout(t_6132));
compressor_4_2 u2_2088(.a(s_225_15), .b(s_225_14), .c(s_225_13), .d(s_225_12), .cin(t_6123), .o(t_6133), .co(t_6134), .cout(t_6135));
compressor_4_2 u2_2089(.a(s_226_3), .b(s_226_2), .c(s_226_1), .d(s_226_0), .cin(t_6126), .o(t_6136), .co(t_6137), .cout(t_6138));
compressor_4_2 u2_2090(.a(s_226_7), .b(s_226_6), .c(s_226_5), .d(s_226_4), .cin(t_6129), .o(t_6139), .co(t_6140), .cout(t_6141));
compressor_4_2 u2_2091(.a(s_226_11), .b(s_226_10), .c(s_226_9), .d(s_226_8), .cin(t_6132), .o(t_6142), .co(t_6143), .cout(t_6144));
compressor_4_2 u2_2092(.a(s_226_15), .b(s_226_14), .c(s_226_13), .d(s_226_12), .cin(t_6135), .o(t_6145), .co(t_6146), .cout(t_6147));
compressor_4_2 u2_2093(.a(s_227_3), .b(s_227_2), .c(s_227_1), .d(s_227_0), .cin(t_6138), .o(t_6148), .co(t_6149), .cout(t_6150));
compressor_4_2 u2_2094(.a(s_227_7), .b(s_227_6), .c(s_227_5), .d(s_227_4), .cin(t_6141), .o(t_6151), .co(t_6152), .cout(t_6153));
compressor_4_2 u2_2095(.a(s_227_11), .b(s_227_10), .c(s_227_9), .d(s_227_8), .cin(t_6144), .o(t_6154), .co(t_6155), .cout(t_6156));
compressor_4_2 u2_2096(.a(s_227_15), .b(s_227_14), .c(s_227_13), .d(s_227_12), .cin(t_6147), .o(t_6157), .co(t_6158), .cout(t_6159));
compressor_4_2 u2_2097(.a(s_228_3), .b(s_228_2), .c(s_228_1), .d(s_228_0), .cin(t_6150), .o(t_6160), .co(t_6161), .cout(t_6162));
compressor_4_2 u2_2098(.a(s_228_7), .b(s_228_6), .c(s_228_5), .d(s_228_4), .cin(t_6153), .o(t_6163), .co(t_6164), .cout(t_6165));
compressor_4_2 u2_2099(.a(s_228_11), .b(s_228_10), .c(s_228_9), .d(s_228_8), .cin(t_6156), .o(t_6166), .co(t_6167), .cout(t_6168));
compressor_3_2 u1_2100(.a(s_228_13), .b(s_228_12), .cin(t_6159), .o(t_6169), .cout(t_6170));
compressor_4_2 u2_2101(.a(s_229_3), .b(s_229_2), .c(s_229_1), .d(s_229_0), .cin(t_6162), .o(t_6171), .co(t_6172), .cout(t_6173));
compressor_4_2 u2_2102(.a(s_229_7), .b(s_229_6), .c(s_229_5), .d(s_229_4), .cin(t_6165), .o(t_6174), .co(t_6175), .cout(t_6176));
compressor_4_2 u2_2103(.a(s_229_11), .b(s_229_10), .c(s_229_9), .d(s_229_8), .cin(t_6168), .o(t_6177), .co(t_6178), .cout(t_6179));
compressor_3_2 u1_2104(.a(s_229_14), .b(s_229_13), .cin(s_229_12), .o(t_6180), .cout(t_6181));
compressor_4_2 u2_2105(.a(s_230_3), .b(s_230_2), .c(s_230_1), .d(s_230_0), .cin(t_6173), .o(t_6182), .co(t_6183), .cout(t_6184));
compressor_4_2 u2_2106(.a(s_230_7), .b(s_230_6), .c(s_230_5), .d(s_230_4), .cin(t_6176), .o(t_6185), .co(t_6186), .cout(t_6187));
compressor_4_2 u2_2107(.a(s_230_11), .b(s_230_10), .c(s_230_9), .d(s_230_8), .cin(t_6179), .o(t_6188), .co(t_6189), .cout(t_6190));
half_adder u0_2108(.a(s_230_13), .b(s_230_12), .o(t_6191), .cout(t_6192));
compressor_4_2 u2_2109(.a(s_231_3), .b(s_231_2), .c(s_231_1), .d(s_231_0), .cin(t_6184), .o(t_6193), .co(t_6194), .cout(t_6195));
compressor_4_2 u2_2110(.a(s_231_7), .b(s_231_6), .c(s_231_5), .d(s_231_4), .cin(t_6187), .o(t_6196), .co(t_6197), .cout(t_6198));
compressor_4_2 u2_2111(.a(s_231_11), .b(s_231_10), .c(s_231_9), .d(s_231_8), .cin(t_6190), .o(t_6199), .co(t_6200), .cout(t_6201));
half_adder u0_2112(.a(s_231_13), .b(s_231_12), .o(t_6202), .cout(t_6203));
compressor_4_2 u2_2113(.a(s_232_3), .b(s_232_2), .c(s_232_1), .d(s_232_0), .cin(t_6195), .o(t_6204), .co(t_6205), .cout(t_6206));
compressor_4_2 u2_2114(.a(s_232_7), .b(s_232_6), .c(s_232_5), .d(s_232_4), .cin(t_6198), .o(t_6207), .co(t_6208), .cout(t_6209));
compressor_4_2 u2_2115(.a(s_232_11), .b(s_232_10), .c(s_232_9), .d(s_232_8), .cin(t_6201), .o(t_6210), .co(t_6211), .cout(t_6212));
compressor_4_2 u2_2116(.a(s_233_3), .b(s_233_2), .c(s_233_1), .d(s_233_0), .cin(t_6206), .o(t_6213), .co(t_6214), .cout(t_6215));
compressor_4_2 u2_2117(.a(s_233_7), .b(s_233_6), .c(s_233_5), .d(s_233_4), .cin(t_6209), .o(t_6216), .co(t_6217), .cout(t_6218));
compressor_4_2 u2_2118(.a(s_233_11), .b(s_233_10), .c(s_233_9), .d(s_233_8), .cin(t_6212), .o(t_6219), .co(t_6220), .cout(t_6221));
compressor_4_2 u2_2119(.a(s_234_3), .b(s_234_2), .c(s_234_1), .d(s_234_0), .cin(t_6215), .o(t_6222), .co(t_6223), .cout(t_6224));
compressor_4_2 u2_2120(.a(s_234_7), .b(s_234_6), .c(s_234_5), .d(s_234_4), .cin(t_6218), .o(t_6225), .co(t_6226), .cout(t_6227));
compressor_4_2 u2_2121(.a(s_234_11), .b(s_234_10), .c(s_234_9), .d(s_234_8), .cin(t_6221), .o(t_6228), .co(t_6229), .cout(t_6230));
compressor_4_2 u2_2122(.a(s_235_3), .b(s_235_2), .c(s_235_1), .d(s_235_0), .cin(t_6224), .o(t_6231), .co(t_6232), .cout(t_6233));
compressor_4_2 u2_2123(.a(s_235_7), .b(s_235_6), .c(s_235_5), .d(s_235_4), .cin(t_6227), .o(t_6234), .co(t_6235), .cout(t_6236));
compressor_4_2 u2_2124(.a(s_235_11), .b(s_235_10), .c(s_235_9), .d(s_235_8), .cin(t_6230), .o(t_6237), .co(t_6238), .cout(t_6239));
compressor_4_2 u2_2125(.a(s_236_3), .b(s_236_2), .c(s_236_1), .d(s_236_0), .cin(t_6233), .o(t_6240), .co(t_6241), .cout(t_6242));
compressor_4_2 u2_2126(.a(s_236_7), .b(s_236_6), .c(s_236_5), .d(s_236_4), .cin(t_6236), .o(t_6243), .co(t_6244), .cout(t_6245));
compressor_3_2 u1_2127(.a(s_236_9), .b(s_236_8), .cin(t_6239), .o(t_6246), .cout(t_6247));
compressor_4_2 u2_2128(.a(s_237_3), .b(s_237_2), .c(s_237_1), .d(s_237_0), .cin(t_6242), .o(t_6248), .co(t_6249), .cout(t_6250));
compressor_4_2 u2_2129(.a(s_237_7), .b(s_237_6), .c(s_237_5), .d(s_237_4), .cin(t_6245), .o(t_6251), .co(t_6252), .cout(t_6253));
compressor_3_2 u1_2130(.a(s_237_10), .b(s_237_9), .cin(s_237_8), .o(t_6254), .cout(t_6255));
compressor_4_2 u2_2131(.a(s_238_3), .b(s_238_2), .c(s_238_1), .d(s_238_0), .cin(t_6250), .o(t_6256), .co(t_6257), .cout(t_6258));
compressor_4_2 u2_2132(.a(s_238_7), .b(s_238_6), .c(s_238_5), .d(s_238_4), .cin(t_6253), .o(t_6259), .co(t_6260), .cout(t_6261));
half_adder u0_2133(.a(s_238_9), .b(s_238_8), .o(t_6262), .cout(t_6263));
compressor_4_2 u2_2134(.a(s_239_3), .b(s_239_2), .c(s_239_1), .d(s_239_0), .cin(t_6258), .o(t_6264), .co(t_6265), .cout(t_6266));
compressor_4_2 u2_2135(.a(s_239_7), .b(s_239_6), .c(s_239_5), .d(s_239_4), .cin(t_6261), .o(t_6267), .co(t_6268), .cout(t_6269));
half_adder u0_2136(.a(s_239_9), .b(s_239_8), .o(t_6270), .cout(t_6271));
compressor_4_2 u2_2137(.a(s_240_3), .b(s_240_2), .c(s_240_1), .d(s_240_0), .cin(t_6266), .o(t_6272), .co(t_6273), .cout(t_6274));
compressor_4_2 u2_2138(.a(s_240_7), .b(s_240_6), .c(s_240_5), .d(s_240_4), .cin(t_6269), .o(t_6275), .co(t_6276), .cout(t_6277));
compressor_4_2 u2_2139(.a(s_241_3), .b(s_241_2), .c(s_241_1), .d(s_241_0), .cin(t_6274), .o(t_6278), .co(t_6279), .cout(t_6280));
compressor_4_2 u2_2140(.a(s_241_7), .b(s_241_6), .c(s_241_5), .d(s_241_4), .cin(t_6277), .o(t_6281), .co(t_6282), .cout(t_6283));
compressor_4_2 u2_2141(.a(s_242_3), .b(s_242_2), .c(s_242_1), .d(s_242_0), .cin(t_6280), .o(t_6284), .co(t_6285), .cout(t_6286));
compressor_4_2 u2_2142(.a(s_242_7), .b(s_242_6), .c(s_242_5), .d(s_242_4), .cin(t_6283), .o(t_6287), .co(t_6288), .cout(t_6289));
compressor_4_2 u2_2143(.a(s_243_3), .b(s_243_2), .c(s_243_1), .d(s_243_0), .cin(t_6286), .o(t_6290), .co(t_6291), .cout(t_6292));
compressor_4_2 u2_2144(.a(s_243_7), .b(s_243_6), .c(s_243_5), .d(s_243_4), .cin(t_6289), .o(t_6293), .co(t_6294), .cout(t_6295));
compressor_4_2 u2_2145(.a(s_244_3), .b(s_244_2), .c(s_244_1), .d(s_244_0), .cin(t_6292), .o(t_6296), .co(t_6297), .cout(t_6298));
compressor_3_2 u1_2146(.a(s_244_5), .b(s_244_4), .cin(t_6295), .o(t_6299), .cout(t_6300));
compressor_4_2 u2_2147(.a(s_245_3), .b(s_245_2), .c(s_245_1), .d(s_245_0), .cin(t_6298), .o(t_6301), .co(t_6302), .cout(t_6303));
compressor_3_2 u1_2148(.a(s_245_6), .b(s_245_5), .cin(s_245_4), .o(t_6304), .cout(t_6305));
compressor_4_2 u2_2149(.a(s_246_3), .b(s_246_2), .c(s_246_1), .d(s_246_0), .cin(t_6303), .o(t_6306), .co(t_6307), .cout(t_6308));
half_adder u0_2150(.a(s_246_5), .b(s_246_4), .o(t_6309), .cout(t_6310));
compressor_4_2 u2_2151(.a(s_247_3), .b(s_247_2), .c(s_247_1), .d(s_247_0), .cin(t_6308), .o(t_6311), .co(t_6312), .cout(t_6313));
half_adder u0_2152(.a(s_247_5), .b(s_247_4), .o(t_6314), .cout(t_6315));
compressor_4_2 u2_2153(.a(s_248_3), .b(s_248_2), .c(s_248_1), .d(s_248_0), .cin(t_6313), .o(t_6316), .co(t_6317), .cout(t_6318));
compressor_4_2 u2_2154(.a(s_249_3), .b(s_249_2), .c(s_249_1), .d(s_249_0), .cin(t_6318), .o(t_6319), .co(t_6320), .cout(t_6321));
compressor_4_2 u2_2155(.a(s_250_3), .b(s_250_2), .c(s_250_1), .d(s_250_0), .cin(t_6321), .o(t_6322), .co(t_6323), .cout(t_6324));
compressor_4_2 u2_2156(.a(s_251_3), .b(s_251_2), .c(s_251_1), .d(s_251_0), .cin(t_6324), .o(t_6325), .co(t_6326), .cout(t_6327));
compressor_3_2 u1_2157(.a(s_252_1), .b(s_252_0), .cin(t_6327), .o(t_6328), .cout(t_6329));
compressor_3_2 u1_2158(.a(s_253_2), .b(s_253_1), .cin(s_253_0), .o(t_6330), .cout(t_6331));
half_adder u0_2159(.a(s_254_1), .b(s_254_0), .o(t_6332), .cout(t_6333));
half_adder u0_2160(.a(s_255_1), .b(s_255_0), .o(t_6334), .cout());

/* u0_2161 Output nets */
wire t_6335,   t_6336;
/* u0_2162 Output nets */
wire t_6337,   t_6338;
/* u1_2163 Output nets */
wire t_6339,   t_6340;
/* u0_2164 Output nets */
wire t_6341,   t_6342;
/* u0_2165 Output nets */
wire t_6343,   t_6344;
/* u0_2166 Output nets */
wire t_6345,   t_6346;
/* u1_2167 Output nets */
wire t_6347,   t_6348;
/* u1_2168 Output nets */
wire t_6349,   t_6350;
/* u1_2169 Output nets */
wire t_6351,   t_6352;
/* u1_2170 Output nets */
wire t_6353,   t_6354;
/* u2_2171 Output nets */
wire t_6355,   t_6356,   t_6357;
/* u2_2172 Output nets */
wire t_6358,   t_6359,   t_6360;
/* u2_2173 Output nets */
wire t_6361,   t_6362,   t_6363;
/* u2_2174 Output nets */
wire t_6364,   t_6365,   t_6366;
/* u2_2175 Output nets */
wire t_6367,   t_6368,   t_6369;
/* u2_2176 Output nets */
wire t_6370,   t_6371,   t_6372;
/* u0_2177 Output nets */
wire t_6373,   t_6374;
/* u2_2178 Output nets */
wire t_6375,   t_6376,   t_6377;
/* u2_2179 Output nets */
wire t_6378,   t_6379,   t_6380;
/* u0_2180 Output nets */
wire t_6381,   t_6382;
/* u2_2181 Output nets */
wire t_6383,   t_6384,   t_6385;
/* u1_2182 Output nets */
wire t_6386,   t_6387;
/* u2_2183 Output nets */
wire t_6388,   t_6389,   t_6390;
/* u0_2184 Output nets */
wire t_6391,   t_6392;
/* u2_2185 Output nets */
wire t_6393,   t_6394,   t_6395;
/* u0_2186 Output nets */
wire t_6396,   t_6397;
/* u2_2187 Output nets */
wire t_6398,   t_6399,   t_6400;
/* u0_2188 Output nets */
wire t_6401,   t_6402;
/* u2_2189 Output nets */
wire t_6403,   t_6404,   t_6405;
/* u1_2190 Output nets */
wire t_6406,   t_6407;
/* u2_2191 Output nets */
wire t_6408,   t_6409,   t_6410;
/* u1_2192 Output nets */
wire t_6411,   t_6412;
/* u2_2193 Output nets */
wire t_6413,   t_6414,   t_6415;
/* u1_2194 Output nets */
wire t_6416,   t_6417;
/* u2_2195 Output nets */
wire t_6418,   t_6419,   t_6420;
/* u1_2196 Output nets */
wire t_6421,   t_6422;
/* u2_2197 Output nets */
wire t_6423,   t_6424,   t_6425;
/* u2_2198 Output nets */
wire t_6426,   t_6427,   t_6428;
/* u2_2199 Output nets */
wire t_6429,   t_6430,   t_6431;
/* u2_2200 Output nets */
wire t_6432,   t_6433,   t_6434;
/* u2_2201 Output nets */
wire t_6435,   t_6436,   t_6437;
/* u2_2202 Output nets */
wire t_6438,   t_6439,   t_6440;
/* u2_2203 Output nets */
wire t_6441,   t_6442,   t_6443;
/* u2_2204 Output nets */
wire t_6444,   t_6445,   t_6446;
/* u2_2205 Output nets */
wire t_6447,   t_6448,   t_6449;
/* u2_2206 Output nets */
wire t_6450,   t_6451,   t_6452;
/* u2_2207 Output nets */
wire t_6453,   t_6454,   t_6455;
/* u2_2208 Output nets */
wire t_6456,   t_6457,   t_6458;
/* u0_2209 Output nets */
wire t_6459,   t_6460;
/* u2_2210 Output nets */
wire t_6461,   t_6462,   t_6463;
/* u2_2211 Output nets */
wire t_6464,   t_6465,   t_6466;
/* u2_2212 Output nets */
wire t_6467,   t_6468,   t_6469;
/* u2_2213 Output nets */
wire t_6470,   t_6471,   t_6472;
/* u0_2214 Output nets */
wire t_6473,   t_6474;
/* u2_2215 Output nets */
wire t_6475,   t_6476,   t_6477;
/* u2_2216 Output nets */
wire t_6478,   t_6479,   t_6480;
/* u1_2217 Output nets */
wire t_6481,   t_6482;
/* u2_2218 Output nets */
wire t_6483,   t_6484,   t_6485;
/* u2_2219 Output nets */
wire t_6486,   t_6487,   t_6488;
/* u0_2220 Output nets */
wire t_6489,   t_6490;
/* u2_2221 Output nets */
wire t_6491,   t_6492,   t_6493;
/* u2_2222 Output nets */
wire t_6494,   t_6495,   t_6496;
/* u0_2223 Output nets */
wire t_6497,   t_6498;
/* u2_2224 Output nets */
wire t_6499,   t_6500,   t_6501;
/* u2_2225 Output nets */
wire t_6502,   t_6503,   t_6504;
/* u0_2226 Output nets */
wire t_6505,   t_6506;
/* u2_2227 Output nets */
wire t_6507,   t_6508,   t_6509;
/* u2_2228 Output nets */
wire t_6510,   t_6511,   t_6512;
/* u1_2229 Output nets */
wire t_6513,   t_6514;
/* u2_2230 Output nets */
wire t_6515,   t_6516,   t_6517;
/* u2_2231 Output nets */
wire t_6518,   t_6519,   t_6520;
/* u1_2232 Output nets */
wire t_6521,   t_6522;
/* u2_2233 Output nets */
wire t_6523,   t_6524,   t_6525;
/* u2_2234 Output nets */
wire t_6526,   t_6527,   t_6528;
/* u1_2235 Output nets */
wire t_6529,   t_6530;
/* u2_2236 Output nets */
wire t_6531,   t_6532,   t_6533;
/* u2_2237 Output nets */
wire t_6534,   t_6535,   t_6536;
/* u1_2238 Output nets */
wire t_6537,   t_6538;
/* u2_2239 Output nets */
wire t_6539,   t_6540,   t_6541;
/* u2_2240 Output nets */
wire t_6542,   t_6543,   t_6544;
/* u2_2241 Output nets */
wire t_6545,   t_6546,   t_6547;
/* u2_2242 Output nets */
wire t_6548,   t_6549,   t_6550;
/* u2_2243 Output nets */
wire t_6551,   t_6552,   t_6553;
/* u2_2244 Output nets */
wire t_6554,   t_6555,   t_6556;
/* u2_2245 Output nets */
wire t_6557,   t_6558,   t_6559;
/* u2_2246 Output nets */
wire t_6560,   t_6561,   t_6562;
/* u2_2247 Output nets */
wire t_6563,   t_6564,   t_6565;
/* u2_2248 Output nets */
wire t_6566,   t_6567,   t_6568;
/* u2_2249 Output nets */
wire t_6569,   t_6570,   t_6571;
/* u2_2250 Output nets */
wire t_6572,   t_6573,   t_6574;
/* u2_2251 Output nets */
wire t_6575,   t_6576,   t_6577;
/* u2_2252 Output nets */
wire t_6578,   t_6579,   t_6580;
/* u2_2253 Output nets */
wire t_6581,   t_6582,   t_6583;
/* u2_2254 Output nets */
wire t_6584,   t_6585,   t_6586;
/* u2_2255 Output nets */
wire t_6587,   t_6588,   t_6589;
/* u2_2256 Output nets */
wire t_6590,   t_6591,   t_6592;
/* u0_2257 Output nets */
wire t_6593,   t_6594;
/* u2_2258 Output nets */
wire t_6595,   t_6596,   t_6597;
/* u2_2259 Output nets */
wire t_6598,   t_6599,   t_6600;
/* u2_2260 Output nets */
wire t_6601,   t_6602,   t_6603;
/* u2_2261 Output nets */
wire t_6604,   t_6605,   t_6606;
/* u2_2262 Output nets */
wire t_6607,   t_6608,   t_6609;
/* u2_2263 Output nets */
wire t_6610,   t_6611,   t_6612;
/* u0_2264 Output nets */
wire t_6613,   t_6614;
/* u2_2265 Output nets */
wire t_6615,   t_6616,   t_6617;
/* u2_2266 Output nets */
wire t_6618,   t_6619,   t_6620;
/* u2_2267 Output nets */
wire t_6621,   t_6622,   t_6623;
/* u1_2268 Output nets */
wire t_6624,   t_6625;
/* u2_2269 Output nets */
wire t_6626,   t_6627,   t_6628;
/* u2_2270 Output nets */
wire t_6629,   t_6630,   t_6631;
/* u2_2271 Output nets */
wire t_6632,   t_6633,   t_6634;
/* u0_2272 Output nets */
wire t_6635,   t_6636;
/* u2_2273 Output nets */
wire t_6637,   t_6638,   t_6639;
/* u2_2274 Output nets */
wire t_6640,   t_6641,   t_6642;
/* u2_2275 Output nets */
wire t_6643,   t_6644,   t_6645;
/* u0_2276 Output nets */
wire t_6646,   t_6647;
/* u2_2277 Output nets */
wire t_6648,   t_6649,   t_6650;
/* u2_2278 Output nets */
wire t_6651,   t_6652,   t_6653;
/* u2_2279 Output nets */
wire t_6654,   t_6655,   t_6656;
/* u0_2280 Output nets */
wire t_6657,   t_6658;
/* u2_2281 Output nets */
wire t_6659,   t_6660,   t_6661;
/* u2_2282 Output nets */
wire t_6662,   t_6663,   t_6664;
/* u2_2283 Output nets */
wire t_6665,   t_6666,   t_6667;
/* u1_2284 Output nets */
wire t_6668,   t_6669;
/* u2_2285 Output nets */
wire t_6670,   t_6671,   t_6672;
/* u2_2286 Output nets */
wire t_6673,   t_6674,   t_6675;
/* u2_2287 Output nets */
wire t_6676,   t_6677,   t_6678;
/* u1_2288 Output nets */
wire t_6679,   t_6680;
/* u2_2289 Output nets */
wire t_6681,   t_6682,   t_6683;
/* u2_2290 Output nets */
wire t_6684,   t_6685,   t_6686;
/* u2_2291 Output nets */
wire t_6687,   t_6688,   t_6689;
/* u1_2292 Output nets */
wire t_6690,   t_6691;
/* u2_2293 Output nets */
wire t_6692,   t_6693,   t_6694;
/* u2_2294 Output nets */
wire t_6695,   t_6696,   t_6697;
/* u2_2295 Output nets */
wire t_6698,   t_6699,   t_6700;
/* u1_2296 Output nets */
wire t_6701,   t_6702;
/* u2_2297 Output nets */
wire t_6703,   t_6704,   t_6705;
/* u2_2298 Output nets */
wire t_6706,   t_6707,   t_6708;
/* u2_2299 Output nets */
wire t_6709,   t_6710,   t_6711;
/* u2_2300 Output nets */
wire t_6712,   t_6713,   t_6714;
/* u2_2301 Output nets */
wire t_6715,   t_6716,   t_6717;
/* u2_2302 Output nets */
wire t_6718,   t_6719,   t_6720;
/* u2_2303 Output nets */
wire t_6721,   t_6722,   t_6723;
/* u2_2304 Output nets */
wire t_6724,   t_6725,   t_6726;
/* u2_2305 Output nets */
wire t_6727,   t_6728,   t_6729;
/* u2_2306 Output nets */
wire t_6730,   t_6731,   t_6732;
/* u2_2307 Output nets */
wire t_6733,   t_6734,   t_6735;
/* u2_2308 Output nets */
wire t_6736,   t_6737,   t_6738;
/* u2_2309 Output nets */
wire t_6739,   t_6740,   t_6741;
/* u2_2310 Output nets */
wire t_6742,   t_6743,   t_6744;
/* u2_2311 Output nets */
wire t_6745,   t_6746,   t_6747;
/* u2_2312 Output nets */
wire t_6748,   t_6749,   t_6750;
/* u2_2313 Output nets */
wire t_6751,   t_6752,   t_6753;
/* u2_2314 Output nets */
wire t_6754,   t_6755,   t_6756;
/* u2_2315 Output nets */
wire t_6757,   t_6758,   t_6759;
/* u2_2316 Output nets */
wire t_6760,   t_6761,   t_6762;
/* u2_2317 Output nets */
wire t_6763,   t_6764,   t_6765;
/* u2_2318 Output nets */
wire t_6766,   t_6767,   t_6768;
/* u2_2319 Output nets */
wire t_6769,   t_6770,   t_6771;
/* u2_2320 Output nets */
wire t_6772,   t_6773,   t_6774;
/* u0_2321 Output nets */
wire t_6775,   t_6776;
/* u2_2322 Output nets */
wire t_6777,   t_6778,   t_6779;
/* u2_2323 Output nets */
wire t_6780,   t_6781,   t_6782;
/* u2_2324 Output nets */
wire t_6783,   t_6784,   t_6785;
/* u2_2325 Output nets */
wire t_6786,   t_6787,   t_6788;
/* u2_2326 Output nets */
wire t_6789,   t_6790,   t_6791;
/* u2_2327 Output nets */
wire t_6792,   t_6793,   t_6794;
/* u2_2328 Output nets */
wire t_6795,   t_6796,   t_6797;
/* u2_2329 Output nets */
wire t_6798,   t_6799,   t_6800;
/* u0_2330 Output nets */
wire t_6801,   t_6802;
/* u2_2331 Output nets */
wire t_6803,   t_6804,   t_6805;
/* u2_2332 Output nets */
wire t_6806,   t_6807,   t_6808;
/* u2_2333 Output nets */
wire t_6809,   t_6810,   t_6811;
/* u2_2334 Output nets */
wire t_6812,   t_6813,   t_6814;
/* u1_2335 Output nets */
wire t_6815,   t_6816;
/* u2_2336 Output nets */
wire t_6817,   t_6818,   t_6819;
/* u2_2337 Output nets */
wire t_6820,   t_6821,   t_6822;
/* u2_2338 Output nets */
wire t_6823,   t_6824,   t_6825;
/* u2_2339 Output nets */
wire t_6826,   t_6827,   t_6828;
/* u0_2340 Output nets */
wire t_6829,   t_6830;
/* u2_2341 Output nets */
wire t_6831,   t_6832,   t_6833;
/* u2_2342 Output nets */
wire t_6834,   t_6835,   t_6836;
/* u2_2343 Output nets */
wire t_6837,   t_6838,   t_6839;
/* u2_2344 Output nets */
wire t_6840,   t_6841,   t_6842;
/* u0_2345 Output nets */
wire t_6843,   t_6844;
/* u2_2346 Output nets */
wire t_6845,   t_6846,   t_6847;
/* u2_2347 Output nets */
wire t_6848,   t_6849,   t_6850;
/* u2_2348 Output nets */
wire t_6851,   t_6852,   t_6853;
/* u2_2349 Output nets */
wire t_6854,   t_6855,   t_6856;
/* u0_2350 Output nets */
wire t_6857,   t_6858;
/* u2_2351 Output nets */
wire t_6859,   t_6860,   t_6861;
/* u2_2352 Output nets */
wire t_6862,   t_6863,   t_6864;
/* u2_2353 Output nets */
wire t_6865,   t_6866,   t_6867;
/* u2_2354 Output nets */
wire t_6868,   t_6869,   t_6870;
/* u1_2355 Output nets */
wire t_6871,   t_6872;
/* u2_2356 Output nets */
wire t_6873,   t_6874,   t_6875;
/* u2_2357 Output nets */
wire t_6876,   t_6877,   t_6878;
/* u2_2358 Output nets */
wire t_6879,   t_6880,   t_6881;
/* u2_2359 Output nets */
wire t_6882,   t_6883,   t_6884;
/* u1_2360 Output nets */
wire t_6885,   t_6886;
/* u2_2361 Output nets */
wire t_6887,   t_6888,   t_6889;
/* u2_2362 Output nets */
wire t_6890,   t_6891,   t_6892;
/* u2_2363 Output nets */
wire t_6893,   t_6894,   t_6895;
/* u2_2364 Output nets */
wire t_6896,   t_6897,   t_6898;
/* u1_2365 Output nets */
wire t_6899,   t_6900;
/* u2_2366 Output nets */
wire t_6901,   t_6902,   t_6903;
/* u2_2367 Output nets */
wire t_6904,   t_6905,   t_6906;
/* u2_2368 Output nets */
wire t_6907,   t_6908,   t_6909;
/* u2_2369 Output nets */
wire t_6910,   t_6911,   t_6912;
/* u1_2370 Output nets */
wire t_6913,   t_6914;
/* u2_2371 Output nets */
wire t_6915,   t_6916,   t_6917;
/* u2_2372 Output nets */
wire t_6918,   t_6919,   t_6920;
/* u2_2373 Output nets */
wire t_6921,   t_6922,   t_6923;
/* u2_2374 Output nets */
wire t_6924,   t_6925,   t_6926;
/* u2_2375 Output nets */
wire t_6927,   t_6928,   t_6929;
/* u2_2376 Output nets */
wire t_6930,   t_6931,   t_6932;
/* u2_2377 Output nets */
wire t_6933,   t_6934,   t_6935;
/* u2_2378 Output nets */
wire t_6936,   t_6937,   t_6938;
/* u2_2379 Output nets */
wire t_6939,   t_6940,   t_6941;
/* u2_2380 Output nets */
wire t_6942,   t_6943,   t_6944;
/* u2_2381 Output nets */
wire t_6945,   t_6946,   t_6947;
/* u2_2382 Output nets */
wire t_6948,   t_6949,   t_6950;
/* u2_2383 Output nets */
wire t_6951,   t_6952,   t_6953;
/* u2_2384 Output nets */
wire t_6954,   t_6955,   t_6956;
/* u2_2385 Output nets */
wire t_6957,   t_6958,   t_6959;
/* u2_2386 Output nets */
wire t_6960,   t_6961,   t_6962;
/* u2_2387 Output nets */
wire t_6963,   t_6964,   t_6965;
/* u2_2388 Output nets */
wire t_6966,   t_6967,   t_6968;
/* u2_2389 Output nets */
wire t_6969,   t_6970,   t_6971;
/* u2_2390 Output nets */
wire t_6972,   t_6973,   t_6974;
/* u2_2391 Output nets */
wire t_6975,   t_6976,   t_6977;
/* u2_2392 Output nets */
wire t_6978,   t_6979,   t_6980;
/* u2_2393 Output nets */
wire t_6981,   t_6982,   t_6983;
/* u2_2394 Output nets */
wire t_6984,   t_6985,   t_6986;
/* u2_2395 Output nets */
wire t_6987,   t_6988,   t_6989;
/* u2_2396 Output nets */
wire t_6990,   t_6991,   t_6992;
/* u2_2397 Output nets */
wire t_6993,   t_6994,   t_6995;
/* u2_2398 Output nets */
wire t_6996,   t_6997,   t_6998;
/* u2_2399 Output nets */
wire t_6999,   t_7000,   t_7001;
/* u2_2400 Output nets */
wire t_7002,   t_7003,   t_7004;
/* u0_2401 Output nets */
wire t_7005,   t_7006;
/* u2_2402 Output nets */
wire t_7007,   t_7008,   t_7009;
/* u2_2403 Output nets */
wire t_7010,   t_7011,   t_7012;
/* u2_2404 Output nets */
wire t_7013,   t_7014,   t_7015;
/* u2_2405 Output nets */
wire t_7016,   t_7017,   t_7018;
/* u2_2406 Output nets */
wire t_7019,   t_7020,   t_7021;
/* u2_2407 Output nets */
wire t_7022,   t_7023,   t_7024;
/* u2_2408 Output nets */
wire t_7025,   t_7026,   t_7027;
/* u2_2409 Output nets */
wire t_7028,   t_7029,   t_7030;
/* u2_2410 Output nets */
wire t_7031,   t_7032,   t_7033;
/* u2_2411 Output nets */
wire t_7034,   t_7035,   t_7036;
/* u0_2412 Output nets */
wire t_7037,   t_7038;
/* u2_2413 Output nets */
wire t_7039,   t_7040,   t_7041;
/* u2_2414 Output nets */
wire t_7042,   t_7043,   t_7044;
/* u2_2415 Output nets */
wire t_7045,   t_7046,   t_7047;
/* u2_2416 Output nets */
wire t_7048,   t_7049,   t_7050;
/* u2_2417 Output nets */
wire t_7051,   t_7052,   t_7053;
/* u1_2418 Output nets */
wire t_7054,   t_7055;
/* u2_2419 Output nets */
wire t_7056,   t_7057,   t_7058;
/* u2_2420 Output nets */
wire t_7059,   t_7060,   t_7061;
/* u2_2421 Output nets */
wire t_7062,   t_7063,   t_7064;
/* u2_2422 Output nets */
wire t_7065,   t_7066,   t_7067;
/* u2_2423 Output nets */
wire t_7068,   t_7069,   t_7070;
/* u0_2424 Output nets */
wire t_7071,   t_7072;
/* u2_2425 Output nets */
wire t_7073,   t_7074,   t_7075;
/* u2_2426 Output nets */
wire t_7076,   t_7077,   t_7078;
/* u2_2427 Output nets */
wire t_7079,   t_7080,   t_7081;
/* u2_2428 Output nets */
wire t_7082,   t_7083,   t_7084;
/* u2_2429 Output nets */
wire t_7085,   t_7086,   t_7087;
/* u0_2430 Output nets */
wire t_7088,   t_7089;
/* u2_2431 Output nets */
wire t_7090,   t_7091,   t_7092;
/* u2_2432 Output nets */
wire t_7093,   t_7094,   t_7095;
/* u2_2433 Output nets */
wire t_7096,   t_7097,   t_7098;
/* u2_2434 Output nets */
wire t_7099,   t_7100,   t_7101;
/* u2_2435 Output nets */
wire t_7102,   t_7103,   t_7104;
/* u0_2436 Output nets */
wire t_7105,   t_7106;
/* u2_2437 Output nets */
wire t_7107,   t_7108,   t_7109;
/* u2_2438 Output nets */
wire t_7110,   t_7111,   t_7112;
/* u2_2439 Output nets */
wire t_7113,   t_7114,   t_7115;
/* u2_2440 Output nets */
wire t_7116,   t_7117,   t_7118;
/* u2_2441 Output nets */
wire t_7119,   t_7120,   t_7121;
/* u1_2442 Output nets */
wire t_7122,   t_7123;
/* u2_2443 Output nets */
wire t_7124,   t_7125,   t_7126;
/* u2_2444 Output nets */
wire t_7127,   t_7128,   t_7129;
/* u2_2445 Output nets */
wire t_7130,   t_7131,   t_7132;
/* u2_2446 Output nets */
wire t_7133,   t_7134,   t_7135;
/* u2_2447 Output nets */
wire t_7136,   t_7137,   t_7138;
/* u1_2448 Output nets */
wire t_7139,   t_7140;
/* u2_2449 Output nets */
wire t_7141,   t_7142,   t_7143;
/* u2_2450 Output nets */
wire t_7144,   t_7145,   t_7146;
/* u2_2451 Output nets */
wire t_7147,   t_7148,   t_7149;
/* u2_2452 Output nets */
wire t_7150,   t_7151,   t_7152;
/* u2_2453 Output nets */
wire t_7153,   t_7154,   t_7155;
/* u1_2454 Output nets */
wire t_7156,   t_7157;
/* u2_2455 Output nets */
wire t_7158,   t_7159,   t_7160;
/* u2_2456 Output nets */
wire t_7161,   t_7162,   t_7163;
/* u2_2457 Output nets */
wire t_7164,   t_7165,   t_7166;
/* u2_2458 Output nets */
wire t_7167,   t_7168,   t_7169;
/* u2_2459 Output nets */
wire t_7170,   t_7171,   t_7172;
/* u1_2460 Output nets */
wire t_7173,   t_7174;
/* u2_2461 Output nets */
wire t_7175,   t_7176,   t_7177;
/* u2_2462 Output nets */
wire t_7178,   t_7179,   t_7180;
/* u2_2463 Output nets */
wire t_7181,   t_7182,   t_7183;
/* u2_2464 Output nets */
wire t_7184,   t_7185,   t_7186;
/* u2_2465 Output nets */
wire t_7187,   t_7188,   t_7189;
/* u2_2466 Output nets */
wire t_7190,   t_7191,   t_7192;
/* u2_2467 Output nets */
wire t_7193,   t_7194,   t_7195;
/* u2_2468 Output nets */
wire t_7196,   t_7197,   t_7198;
/* u2_2469 Output nets */
wire t_7199,   t_7200,   t_7201;
/* u2_2470 Output nets */
wire t_7202,   t_7203,   t_7204;
/* u2_2471 Output nets */
wire t_7205,   t_7206,   t_7207;
/* u2_2472 Output nets */
wire t_7208,   t_7209,   t_7210;
/* u2_2473 Output nets */
wire t_7211,   t_7212,   t_7213;
/* u2_2474 Output nets */
wire t_7214,   t_7215,   t_7216;
/* u2_2475 Output nets */
wire t_7217,   t_7218,   t_7219;
/* u2_2476 Output nets */
wire t_7220,   t_7221,   t_7222;
/* u2_2477 Output nets */
wire t_7223,   t_7224,   t_7225;
/* u2_2478 Output nets */
wire t_7226,   t_7227,   t_7228;
/* u2_2479 Output nets */
wire t_7229,   t_7230,   t_7231;
/* u2_2480 Output nets */
wire t_7232,   t_7233,   t_7234;
/* u2_2481 Output nets */
wire t_7235,   t_7236,   t_7237;
/* u2_2482 Output nets */
wire t_7238,   t_7239,   t_7240;
/* u2_2483 Output nets */
wire t_7241,   t_7242,   t_7243;
/* u2_2484 Output nets */
wire t_7244,   t_7245,   t_7246;
/* u2_2485 Output nets */
wire t_7247,   t_7248,   t_7249;
/* u2_2486 Output nets */
wire t_7250,   t_7251,   t_7252;
/* u2_2487 Output nets */
wire t_7253,   t_7254,   t_7255;
/* u2_2488 Output nets */
wire t_7256,   t_7257,   t_7258;
/* u2_2489 Output nets */
wire t_7259,   t_7260,   t_7261;
/* u2_2490 Output nets */
wire t_7262,   t_7263,   t_7264;
/* u2_2491 Output nets */
wire t_7265,   t_7266,   t_7267;
/* u2_2492 Output nets */
wire t_7268,   t_7269,   t_7270;
/* u2_2493 Output nets */
wire t_7271,   t_7272,   t_7273;
/* u2_2494 Output nets */
wire t_7274,   t_7275,   t_7276;
/* u2_2495 Output nets */
wire t_7277,   t_7278,   t_7279;
/* u2_2496 Output nets */
wire t_7280,   t_7281,   t_7282;
/* u0_2497 Output nets */
wire t_7283,   t_7284;
/* u2_2498 Output nets */
wire t_7285,   t_7286,   t_7287;
/* u2_2499 Output nets */
wire t_7288,   t_7289,   t_7290;
/* u2_2500 Output nets */
wire t_7291,   t_7292,   t_7293;
/* u2_2501 Output nets */
wire t_7294,   t_7295,   t_7296;
/* u2_2502 Output nets */
wire t_7297,   t_7298,   t_7299;
/* u2_2503 Output nets */
wire t_7300,   t_7301,   t_7302;
/* u2_2504 Output nets */
wire t_7303,   t_7304,   t_7305;
/* u2_2505 Output nets */
wire t_7306,   t_7307,   t_7308;
/* u2_2506 Output nets */
wire t_7309,   t_7310,   t_7311;
/* u2_2507 Output nets */
wire t_7312,   t_7313,   t_7314;
/* u2_2508 Output nets */
wire t_7315,   t_7316,   t_7317;
/* u2_2509 Output nets */
wire t_7318,   t_7319,   t_7320;
/* u0_2510 Output nets */
wire t_7321,   t_7322;
/* u2_2511 Output nets */
wire t_7323,   t_7324,   t_7325;
/* u2_2512 Output nets */
wire t_7326,   t_7327,   t_7328;
/* u2_2513 Output nets */
wire t_7329,   t_7330,   t_7331;
/* u2_2514 Output nets */
wire t_7332,   t_7333,   t_7334;
/* u2_2515 Output nets */
wire t_7335,   t_7336,   t_7337;
/* u2_2516 Output nets */
wire t_7338,   t_7339,   t_7340;
/* u1_2517 Output nets */
wire t_7341,   t_7342;
/* u2_2518 Output nets */
wire t_7343,   t_7344,   t_7345;
/* u2_2519 Output nets */
wire t_7346,   t_7347,   t_7348;
/* u2_2520 Output nets */
wire t_7349,   t_7350,   t_7351;
/* u2_2521 Output nets */
wire t_7352,   t_7353,   t_7354;
/* u2_2522 Output nets */
wire t_7355,   t_7356,   t_7357;
/* u2_2523 Output nets */
wire t_7358,   t_7359,   t_7360;
/* u0_2524 Output nets */
wire t_7361,   t_7362;
/* u2_2525 Output nets */
wire t_7363,   t_7364,   t_7365;
/* u2_2526 Output nets */
wire t_7366,   t_7367,   t_7368;
/* u2_2527 Output nets */
wire t_7369,   t_7370,   t_7371;
/* u2_2528 Output nets */
wire t_7372,   t_7373,   t_7374;
/* u2_2529 Output nets */
wire t_7375,   t_7376,   t_7377;
/* u2_2530 Output nets */
wire t_7378,   t_7379,   t_7380;
/* u0_2531 Output nets */
wire t_7381,   t_7382;
/* u2_2532 Output nets */
wire t_7383,   t_7384,   t_7385;
/* u2_2533 Output nets */
wire t_7386,   t_7387,   t_7388;
/* u2_2534 Output nets */
wire t_7389,   t_7390,   t_7391;
/* u2_2535 Output nets */
wire t_7392,   t_7393,   t_7394;
/* u2_2536 Output nets */
wire t_7395,   t_7396,   t_7397;
/* u2_2537 Output nets */
wire t_7398,   t_7399,   t_7400;
/* u0_2538 Output nets */
wire t_7401,   t_7402;
/* u2_2539 Output nets */
wire t_7403,   t_7404,   t_7405;
/* u2_2540 Output nets */
wire t_7406,   t_7407,   t_7408;
/* u2_2541 Output nets */
wire t_7409,   t_7410,   t_7411;
/* u2_2542 Output nets */
wire t_7412,   t_7413,   t_7414;
/* u2_2543 Output nets */
wire t_7415,   t_7416,   t_7417;
/* u2_2544 Output nets */
wire t_7418,   t_7419,   t_7420;
/* u1_2545 Output nets */
wire t_7421,   t_7422;
/* u2_2546 Output nets */
wire t_7423,   t_7424,   t_7425;
/* u2_2547 Output nets */
wire t_7426,   t_7427,   t_7428;
/* u2_2548 Output nets */
wire t_7429,   t_7430,   t_7431;
/* u2_2549 Output nets */
wire t_7432,   t_7433,   t_7434;
/* u2_2550 Output nets */
wire t_7435,   t_7436,   t_7437;
/* u2_2551 Output nets */
wire t_7438,   t_7439,   t_7440;
/* u1_2552 Output nets */
wire t_7441,   t_7442;
/* u2_2553 Output nets */
wire t_7443,   t_7444,   t_7445;
/* u2_2554 Output nets */
wire t_7446,   t_7447,   t_7448;
/* u2_2555 Output nets */
wire t_7449,   t_7450,   t_7451;
/* u2_2556 Output nets */
wire t_7452,   t_7453,   t_7454;
/* u2_2557 Output nets */
wire t_7455,   t_7456,   t_7457;
/* u2_2558 Output nets */
wire t_7458,   t_7459,   t_7460;
/* u1_2559 Output nets */
wire t_7461,   t_7462;
/* u2_2560 Output nets */
wire t_7463,   t_7464,   t_7465;
/* u2_2561 Output nets */
wire t_7466,   t_7467,   t_7468;
/* u2_2562 Output nets */
wire t_7469,   t_7470,   t_7471;
/* u2_2563 Output nets */
wire t_7472,   t_7473,   t_7474;
/* u2_2564 Output nets */
wire t_7475,   t_7476,   t_7477;
/* u2_2565 Output nets */
wire t_7478,   t_7479,   t_7480;
/* u1_2566 Output nets */
wire t_7481,   t_7482;
/* u2_2567 Output nets */
wire t_7483,   t_7484,   t_7485;
/* u2_2568 Output nets */
wire t_7486,   t_7487,   t_7488;
/* u2_2569 Output nets */
wire t_7489,   t_7490,   t_7491;
/* u2_2570 Output nets */
wire t_7492,   t_7493,   t_7494;
/* u2_2571 Output nets */
wire t_7495,   t_7496,   t_7497;
/* u2_2572 Output nets */
wire t_7498,   t_7499,   t_7500;
/* u2_2573 Output nets */
wire t_7501,   t_7502,   t_7503;
/* u2_2574 Output nets */
wire t_7504,   t_7505,   t_7506;
/* u2_2575 Output nets */
wire t_7507,   t_7508,   t_7509;
/* u2_2576 Output nets */
wire t_7510,   t_7511,   t_7512;
/* u2_2577 Output nets */
wire t_7513,   t_7514,   t_7515;
/* u2_2578 Output nets */
wire t_7516,   t_7517,   t_7518;
/* u2_2579 Output nets */
wire t_7519,   t_7520,   t_7521;
/* u2_2580 Output nets */
wire t_7522,   t_7523,   t_7524;
/* u2_2581 Output nets */
wire t_7525,   t_7526,   t_7527;
/* u2_2582 Output nets */
wire t_7528,   t_7529,   t_7530;
/* u2_2583 Output nets */
wire t_7531,   t_7532,   t_7533;
/* u2_2584 Output nets */
wire t_7534,   t_7535,   t_7536;
/* u2_2585 Output nets */
wire t_7537,   t_7538,   t_7539;
/* u2_2586 Output nets */
wire t_7540,   t_7541,   t_7542;
/* u2_2587 Output nets */
wire t_7543,   t_7544,   t_7545;
/* u2_2588 Output nets */
wire t_7546,   t_7547,   t_7548;
/* u2_2589 Output nets */
wire t_7549,   t_7550,   t_7551;
/* u2_2590 Output nets */
wire t_7552,   t_7553,   t_7554;
/* u2_2591 Output nets */
wire t_7555,   t_7556,   t_7557;
/* u2_2592 Output nets */
wire t_7558,   t_7559,   t_7560;
/* u2_2593 Output nets */
wire t_7561,   t_7562,   t_7563;
/* u2_2594 Output nets */
wire t_7564,   t_7565,   t_7566;
/* u2_2595 Output nets */
wire t_7567,   t_7568,   t_7569;
/* u2_2596 Output nets */
wire t_7570,   t_7571,   t_7572;
/* u2_2597 Output nets */
wire t_7573,   t_7574,   t_7575;
/* u2_2598 Output nets */
wire t_7576,   t_7577,   t_7578;
/* u2_2599 Output nets */
wire t_7579,   t_7580,   t_7581;
/* u2_2600 Output nets */
wire t_7582,   t_7583,   t_7584;
/* u2_2601 Output nets */
wire t_7585,   t_7586,   t_7587;
/* u2_2602 Output nets */
wire t_7588,   t_7589,   t_7590;
/* u2_2603 Output nets */
wire t_7591,   t_7592,   t_7593;
/* u2_2604 Output nets */
wire t_7594,   t_7595,   t_7596;
/* u2_2605 Output nets */
wire t_7597,   t_7598,   t_7599;
/* u2_2606 Output nets */
wire t_7600,   t_7601,   t_7602;
/* u2_2607 Output nets */
wire t_7603,   t_7604,   t_7605;
/* u2_2608 Output nets */
wire t_7606,   t_7607,   t_7608;
/* u0_2609 Output nets */
wire t_7609,   t_7610;
/* u2_2610 Output nets */
wire t_7611,   t_7612,   t_7613;
/* u2_2611 Output nets */
wire t_7614,   t_7615,   t_7616;
/* u2_2612 Output nets */
wire t_7617,   t_7618,   t_7619;
/* u2_2613 Output nets */
wire t_7620,   t_7621,   t_7622;
/* u2_2614 Output nets */
wire t_7623,   t_7624,   t_7625;
/* u2_2615 Output nets */
wire t_7626,   t_7627,   t_7628;
/* u2_2616 Output nets */
wire t_7629,   t_7630,   t_7631;
/* u2_2617 Output nets */
wire t_7632,   t_7633,   t_7634;
/* u2_2618 Output nets */
wire t_7635,   t_7636,   t_7637;
/* u2_2619 Output nets */
wire t_7638,   t_7639,   t_7640;
/* u2_2620 Output nets */
wire t_7641,   t_7642,   t_7643;
/* u2_2621 Output nets */
wire t_7644,   t_7645,   t_7646;
/* u2_2622 Output nets */
wire t_7647,   t_7648,   t_7649;
/* u2_2623 Output nets */
wire t_7650,   t_7651,   t_7652;
/* u0_2624 Output nets */
wire t_7653,   t_7654;
/* u2_2625 Output nets */
wire t_7655,   t_7656,   t_7657;
/* u2_2626 Output nets */
wire t_7658,   t_7659,   t_7660;
/* u2_2627 Output nets */
wire t_7661,   t_7662,   t_7663;
/* u2_2628 Output nets */
wire t_7664,   t_7665,   t_7666;
/* u2_2629 Output nets */
wire t_7667,   t_7668,   t_7669;
/* u2_2630 Output nets */
wire t_7670,   t_7671,   t_7672;
/* u2_2631 Output nets */
wire t_7673,   t_7674,   t_7675;
/* u1_2632 Output nets */
wire t_7676,   t_7677;
/* u2_2633 Output nets */
wire t_7678,   t_7679,   t_7680;
/* u2_2634 Output nets */
wire t_7681,   t_7682,   t_7683;
/* u2_2635 Output nets */
wire t_7684,   t_7685,   t_7686;
/* u2_2636 Output nets */
wire t_7687,   t_7688,   t_7689;
/* u2_2637 Output nets */
wire t_7690,   t_7691,   t_7692;
/* u2_2638 Output nets */
wire t_7693,   t_7694,   t_7695;
/* u2_2639 Output nets */
wire t_7696,   t_7697,   t_7698;
/* u0_2640 Output nets */
wire t_7699,   t_7700;
/* u2_2641 Output nets */
wire t_7701,   t_7702,   t_7703;
/* u2_2642 Output nets */
wire t_7704,   t_7705,   t_7706;
/* u2_2643 Output nets */
wire t_7707,   t_7708,   t_7709;
/* u2_2644 Output nets */
wire t_7710,   t_7711,   t_7712;
/* u2_2645 Output nets */
wire t_7713,   t_7714,   t_7715;
/* u2_2646 Output nets */
wire t_7716,   t_7717,   t_7718;
/* u2_2647 Output nets */
wire t_7719,   t_7720,   t_7721;
/* u0_2648 Output nets */
wire t_7722,   t_7723;
/* u2_2649 Output nets */
wire t_7724,   t_7725,   t_7726;
/* u2_2650 Output nets */
wire t_7727,   t_7728,   t_7729;
/* u2_2651 Output nets */
wire t_7730,   t_7731,   t_7732;
/* u2_2652 Output nets */
wire t_7733,   t_7734,   t_7735;
/* u2_2653 Output nets */
wire t_7736,   t_7737,   t_7738;
/* u2_2654 Output nets */
wire t_7739,   t_7740,   t_7741;
/* u2_2655 Output nets */
wire t_7742,   t_7743,   t_7744;
/* u0_2656 Output nets */
wire t_7745,   t_7746;
/* u2_2657 Output nets */
wire t_7747,   t_7748,   t_7749;
/* u2_2658 Output nets */
wire t_7750,   t_7751,   t_7752;
/* u2_2659 Output nets */
wire t_7753,   t_7754,   t_7755;
/* u2_2660 Output nets */
wire t_7756,   t_7757,   t_7758;
/* u2_2661 Output nets */
wire t_7759,   t_7760,   t_7761;
/* u2_2662 Output nets */
wire t_7762,   t_7763,   t_7764;
/* u2_2663 Output nets */
wire t_7765,   t_7766,   t_7767;
/* u1_2664 Output nets */
wire t_7768,   t_7769;
/* u2_2665 Output nets */
wire t_7770,   t_7771,   t_7772;
/* u2_2666 Output nets */
wire t_7773,   t_7774,   t_7775;
/* u2_2667 Output nets */
wire t_7776,   t_7777,   t_7778;
/* u2_2668 Output nets */
wire t_7779,   t_7780,   t_7781;
/* u2_2669 Output nets */
wire t_7782,   t_7783,   t_7784;
/* u2_2670 Output nets */
wire t_7785,   t_7786,   t_7787;
/* u2_2671 Output nets */
wire t_7788,   t_7789,   t_7790;
/* u1_2672 Output nets */
wire t_7791,   t_7792;
/* u2_2673 Output nets */
wire t_7793,   t_7794,   t_7795;
/* u2_2674 Output nets */
wire t_7796,   t_7797,   t_7798;
/* u2_2675 Output nets */
wire t_7799,   t_7800,   t_7801;
/* u2_2676 Output nets */
wire t_7802,   t_7803,   t_7804;
/* u2_2677 Output nets */
wire t_7805,   t_7806,   t_7807;
/* u2_2678 Output nets */
wire t_7808,   t_7809,   t_7810;
/* u2_2679 Output nets */
wire t_7811,   t_7812,   t_7813;
/* u1_2680 Output nets */
wire t_7814,   t_7815;
/* u2_2681 Output nets */
wire t_7816,   t_7817,   t_7818;
/* u2_2682 Output nets */
wire t_7819,   t_7820,   t_7821;
/* u2_2683 Output nets */
wire t_7822,   t_7823,   t_7824;
/* u2_2684 Output nets */
wire t_7825,   t_7826,   t_7827;
/* u2_2685 Output nets */
wire t_7828,   t_7829,   t_7830;
/* u2_2686 Output nets */
wire t_7831,   t_7832,   t_7833;
/* u2_2687 Output nets */
wire t_7834,   t_7835,   t_7836;
/* u1_2688 Output nets */
wire t_7837,   t_7838;
/* u2_2689 Output nets */
wire t_7839,   t_7840,   t_7841;
/* u2_2690 Output nets */
wire t_7842,   t_7843,   t_7844;
/* u2_2691 Output nets */
wire t_7845,   t_7846,   t_7847;
/* u2_2692 Output nets */
wire t_7848,   t_7849,   t_7850;
/* u2_2693 Output nets */
wire t_7851,   t_7852,   t_7853;
/* u2_2694 Output nets */
wire t_7854,   t_7855,   t_7856;
/* u2_2695 Output nets */
wire t_7857,   t_7858,   t_7859;
/* u2_2696 Output nets */
wire t_7860,   t_7861,   t_7862;
/* u2_2697 Output nets */
wire t_7863,   t_7864,   t_7865;
/* u2_2698 Output nets */
wire t_7866,   t_7867,   t_7868;
/* u2_2699 Output nets */
wire t_7869,   t_7870,   t_7871;
/* u2_2700 Output nets */
wire t_7872,   t_7873,   t_7874;
/* u2_2701 Output nets */
wire t_7875,   t_7876,   t_7877;
/* u2_2702 Output nets */
wire t_7878,   t_7879,   t_7880;
/* u2_2703 Output nets */
wire t_7881,   t_7882,   t_7883;
/* u2_2704 Output nets */
wire t_7884,   t_7885,   t_7886;
/* u2_2705 Output nets */
wire t_7887,   t_7888,   t_7889;
/* u2_2706 Output nets */
wire t_7890,   t_7891,   t_7892;
/* u2_2707 Output nets */
wire t_7893,   t_7894,   t_7895;
/* u2_2708 Output nets */
wire t_7896,   t_7897,   t_7898;
/* u2_2709 Output nets */
wire t_7899,   t_7900,   t_7901;
/* u2_2710 Output nets */
wire t_7902,   t_7903,   t_7904;
/* u2_2711 Output nets */
wire t_7905,   t_7906,   t_7907;
/* u2_2712 Output nets */
wire t_7908,   t_7909,   t_7910;
/* u2_2713 Output nets */
wire t_7911,   t_7912,   t_7913;
/* u2_2714 Output nets */
wire t_7914,   t_7915,   t_7916;
/* u2_2715 Output nets */
wire t_7917,   t_7918,   t_7919;
/* u2_2716 Output nets */
wire t_7920,   t_7921,   t_7922;
/* u2_2717 Output nets */
wire t_7923,   t_7924,   t_7925;
/* u2_2718 Output nets */
wire t_7926,   t_7927,   t_7928;
/* u2_2719 Output nets */
wire t_7929,   t_7930,   t_7931;
/* u2_2720 Output nets */
wire t_7932,   t_7933,   t_7934;
/* u2_2721 Output nets */
wire t_7935,   t_7936,   t_7937;
/* u2_2722 Output nets */
wire t_7938,   t_7939,   t_7940;
/* u2_2723 Output nets */
wire t_7941,   t_7942,   t_7943;
/* u2_2724 Output nets */
wire t_7944,   t_7945,   t_7946;
/* u2_2725 Output nets */
wire t_7947,   t_7948,   t_7949;
/* u2_2726 Output nets */
wire t_7950,   t_7951,   t_7952;
/* u2_2727 Output nets */
wire t_7953,   t_7954,   t_7955;
/* u2_2728 Output nets */
wire t_7956,   t_7957,   t_7958;
/* u2_2729 Output nets */
wire t_7959,   t_7960,   t_7961;
/* u2_2730 Output nets */
wire t_7962,   t_7963,   t_7964;
/* u2_2731 Output nets */
wire t_7965,   t_7966,   t_7967;
/* u2_2732 Output nets */
wire t_7968,   t_7969,   t_7970;
/* u2_2733 Output nets */
wire t_7971,   t_7972,   t_7973;
/* u2_2734 Output nets */
wire t_7974,   t_7975,   t_7976;
/* u2_2735 Output nets */
wire t_7977,   t_7978,   t_7979;
/* u2_2736 Output nets */
wire t_7980,   t_7981,   t_7982;
/* u2_2737 Output nets */
wire t_7983,   t_7984,   t_7985;
/* u2_2738 Output nets */
wire t_7986,   t_7987,   t_7988;
/* u2_2739 Output nets */
wire t_7989,   t_7990,   t_7991;
/* u2_2740 Output nets */
wire t_7992,   t_7993,   t_7994;
/* u2_2741 Output nets */
wire t_7995,   t_7996,   t_7997;
/* u2_2742 Output nets */
wire t_7998,   t_7999,   t_8000;
/* u2_2743 Output nets */
wire t_8001,   t_8002,   t_8003;
/* u2_2744 Output nets */
wire t_8004,   t_8005,   t_8006;
/* u2_2745 Output nets */
wire t_8007,   t_8008,   t_8009;
/* u2_2746 Output nets */
wire t_8010,   t_8011,   t_8012;
/* u2_2747 Output nets */
wire t_8013,   t_8014,   t_8015;
/* u2_2748 Output nets */
wire t_8016,   t_8017,   t_8018;
/* u2_2749 Output nets */
wire t_8019,   t_8020,   t_8021;
/* u2_2750 Output nets */
wire t_8022,   t_8023,   t_8024;
/* u2_2751 Output nets */
wire t_8025,   t_8026,   t_8027;
/* u2_2752 Output nets */
wire t_8028,   t_8029,   t_8030;
/* u2_2753 Output nets */
wire t_8031,   t_8032,   t_8033;
/* u2_2754 Output nets */
wire t_8034,   t_8035,   t_8036;
/* u2_2755 Output nets */
wire t_8037,   t_8038,   t_8039;
/* u2_2756 Output nets */
wire t_8040,   t_8041,   t_8042;
/* u2_2757 Output nets */
wire t_8043,   t_8044,   t_8045;
/* u2_2758 Output nets */
wire t_8046,   t_8047,   t_8048;
/* u2_2759 Output nets */
wire t_8049,   t_8050,   t_8051;
/* u2_2760 Output nets */
wire t_8052,   t_8053,   t_8054;
/* u2_2761 Output nets */
wire t_8055,   t_8056,   t_8057;
/* u2_2762 Output nets */
wire t_8058,   t_8059,   t_8060;
/* u2_2763 Output nets */
wire t_8061,   t_8062,   t_8063;
/* u2_2764 Output nets */
wire t_8064,   t_8065,   t_8066;
/* u2_2765 Output nets */
wire t_8067,   t_8068,   t_8069;
/* u2_2766 Output nets */
wire t_8070,   t_8071,   t_8072;
/* u2_2767 Output nets */
wire t_8073,   t_8074,   t_8075;
/* u2_2768 Output nets */
wire t_8076,   t_8077,   t_8078;
/* u2_2769 Output nets */
wire t_8079,   t_8080,   t_8081;
/* u2_2770 Output nets */
wire t_8082,   t_8083,   t_8084;
/* u2_2771 Output nets */
wire t_8085,   t_8086,   t_8087;
/* u2_2772 Output nets */
wire t_8088,   t_8089,   t_8090;
/* u2_2773 Output nets */
wire t_8091,   t_8092,   t_8093;
/* u2_2774 Output nets */
wire t_8094,   t_8095,   t_8096;
/* u2_2775 Output nets */
wire t_8097,   t_8098,   t_8099;
/* u2_2776 Output nets */
wire t_8100,   t_8101,   t_8102;
/* u2_2777 Output nets */
wire t_8103,   t_8104,   t_8105;
/* u2_2778 Output nets */
wire t_8106,   t_8107,   t_8108;
/* u2_2779 Output nets */
wire t_8109,   t_8110,   t_8111;
/* u2_2780 Output nets */
wire t_8112,   t_8113,   t_8114;
/* u2_2781 Output nets */
wire t_8115,   t_8116,   t_8117;
/* u2_2782 Output nets */
wire t_8118,   t_8119,   t_8120;
/* u2_2783 Output nets */
wire t_8121,   t_8122,   t_8123;
/* u2_2784 Output nets */
wire t_8124,   t_8125,   t_8126;
/* u2_2785 Output nets */
wire t_8127,   t_8128,   t_8129;
/* u2_2786 Output nets */
wire t_8130,   t_8131,   t_8132;
/* u2_2787 Output nets */
wire t_8133,   t_8134,   t_8135;
/* u2_2788 Output nets */
wire t_8136,   t_8137,   t_8138;
/* u2_2789 Output nets */
wire t_8139,   t_8140,   t_8141;
/* u2_2790 Output nets */
wire t_8142,   t_8143,   t_8144;
/* u2_2791 Output nets */
wire t_8145,   t_8146,   t_8147;
/* u2_2792 Output nets */
wire t_8148,   t_8149,   t_8150;
/* u2_2793 Output nets */
wire t_8151,   t_8152,   t_8153;
/* u2_2794 Output nets */
wire t_8154,   t_8155,   t_8156;
/* u2_2795 Output nets */
wire t_8157,   t_8158,   t_8159;
/* u2_2796 Output nets */
wire t_8160,   t_8161,   t_8162;
/* u2_2797 Output nets */
wire t_8163,   t_8164,   t_8165;
/* u2_2798 Output nets */
wire t_8166,   t_8167,   t_8168;
/* u2_2799 Output nets */
wire t_8169,   t_8170,   t_8171;
/* u1_2800 Output nets */
wire t_8172,   t_8173;
/* u2_2801 Output nets */
wire t_8174,   t_8175,   t_8176;
/* u2_2802 Output nets */
wire t_8177,   t_8178,   t_8179;
/* u2_2803 Output nets */
wire t_8180,   t_8181,   t_8182;
/* u2_2804 Output nets */
wire t_8183,   t_8184,   t_8185;
/* u2_2805 Output nets */
wire t_8186,   t_8187,   t_8188;
/* u2_2806 Output nets */
wire t_8189,   t_8190,   t_8191;
/* u2_2807 Output nets */
wire t_8192,   t_8193,   t_8194;
/* u0_2808 Output nets */
wire t_8195,   t_8196;
/* u2_2809 Output nets */
wire t_8197,   t_8198,   t_8199;
/* u2_2810 Output nets */
wire t_8200,   t_8201,   t_8202;
/* u2_2811 Output nets */
wire t_8203,   t_8204,   t_8205;
/* u2_2812 Output nets */
wire t_8206,   t_8207,   t_8208;
/* u2_2813 Output nets */
wire t_8209,   t_8210,   t_8211;
/* u2_2814 Output nets */
wire t_8212,   t_8213,   t_8214;
/* u2_2815 Output nets */
wire t_8215,   t_8216,   t_8217;
/* u0_2816 Output nets */
wire t_8218,   t_8219;
/* u2_2817 Output nets */
wire t_8220,   t_8221,   t_8222;
/* u2_2818 Output nets */
wire t_8223,   t_8224,   t_8225;
/* u2_2819 Output nets */
wire t_8226,   t_8227,   t_8228;
/* u2_2820 Output nets */
wire t_8229,   t_8230,   t_8231;
/* u2_2821 Output nets */
wire t_8232,   t_8233,   t_8234;
/* u2_2822 Output nets */
wire t_8235,   t_8236,   t_8237;
/* u2_2823 Output nets */
wire t_8238,   t_8239,   t_8240;
/* u1_2824 Output nets */
wire t_8241,   t_8242;
/* u2_2825 Output nets */
wire t_8243,   t_8244,   t_8245;
/* u2_2826 Output nets */
wire t_8246,   t_8247,   t_8248;
/* u2_2827 Output nets */
wire t_8249,   t_8250,   t_8251;
/* u2_2828 Output nets */
wire t_8252,   t_8253,   t_8254;
/* u2_2829 Output nets */
wire t_8255,   t_8256,   t_8257;
/* u2_2830 Output nets */
wire t_8258,   t_8259,   t_8260;
/* u2_2831 Output nets */
wire t_8261,   t_8262,   t_8263;
/* u0_2832 Output nets */
wire t_8264,   t_8265;
/* u2_2833 Output nets */
wire t_8266,   t_8267,   t_8268;
/* u2_2834 Output nets */
wire t_8269,   t_8270,   t_8271;
/* u2_2835 Output nets */
wire t_8272,   t_8273,   t_8274;
/* u2_2836 Output nets */
wire t_8275,   t_8276,   t_8277;
/* u2_2837 Output nets */
wire t_8278,   t_8279,   t_8280;
/* u2_2838 Output nets */
wire t_8281,   t_8282,   t_8283;
/* u2_2839 Output nets */
wire t_8284,   t_8285,   t_8286;
/* u0_2840 Output nets */
wire t_8287,   t_8288;
/* u2_2841 Output nets */
wire t_8289,   t_8290,   t_8291;
/* u2_2842 Output nets */
wire t_8292,   t_8293,   t_8294;
/* u2_2843 Output nets */
wire t_8295,   t_8296,   t_8297;
/* u2_2844 Output nets */
wire t_8298,   t_8299,   t_8300;
/* u2_2845 Output nets */
wire t_8301,   t_8302,   t_8303;
/* u2_2846 Output nets */
wire t_8304,   t_8305,   t_8306;
/* u2_2847 Output nets */
wire t_8307,   t_8308,   t_8309;
/* u0_2848 Output nets */
wire t_8310,   t_8311;
/* u2_2849 Output nets */
wire t_8312,   t_8313,   t_8314;
/* u2_2850 Output nets */
wire t_8315,   t_8316,   t_8317;
/* u2_2851 Output nets */
wire t_8318,   t_8319,   t_8320;
/* u2_2852 Output nets */
wire t_8321,   t_8322,   t_8323;
/* u2_2853 Output nets */
wire t_8324,   t_8325,   t_8326;
/* u2_2854 Output nets */
wire t_8327,   t_8328,   t_8329;
/* u2_2855 Output nets */
wire t_8330,   t_8331,   t_8332;
/* u0_2856 Output nets */
wire t_8333,   t_8334;
/* u2_2857 Output nets */
wire t_8335,   t_8336,   t_8337;
/* u2_2858 Output nets */
wire t_8338,   t_8339,   t_8340;
/* u2_2859 Output nets */
wire t_8341,   t_8342,   t_8343;
/* u2_2860 Output nets */
wire t_8344,   t_8345,   t_8346;
/* u2_2861 Output nets */
wire t_8347,   t_8348,   t_8349;
/* u2_2862 Output nets */
wire t_8350,   t_8351,   t_8352;
/* u2_2863 Output nets */
wire t_8353,   t_8354,   t_8355;
/* u2_2864 Output nets */
wire t_8356,   t_8357,   t_8358;
/* u2_2865 Output nets */
wire t_8359,   t_8360,   t_8361;
/* u2_2866 Output nets */
wire t_8362,   t_8363,   t_8364;
/* u2_2867 Output nets */
wire t_8365,   t_8366,   t_8367;
/* u2_2868 Output nets */
wire t_8368,   t_8369,   t_8370;
/* u2_2869 Output nets */
wire t_8371,   t_8372,   t_8373;
/* u2_2870 Output nets */
wire t_8374,   t_8375,   t_8376;
/* u2_2871 Output nets */
wire t_8377,   t_8378,   t_8379;
/* u2_2872 Output nets */
wire t_8380,   t_8381,   t_8382;
/* u2_2873 Output nets */
wire t_8383,   t_8384,   t_8385;
/* u2_2874 Output nets */
wire t_8386,   t_8387,   t_8388;
/* u2_2875 Output nets */
wire t_8389,   t_8390,   t_8391;
/* u2_2876 Output nets */
wire t_8392,   t_8393,   t_8394;
/* u2_2877 Output nets */
wire t_8395,   t_8396,   t_8397;
/* u2_2878 Output nets */
wire t_8398,   t_8399,   t_8400;
/* u2_2879 Output nets */
wire t_8401,   t_8402,   t_8403;
/* u2_2880 Output nets */
wire t_8404,   t_8405,   t_8406;
/* u2_2881 Output nets */
wire t_8407,   t_8408,   t_8409;
/* u2_2882 Output nets */
wire t_8410,   t_8411,   t_8412;
/* u2_2883 Output nets */
wire t_8413,   t_8414,   t_8415;
/* u2_2884 Output nets */
wire t_8416,   t_8417,   t_8418;
/* u2_2885 Output nets */
wire t_8419,   t_8420,   t_8421;
/* u2_2886 Output nets */
wire t_8422,   t_8423,   t_8424;
/* u2_2887 Output nets */
wire t_8425,   t_8426,   t_8427;
/* u2_2888 Output nets */
wire t_8428,   t_8429,   t_8430;
/* u2_2889 Output nets */
wire t_8431,   t_8432,   t_8433;
/* u2_2890 Output nets */
wire t_8434,   t_8435,   t_8436;
/* u2_2891 Output nets */
wire t_8437,   t_8438,   t_8439;
/* u2_2892 Output nets */
wire t_8440,   t_8441,   t_8442;
/* u2_2893 Output nets */
wire t_8443,   t_8444,   t_8445;
/* u2_2894 Output nets */
wire t_8446,   t_8447,   t_8448;
/* u2_2895 Output nets */
wire t_8449,   t_8450,   t_8451;
/* u2_2896 Output nets */
wire t_8452,   t_8453,   t_8454;
/* u2_2897 Output nets */
wire t_8455,   t_8456,   t_8457;
/* u2_2898 Output nets */
wire t_8458,   t_8459,   t_8460;
/* u2_2899 Output nets */
wire t_8461,   t_8462,   t_8463;
/* u2_2900 Output nets */
wire t_8464,   t_8465,   t_8466;
/* u2_2901 Output nets */
wire t_8467,   t_8468,   t_8469;
/* u2_2902 Output nets */
wire t_8470,   t_8471,   t_8472;
/* u2_2903 Output nets */
wire t_8473,   t_8474,   t_8475;
/* u2_2904 Output nets */
wire t_8476,   t_8477,   t_8478;
/* u2_2905 Output nets */
wire t_8479,   t_8480,   t_8481;
/* u2_2906 Output nets */
wire t_8482,   t_8483,   t_8484;
/* u2_2907 Output nets */
wire t_8485,   t_8486,   t_8487;
/* u2_2908 Output nets */
wire t_8488,   t_8489,   t_8490;
/* u2_2909 Output nets */
wire t_8491,   t_8492,   t_8493;
/* u2_2910 Output nets */
wire t_8494,   t_8495,   t_8496;
/* u2_2911 Output nets */
wire t_8497,   t_8498,   t_8499;
/* u2_2912 Output nets */
wire t_8500,   t_8501,   t_8502;
/* u2_2913 Output nets */
wire t_8503,   t_8504,   t_8505;
/* u2_2914 Output nets */
wire t_8506,   t_8507,   t_8508;
/* u2_2915 Output nets */
wire t_8509,   t_8510,   t_8511;
/* u2_2916 Output nets */
wire t_8512,   t_8513,   t_8514;
/* u2_2917 Output nets */
wire t_8515,   t_8516,   t_8517;
/* u2_2918 Output nets */
wire t_8518,   t_8519,   t_8520;
/* u1_2919 Output nets */
wire t_8521,   t_8522;
/* u2_2920 Output nets */
wire t_8523,   t_8524,   t_8525;
/* u2_2921 Output nets */
wire t_8526,   t_8527,   t_8528;
/* u2_2922 Output nets */
wire t_8529,   t_8530,   t_8531;
/* u2_2923 Output nets */
wire t_8532,   t_8533,   t_8534;
/* u2_2924 Output nets */
wire t_8535,   t_8536,   t_8537;
/* u2_2925 Output nets */
wire t_8538,   t_8539,   t_8540;
/* u0_2926 Output nets */
wire t_8541,   t_8542;
/* u2_2927 Output nets */
wire t_8543,   t_8544,   t_8545;
/* u2_2928 Output nets */
wire t_8546,   t_8547,   t_8548;
/* u2_2929 Output nets */
wire t_8549,   t_8550,   t_8551;
/* u2_2930 Output nets */
wire t_8552,   t_8553,   t_8554;
/* u2_2931 Output nets */
wire t_8555,   t_8556,   t_8557;
/* u2_2932 Output nets */
wire t_8558,   t_8559,   t_8560;
/* u0_2933 Output nets */
wire t_8561,   t_8562;
/* u2_2934 Output nets */
wire t_8563,   t_8564,   t_8565;
/* u2_2935 Output nets */
wire t_8566,   t_8567,   t_8568;
/* u2_2936 Output nets */
wire t_8569,   t_8570,   t_8571;
/* u2_2937 Output nets */
wire t_8572,   t_8573,   t_8574;
/* u2_2938 Output nets */
wire t_8575,   t_8576,   t_8577;
/* u2_2939 Output nets */
wire t_8578,   t_8579,   t_8580;
/* u1_2940 Output nets */
wire t_8581,   t_8582;
/* u2_2941 Output nets */
wire t_8583,   t_8584,   t_8585;
/* u2_2942 Output nets */
wire t_8586,   t_8587,   t_8588;
/* u2_2943 Output nets */
wire t_8589,   t_8590,   t_8591;
/* u2_2944 Output nets */
wire t_8592,   t_8593,   t_8594;
/* u2_2945 Output nets */
wire t_8595,   t_8596,   t_8597;
/* u2_2946 Output nets */
wire t_8598,   t_8599,   t_8600;
/* u0_2947 Output nets */
wire t_8601,   t_8602;
/* u2_2948 Output nets */
wire t_8603,   t_8604,   t_8605;
/* u2_2949 Output nets */
wire t_8606,   t_8607,   t_8608;
/* u2_2950 Output nets */
wire t_8609,   t_8610,   t_8611;
/* u2_2951 Output nets */
wire t_8612,   t_8613,   t_8614;
/* u2_2952 Output nets */
wire t_8615,   t_8616,   t_8617;
/* u2_2953 Output nets */
wire t_8618,   t_8619,   t_8620;
/* u0_2954 Output nets */
wire t_8621,   t_8622;
/* u2_2955 Output nets */
wire t_8623,   t_8624,   t_8625;
/* u2_2956 Output nets */
wire t_8626,   t_8627,   t_8628;
/* u2_2957 Output nets */
wire t_8629,   t_8630,   t_8631;
/* u2_2958 Output nets */
wire t_8632,   t_8633,   t_8634;
/* u2_2959 Output nets */
wire t_8635,   t_8636,   t_8637;
/* u2_2960 Output nets */
wire t_8638,   t_8639,   t_8640;
/* u0_2961 Output nets */
wire t_8641,   t_8642;
/* u2_2962 Output nets */
wire t_8643,   t_8644,   t_8645;
/* u2_2963 Output nets */
wire t_8646,   t_8647,   t_8648;
/* u2_2964 Output nets */
wire t_8649,   t_8650,   t_8651;
/* u2_2965 Output nets */
wire t_8652,   t_8653,   t_8654;
/* u2_2966 Output nets */
wire t_8655,   t_8656,   t_8657;
/* u2_2967 Output nets */
wire t_8658,   t_8659,   t_8660;
/* u0_2968 Output nets */
wire t_8661,   t_8662;
/* u2_2969 Output nets */
wire t_8663,   t_8664,   t_8665;
/* u2_2970 Output nets */
wire t_8666,   t_8667,   t_8668;
/* u2_2971 Output nets */
wire t_8669,   t_8670,   t_8671;
/* u2_2972 Output nets */
wire t_8672,   t_8673,   t_8674;
/* u2_2973 Output nets */
wire t_8675,   t_8676,   t_8677;
/* u2_2974 Output nets */
wire t_8678,   t_8679,   t_8680;
/* u2_2975 Output nets */
wire t_8681,   t_8682,   t_8683;
/* u2_2976 Output nets */
wire t_8684,   t_8685,   t_8686;
/* u2_2977 Output nets */
wire t_8687,   t_8688,   t_8689;
/* u2_2978 Output nets */
wire t_8690,   t_8691,   t_8692;
/* u2_2979 Output nets */
wire t_8693,   t_8694,   t_8695;
/* u2_2980 Output nets */
wire t_8696,   t_8697,   t_8698;
/* u2_2981 Output nets */
wire t_8699,   t_8700,   t_8701;
/* u2_2982 Output nets */
wire t_8702,   t_8703,   t_8704;
/* u2_2983 Output nets */
wire t_8705,   t_8706,   t_8707;
/* u2_2984 Output nets */
wire t_8708,   t_8709,   t_8710;
/* u2_2985 Output nets */
wire t_8711,   t_8712,   t_8713;
/* u2_2986 Output nets */
wire t_8714,   t_8715,   t_8716;
/* u2_2987 Output nets */
wire t_8717,   t_8718,   t_8719;
/* u2_2988 Output nets */
wire t_8720,   t_8721,   t_8722;
/* u2_2989 Output nets */
wire t_8723,   t_8724,   t_8725;
/* u2_2990 Output nets */
wire t_8726,   t_8727,   t_8728;
/* u2_2991 Output nets */
wire t_8729,   t_8730,   t_8731;
/* u2_2992 Output nets */
wire t_8732,   t_8733,   t_8734;
/* u2_2993 Output nets */
wire t_8735,   t_8736,   t_8737;
/* u2_2994 Output nets */
wire t_8738,   t_8739,   t_8740;
/* u2_2995 Output nets */
wire t_8741,   t_8742,   t_8743;
/* u2_2996 Output nets */
wire t_8744,   t_8745,   t_8746;
/* u2_2997 Output nets */
wire t_8747,   t_8748,   t_8749;
/* u2_2998 Output nets */
wire t_8750,   t_8751,   t_8752;
/* u2_2999 Output nets */
wire t_8753,   t_8754,   t_8755;
/* u2_3000 Output nets */
wire t_8756,   t_8757,   t_8758;
/* u2_3001 Output nets */
wire t_8759,   t_8760,   t_8761;
/* u2_3002 Output nets */
wire t_8762,   t_8763,   t_8764;
/* u2_3003 Output nets */
wire t_8765,   t_8766,   t_8767;
/* u2_3004 Output nets */
wire t_8768,   t_8769,   t_8770;
/* u2_3005 Output nets */
wire t_8771,   t_8772,   t_8773;
/* u2_3006 Output nets */
wire t_8774,   t_8775,   t_8776;
/* u2_3007 Output nets */
wire t_8777,   t_8778,   t_8779;
/* u2_3008 Output nets */
wire t_8780,   t_8781,   t_8782;
/* u2_3009 Output nets */
wire t_8783,   t_8784,   t_8785;
/* u2_3010 Output nets */
wire t_8786,   t_8787,   t_8788;
/* u2_3011 Output nets */
wire t_8789,   t_8790,   t_8791;
/* u2_3012 Output nets */
wire t_8792,   t_8793,   t_8794;
/* u2_3013 Output nets */
wire t_8795,   t_8796,   t_8797;
/* u2_3014 Output nets */
wire t_8798,   t_8799,   t_8800;
/* u2_3015 Output nets */
wire t_8801,   t_8802,   t_8803;
/* u2_3016 Output nets */
wire t_8804,   t_8805,   t_8806;
/* u2_3017 Output nets */
wire t_8807,   t_8808,   t_8809;
/* u2_3018 Output nets */
wire t_8810,   t_8811,   t_8812;
/* u2_3019 Output nets */
wire t_8813,   t_8814,   t_8815;
/* u2_3020 Output nets */
wire t_8816,   t_8817,   t_8818;
/* u2_3021 Output nets */
wire t_8819,   t_8820,   t_8821;
/* u1_3022 Output nets */
wire t_8822,   t_8823;
/* u2_3023 Output nets */
wire t_8824,   t_8825,   t_8826;
/* u2_3024 Output nets */
wire t_8827,   t_8828,   t_8829;
/* u2_3025 Output nets */
wire t_8830,   t_8831,   t_8832;
/* u2_3026 Output nets */
wire t_8833,   t_8834,   t_8835;
/* u2_3027 Output nets */
wire t_8836,   t_8837,   t_8838;
/* u0_3028 Output nets */
wire t_8839,   t_8840;
/* u2_3029 Output nets */
wire t_8841,   t_8842,   t_8843;
/* u2_3030 Output nets */
wire t_8844,   t_8845,   t_8846;
/* u2_3031 Output nets */
wire t_8847,   t_8848,   t_8849;
/* u2_3032 Output nets */
wire t_8850,   t_8851,   t_8852;
/* u2_3033 Output nets */
wire t_8853,   t_8854,   t_8855;
/* u0_3034 Output nets */
wire t_8856,   t_8857;
/* u2_3035 Output nets */
wire t_8858,   t_8859,   t_8860;
/* u2_3036 Output nets */
wire t_8861,   t_8862,   t_8863;
/* u2_3037 Output nets */
wire t_8864,   t_8865,   t_8866;
/* u2_3038 Output nets */
wire t_8867,   t_8868,   t_8869;
/* u2_3039 Output nets */
wire t_8870,   t_8871,   t_8872;
/* u1_3040 Output nets */
wire t_8873,   t_8874;
/* u2_3041 Output nets */
wire t_8875,   t_8876,   t_8877;
/* u2_3042 Output nets */
wire t_8878,   t_8879,   t_8880;
/* u2_3043 Output nets */
wire t_8881,   t_8882,   t_8883;
/* u2_3044 Output nets */
wire t_8884,   t_8885,   t_8886;
/* u2_3045 Output nets */
wire t_8887,   t_8888,   t_8889;
/* u0_3046 Output nets */
wire t_8890,   t_8891;
/* u2_3047 Output nets */
wire t_8892,   t_8893,   t_8894;
/* u2_3048 Output nets */
wire t_8895,   t_8896,   t_8897;
/* u2_3049 Output nets */
wire t_8898,   t_8899,   t_8900;
/* u2_3050 Output nets */
wire t_8901,   t_8902,   t_8903;
/* u2_3051 Output nets */
wire t_8904,   t_8905,   t_8906;
/* u0_3052 Output nets */
wire t_8907,   t_8908;
/* u2_3053 Output nets */
wire t_8909,   t_8910,   t_8911;
/* u2_3054 Output nets */
wire t_8912,   t_8913,   t_8914;
/* u2_3055 Output nets */
wire t_8915,   t_8916,   t_8917;
/* u2_3056 Output nets */
wire t_8918,   t_8919,   t_8920;
/* u2_3057 Output nets */
wire t_8921,   t_8922,   t_8923;
/* u0_3058 Output nets */
wire t_8924,   t_8925;
/* u2_3059 Output nets */
wire t_8926,   t_8927,   t_8928;
/* u2_3060 Output nets */
wire t_8929,   t_8930,   t_8931;
/* u2_3061 Output nets */
wire t_8932,   t_8933,   t_8934;
/* u2_3062 Output nets */
wire t_8935,   t_8936,   t_8937;
/* u2_3063 Output nets */
wire t_8938,   t_8939,   t_8940;
/* u0_3064 Output nets */
wire t_8941,   t_8942;
/* u2_3065 Output nets */
wire t_8943,   t_8944,   t_8945;
/* u2_3066 Output nets */
wire t_8946,   t_8947,   t_8948;
/* u2_3067 Output nets */
wire t_8949,   t_8950,   t_8951;
/* u2_3068 Output nets */
wire t_8952,   t_8953,   t_8954;
/* u2_3069 Output nets */
wire t_8955,   t_8956,   t_8957;
/* u2_3070 Output nets */
wire t_8958,   t_8959,   t_8960;
/* u2_3071 Output nets */
wire t_8961,   t_8962,   t_8963;
/* u2_3072 Output nets */
wire t_8964,   t_8965,   t_8966;
/* u2_3073 Output nets */
wire t_8967,   t_8968,   t_8969;
/* u2_3074 Output nets */
wire t_8970,   t_8971,   t_8972;
/* u2_3075 Output nets */
wire t_8973,   t_8974,   t_8975;
/* u2_3076 Output nets */
wire t_8976,   t_8977,   t_8978;
/* u2_3077 Output nets */
wire t_8979,   t_8980,   t_8981;
/* u2_3078 Output nets */
wire t_8982,   t_8983,   t_8984;
/* u2_3079 Output nets */
wire t_8985,   t_8986,   t_8987;
/* u2_3080 Output nets */
wire t_8988,   t_8989,   t_8990;
/* u2_3081 Output nets */
wire t_8991,   t_8992,   t_8993;
/* u2_3082 Output nets */
wire t_8994,   t_8995,   t_8996;
/* u2_3083 Output nets */
wire t_8997,   t_8998,   t_8999;
/* u2_3084 Output nets */
wire t_9000,   t_9001,   t_9002;
/* u2_3085 Output nets */
wire t_9003,   t_9004,   t_9005;
/* u2_3086 Output nets */
wire t_9006,   t_9007,   t_9008;
/* u2_3087 Output nets */
wire t_9009,   t_9010,   t_9011;
/* u2_3088 Output nets */
wire t_9012,   t_9013,   t_9014;
/* u2_3089 Output nets */
wire t_9015,   t_9016,   t_9017;
/* u2_3090 Output nets */
wire t_9018,   t_9019,   t_9020;
/* u2_3091 Output nets */
wire t_9021,   t_9022,   t_9023;
/* u2_3092 Output nets */
wire t_9024,   t_9025,   t_9026;
/* u2_3093 Output nets */
wire t_9027,   t_9028,   t_9029;
/* u2_3094 Output nets */
wire t_9030,   t_9031,   t_9032;
/* u2_3095 Output nets */
wire t_9033,   t_9034,   t_9035;
/* u2_3096 Output nets */
wire t_9036,   t_9037,   t_9038;
/* u2_3097 Output nets */
wire t_9039,   t_9040,   t_9041;
/* u2_3098 Output nets */
wire t_9042,   t_9043,   t_9044;
/* u2_3099 Output nets */
wire t_9045,   t_9046,   t_9047;
/* u2_3100 Output nets */
wire t_9048,   t_9049,   t_9050;
/* u2_3101 Output nets */
wire t_9051,   t_9052,   t_9053;
/* u2_3102 Output nets */
wire t_9054,   t_9055,   t_9056;
/* u2_3103 Output nets */
wire t_9057,   t_9058,   t_9059;
/* u2_3104 Output nets */
wire t_9060,   t_9061,   t_9062;
/* u2_3105 Output nets */
wire t_9063,   t_9064,   t_9065;
/* u2_3106 Output nets */
wire t_9066,   t_9067,   t_9068;
/* u2_3107 Output nets */
wire t_9069,   t_9070,   t_9071;
/* u2_3108 Output nets */
wire t_9072,   t_9073,   t_9074;
/* u1_3109 Output nets */
wire t_9075,   t_9076;
/* u2_3110 Output nets */
wire t_9077,   t_9078,   t_9079;
/* u2_3111 Output nets */
wire t_9080,   t_9081,   t_9082;
/* u2_3112 Output nets */
wire t_9083,   t_9084,   t_9085;
/* u2_3113 Output nets */
wire t_9086,   t_9087,   t_9088;
/* u0_3114 Output nets */
wire t_9089,   t_9090;
/* u2_3115 Output nets */
wire t_9091,   t_9092,   t_9093;
/* u2_3116 Output nets */
wire t_9094,   t_9095,   t_9096;
/* u2_3117 Output nets */
wire t_9097,   t_9098,   t_9099;
/* u2_3118 Output nets */
wire t_9100,   t_9101,   t_9102;
/* u0_3119 Output nets */
wire t_9103,   t_9104;
/* u2_3120 Output nets */
wire t_9105,   t_9106,   t_9107;
/* u2_3121 Output nets */
wire t_9108,   t_9109,   t_9110;
/* u2_3122 Output nets */
wire t_9111,   t_9112,   t_9113;
/* u2_3123 Output nets */
wire t_9114,   t_9115,   t_9116;
/* u1_3124 Output nets */
wire t_9117,   t_9118;
/* u2_3125 Output nets */
wire t_9119,   t_9120,   t_9121;
/* u2_3126 Output nets */
wire t_9122,   t_9123,   t_9124;
/* u2_3127 Output nets */
wire t_9125,   t_9126,   t_9127;
/* u2_3128 Output nets */
wire t_9128,   t_9129,   t_9130;
/* u0_3129 Output nets */
wire t_9131,   t_9132;
/* u2_3130 Output nets */
wire t_9133,   t_9134,   t_9135;
/* u2_3131 Output nets */
wire t_9136,   t_9137,   t_9138;
/* u2_3132 Output nets */
wire t_9139,   t_9140,   t_9141;
/* u2_3133 Output nets */
wire t_9142,   t_9143,   t_9144;
/* u0_3134 Output nets */
wire t_9145,   t_9146;
/* u2_3135 Output nets */
wire t_9147,   t_9148,   t_9149;
/* u2_3136 Output nets */
wire t_9150,   t_9151,   t_9152;
/* u2_3137 Output nets */
wire t_9153,   t_9154,   t_9155;
/* u2_3138 Output nets */
wire t_9156,   t_9157,   t_9158;
/* u0_3139 Output nets */
wire t_9159,   t_9160;
/* u2_3140 Output nets */
wire t_9161,   t_9162,   t_9163;
/* u2_3141 Output nets */
wire t_9164,   t_9165,   t_9166;
/* u2_3142 Output nets */
wire t_9167,   t_9168,   t_9169;
/* u2_3143 Output nets */
wire t_9170,   t_9171,   t_9172;
/* u0_3144 Output nets */
wire t_9173,   t_9174;
/* u2_3145 Output nets */
wire t_9175,   t_9176,   t_9177;
/* u2_3146 Output nets */
wire t_9178,   t_9179,   t_9180;
/* u2_3147 Output nets */
wire t_9181,   t_9182,   t_9183;
/* u2_3148 Output nets */
wire t_9184,   t_9185,   t_9186;
/* u2_3149 Output nets */
wire t_9187,   t_9188,   t_9189;
/* u2_3150 Output nets */
wire t_9190,   t_9191,   t_9192;
/* u2_3151 Output nets */
wire t_9193,   t_9194,   t_9195;
/* u2_3152 Output nets */
wire t_9196,   t_9197,   t_9198;
/* u2_3153 Output nets */
wire t_9199,   t_9200,   t_9201;
/* u2_3154 Output nets */
wire t_9202,   t_9203,   t_9204;
/* u2_3155 Output nets */
wire t_9205,   t_9206,   t_9207;
/* u2_3156 Output nets */
wire t_9208,   t_9209,   t_9210;
/* u2_3157 Output nets */
wire t_9211,   t_9212,   t_9213;
/* u2_3158 Output nets */
wire t_9214,   t_9215,   t_9216;
/* u2_3159 Output nets */
wire t_9217,   t_9218,   t_9219;
/* u2_3160 Output nets */
wire t_9220,   t_9221,   t_9222;
/* u2_3161 Output nets */
wire t_9223,   t_9224,   t_9225;
/* u2_3162 Output nets */
wire t_9226,   t_9227,   t_9228;
/* u2_3163 Output nets */
wire t_9229,   t_9230,   t_9231;
/* u2_3164 Output nets */
wire t_9232,   t_9233,   t_9234;
/* u2_3165 Output nets */
wire t_9235,   t_9236,   t_9237;
/* u2_3166 Output nets */
wire t_9238,   t_9239,   t_9240;
/* u2_3167 Output nets */
wire t_9241,   t_9242,   t_9243;
/* u2_3168 Output nets */
wire t_9244,   t_9245,   t_9246;
/* u2_3169 Output nets */
wire t_9247,   t_9248,   t_9249;
/* u2_3170 Output nets */
wire t_9250,   t_9251,   t_9252;
/* u2_3171 Output nets */
wire t_9253,   t_9254,   t_9255;
/* u2_3172 Output nets */
wire t_9256,   t_9257,   t_9258;
/* u2_3173 Output nets */
wire t_9259,   t_9260,   t_9261;
/* u2_3174 Output nets */
wire t_9262,   t_9263,   t_9264;
/* u2_3175 Output nets */
wire t_9265,   t_9266,   t_9267;
/* u2_3176 Output nets */
wire t_9268,   t_9269,   t_9270;
/* u2_3177 Output nets */
wire t_9271,   t_9272,   t_9273;
/* u2_3178 Output nets */
wire t_9274,   t_9275,   t_9276;
/* u2_3179 Output nets */
wire t_9277,   t_9278,   t_9279;
/* u1_3180 Output nets */
wire t_9280,   t_9281;
/* u2_3181 Output nets */
wire t_9282,   t_9283,   t_9284;
/* u2_3182 Output nets */
wire t_9285,   t_9286,   t_9287;
/* u2_3183 Output nets */
wire t_9288,   t_9289,   t_9290;
/* u0_3184 Output nets */
wire t_9291,   t_9292;
/* u2_3185 Output nets */
wire t_9293,   t_9294,   t_9295;
/* u2_3186 Output nets */
wire t_9296,   t_9297,   t_9298;
/* u2_3187 Output nets */
wire t_9299,   t_9300,   t_9301;
/* u0_3188 Output nets */
wire t_9302,   t_9303;
/* u2_3189 Output nets */
wire t_9304,   t_9305,   t_9306;
/* u2_3190 Output nets */
wire t_9307,   t_9308,   t_9309;
/* u2_3191 Output nets */
wire t_9310,   t_9311,   t_9312;
/* u1_3192 Output nets */
wire t_9313,   t_9314;
/* u2_3193 Output nets */
wire t_9315,   t_9316,   t_9317;
/* u2_3194 Output nets */
wire t_9318,   t_9319,   t_9320;
/* u2_3195 Output nets */
wire t_9321,   t_9322,   t_9323;
/* u0_3196 Output nets */
wire t_9324,   t_9325;
/* u2_3197 Output nets */
wire t_9326,   t_9327,   t_9328;
/* u2_3198 Output nets */
wire t_9329,   t_9330,   t_9331;
/* u2_3199 Output nets */
wire t_9332,   t_9333,   t_9334;
/* u0_3200 Output nets */
wire t_9335,   t_9336;
/* u2_3201 Output nets */
wire t_9337,   t_9338,   t_9339;
/* u2_3202 Output nets */
wire t_9340,   t_9341,   t_9342;
/* u2_3203 Output nets */
wire t_9343,   t_9344,   t_9345;
/* u0_3204 Output nets */
wire t_9346,   t_9347;
/* u2_3205 Output nets */
wire t_9348,   t_9349,   t_9350;
/* u2_3206 Output nets */
wire t_9351,   t_9352,   t_9353;
/* u2_3207 Output nets */
wire t_9354,   t_9355,   t_9356;
/* u0_3208 Output nets */
wire t_9357,   t_9358;
/* u2_3209 Output nets */
wire t_9359,   t_9360,   t_9361;
/* u2_3210 Output nets */
wire t_9362,   t_9363,   t_9364;
/* u2_3211 Output nets */
wire t_9365,   t_9366,   t_9367;
/* u2_3212 Output nets */
wire t_9368,   t_9369,   t_9370;
/* u2_3213 Output nets */
wire t_9371,   t_9372,   t_9373;
/* u2_3214 Output nets */
wire t_9374,   t_9375,   t_9376;
/* u2_3215 Output nets */
wire t_9377,   t_9378,   t_9379;
/* u2_3216 Output nets */
wire t_9380,   t_9381,   t_9382;
/* u2_3217 Output nets */
wire t_9383,   t_9384,   t_9385;
/* u2_3218 Output nets */
wire t_9386,   t_9387,   t_9388;
/* u2_3219 Output nets */
wire t_9389,   t_9390,   t_9391;
/* u2_3220 Output nets */
wire t_9392,   t_9393,   t_9394;
/* u2_3221 Output nets */
wire t_9395,   t_9396,   t_9397;
/* u2_3222 Output nets */
wire t_9398,   t_9399,   t_9400;
/* u2_3223 Output nets */
wire t_9401,   t_9402,   t_9403;
/* u2_3224 Output nets */
wire t_9404,   t_9405,   t_9406;
/* u2_3225 Output nets */
wire t_9407,   t_9408,   t_9409;
/* u2_3226 Output nets */
wire t_9410,   t_9411,   t_9412;
/* u2_3227 Output nets */
wire t_9413,   t_9414,   t_9415;
/* u2_3228 Output nets */
wire t_9416,   t_9417,   t_9418;
/* u2_3229 Output nets */
wire t_9419,   t_9420,   t_9421;
/* u2_3230 Output nets */
wire t_9422,   t_9423,   t_9424;
/* u2_3231 Output nets */
wire t_9425,   t_9426,   t_9427;
/* u2_3232 Output nets */
wire t_9428,   t_9429,   t_9430;
/* u2_3233 Output nets */
wire t_9431,   t_9432,   t_9433;
/* u2_3234 Output nets */
wire t_9434,   t_9435,   t_9436;
/* u1_3235 Output nets */
wire t_9437,   t_9438;
/* u2_3236 Output nets */
wire t_9439,   t_9440,   t_9441;
/* u2_3237 Output nets */
wire t_9442,   t_9443,   t_9444;
/* u0_3238 Output nets */
wire t_9445,   t_9446;
/* u2_3239 Output nets */
wire t_9447,   t_9448,   t_9449;
/* u2_3240 Output nets */
wire t_9450,   t_9451,   t_9452;
/* u0_3241 Output nets */
wire t_9453,   t_9454;
/* u2_3242 Output nets */
wire t_9455,   t_9456,   t_9457;
/* u2_3243 Output nets */
wire t_9458,   t_9459,   t_9460;
/* u1_3244 Output nets */
wire t_9461,   t_9462;
/* u2_3245 Output nets */
wire t_9463,   t_9464,   t_9465;
/* u2_3246 Output nets */
wire t_9466,   t_9467,   t_9468;
/* u0_3247 Output nets */
wire t_9469,   t_9470;
/* u2_3248 Output nets */
wire t_9471,   t_9472,   t_9473;
/* u2_3249 Output nets */
wire t_9474,   t_9475,   t_9476;
/* u0_3250 Output nets */
wire t_9477,   t_9478;
/* u2_3251 Output nets */
wire t_9479,   t_9480,   t_9481;
/* u2_3252 Output nets */
wire t_9482,   t_9483,   t_9484;
/* u0_3253 Output nets */
wire t_9485,   t_9486;
/* u2_3254 Output nets */
wire t_9487,   t_9488,   t_9489;
/* u2_3255 Output nets */
wire t_9490,   t_9491,   t_9492;
/* u0_3256 Output nets */
wire t_9493,   t_9494;
/* u2_3257 Output nets */
wire t_9495,   t_9496,   t_9497;
/* u2_3258 Output nets */
wire t_9498,   t_9499,   t_9500;
/* u2_3259 Output nets */
wire t_9501,   t_9502,   t_9503;
/* u2_3260 Output nets */
wire t_9504,   t_9505,   t_9506;
/* u2_3261 Output nets */
wire t_9507,   t_9508,   t_9509;
/* u2_3262 Output nets */
wire t_9510,   t_9511,   t_9512;
/* u2_3263 Output nets */
wire t_9513,   t_9514,   t_9515;
/* u2_3264 Output nets */
wire t_9516,   t_9517,   t_9518;
/* u2_3265 Output nets */
wire t_9519,   t_9520,   t_9521;
/* u2_3266 Output nets */
wire t_9522,   t_9523,   t_9524;
/* u2_3267 Output nets */
wire t_9525,   t_9526,   t_9527;
/* u2_3268 Output nets */
wire t_9528,   t_9529,   t_9530;
/* u2_3269 Output nets */
wire t_9531,   t_9532,   t_9533;
/* u2_3270 Output nets */
wire t_9534,   t_9535,   t_9536;
/* u2_3271 Output nets */
wire t_9537,   t_9538,   t_9539;
/* u2_3272 Output nets */
wire t_9540,   t_9541,   t_9542;
/* u2_3273 Output nets */
wire t_9543,   t_9544,   t_9545;
/* u1_3274 Output nets */
wire t_9546,   t_9547;
/* u2_3275 Output nets */
wire t_9548,   t_9549,   t_9550;
/* u0_3276 Output nets */
wire t_9551,   t_9552;
/* u2_3277 Output nets */
wire t_9553,   t_9554,   t_9555;
/* u0_3278 Output nets */
wire t_9556,   t_9557;
/* u2_3279 Output nets */
wire t_9558,   t_9559,   t_9560;
/* u1_3280 Output nets */
wire t_9561,   t_9562;
/* u2_3281 Output nets */
wire t_9563,   t_9564,   t_9565;
/* u0_3282 Output nets */
wire t_9566,   t_9567;
/* u2_3283 Output nets */
wire t_9568,   t_9569,   t_9570;
/* u0_3284 Output nets */
wire t_9571,   t_9572;
/* u2_3285 Output nets */
wire t_9573,   t_9574,   t_9575;
/* u0_3286 Output nets */
wire t_9576,   t_9577;
/* u2_3287 Output nets */
wire t_9578,   t_9579,   t_9580;
/* u0_3288 Output nets */
wire t_9581,   t_9582;
/* u2_3289 Output nets */
wire t_9583,   t_9584,   t_9585;
/* u2_3290 Output nets */
wire t_9586,   t_9587,   t_9588;
/* u2_3291 Output nets */
wire t_9589,   t_9590,   t_9591;
/* u2_3292 Output nets */
wire t_9592,   t_9593,   t_9594;
/* u2_3293 Output nets */
wire t_9595,   t_9596,   t_9597;
/* u2_3294 Output nets */
wire t_9598,   t_9599,   t_9600;
/* u2_3295 Output nets */
wire t_9601,   t_9602,   t_9603;
/* u2_3296 Output nets */
wire t_9604,   t_9605,   t_9606;
/* u1_3297 Output nets */
wire t_9607,   t_9608;
/* u0_3298 Output nets */
wire t_9609,   t_9610;
/* u0_3299 Output nets */
wire t_9611,   t_9612;
/* u1_3300 Output nets */
wire t_9613,   t_9614;
/* u0_3301 Output nets */
wire t_9615,   t_9616;
/* u0_3302 Output nets */
wire t_9617,   t_9618;
/* u0_3303 Output nets */
wire t_9619;

/* compress stage 2 */
half_adder u0_2161(.a(t_1), .b(s_1_0), .o(t_6335), .cout(t_6336));
half_adder u0_2162(.a(t_4), .b(t_3), .o(t_6337), .cout(t_6338));
compressor_3_2 u1_2163(.a(t_6), .b(t_5), .cin(s_4_3), .o(t_6339), .cout(t_6340));
half_adder u0_2164(.a(t_8), .b(t_7), .o(t_6341), .cout(t_6342));
half_adder u0_2165(.a(t_10), .b(t_9), .o(t_6343), .cout(t_6344));
half_adder u0_2166(.a(t_13), .b(t_11), .o(t_6345), .cout(t_6346));
compressor_3_2 u1_2167(.a(t_19), .b(t_16), .cin(t_14), .o(t_6347), .cout(t_6348));
compressor_3_2 u1_2168(.a(t_20), .b(t_17), .cin(s_9_4), .o(t_6349), .cout(t_6350));
compressor_3_2 u1_2169(.a(t_27), .b(t_24), .cin(t_22), .o(t_6351), .cout(t_6352));
compressor_3_2 u1_2170(.a(t_29), .b(t_28), .cin(t_25), .o(t_6353), .cout(t_6354));
compressor_4_2 u2_2171(.a(t_37), .b(t_34), .c(t_33), .d(t_30), .cin(s_12_7), .o(t_6355), .co(t_6356), .cout(t_6357));
compressor_4_2 u2_2172(.a(t_42), .b(t_39), .c(t_38), .d(t_35), .cin(t_6357), .o(t_6358), .co(t_6359), .cout(t_6360));
compressor_4_2 u2_2173(.a(t_47), .b(t_44), .c(t_43), .d(t_40), .cin(t_6360), .o(t_6361), .co(t_6362), .cout(t_6363));
compressor_4_2 u2_2174(.a(t_53), .b(t_50), .c(t_48), .d(t_45), .cin(t_6363), .o(t_6364), .co(t_6365), .cout(t_6366));
compressor_4_2 u2_2175(.a(t_59), .b(t_56), .c(t_54), .d(t_51), .cin(t_6366), .o(t_6367), .co(t_6368), .cout(t_6369));
compressor_4_2 u2_2176(.a(t_63), .b(t_60), .c(t_57), .d(s_17_8), .cin(t_6369), .o(t_6370), .co(t_6371), .cout(t_6372));
half_adder u0_2177(.a(t_67), .b(t_64), .o(t_6373), .cout(t_6374));
compressor_4_2 u2_2178(.a(t_73), .b(t_70), .c(t_68), .d(t_65), .cin(t_6372), .o(t_6375), .co(t_6376), .cout(t_6377));
compressor_4_2 u2_2179(.a(t_78), .b(t_77), .c(t_74), .d(t_71), .cin(t_6377), .o(t_6378), .co(t_6379), .cout(t_6380));
half_adder u0_2180(.a(t_84), .b(t_81), .o(t_6381), .cout(t_6382));
compressor_4_2 u2_2181(.a(t_85), .b(t_82), .c(t_79), .d(s_20_11), .cin(t_6380), .o(t_6383), .co(t_6384), .cout(t_6385));
compressor_3_2 u1_2182(.a(t_92), .b(t_89), .cin(t_86), .o(t_6386), .cout(t_6387));
compressor_4_2 u2_2183(.a(t_94), .b(t_93), .c(t_90), .d(t_87), .cin(t_6385), .o(t_6388), .co(t_6389), .cout(t_6390));
half_adder u0_2184(.a(t_100), .b(t_97), .o(t_6391), .cout(t_6392));
compressor_4_2 u2_2185(.a(t_102), .b(t_101), .c(t_98), .d(t_95), .cin(t_6390), .o(t_6393), .co(t_6394), .cout(t_6395));
half_adder u0_2186(.a(t_108), .b(t_105), .o(t_6396), .cout(t_6397));
compressor_4_2 u2_2187(.a(t_111), .b(t_109), .c(t_106), .d(t_103), .cin(t_6395), .o(t_6398), .co(t_6399), .cout(t_6400));
half_adder u0_2188(.a(t_117), .b(t_114), .o(t_6401), .cout(t_6402));
compressor_4_2 u2_2189(.a(t_120), .b(t_118), .c(t_115), .d(t_112), .cin(t_6400), .o(t_6403), .co(t_6404), .cout(t_6405));
compressor_3_2 u1_2190(.a(t_129), .b(t_126), .cin(t_123), .o(t_6406), .cout(t_6407));
compressor_4_2 u2_2191(.a(t_127), .b(t_124), .c(t_121), .d(s_25_12), .cin(t_6405), .o(t_6408), .co(t_6409), .cout(t_6410));
compressor_3_2 u1_2192(.a(t_134), .b(t_131), .cin(t_130), .o(t_6411), .cout(t_6412));
compressor_4_2 u2_2193(.a(t_140), .b(t_138), .c(t_135), .d(t_132), .cin(t_6410), .o(t_6413), .co(t_6414), .cout(t_6415));
compressor_3_2 u1_2194(.a(t_149), .b(t_146), .cin(t_143), .o(t_6416), .cout(t_6417));
compressor_4_2 u2_2195(.a(t_150), .b(t_147), .c(t_144), .d(t_141), .cin(t_6415), .o(t_6418), .co(t_6419), .cout(t_6420));
compressor_3_2 u1_2196(.a(t_157), .b(t_154), .cin(t_151), .o(t_6421), .cout(t_6422));
compressor_4_2 u2_2197(.a(t_158), .b(t_155), .c(t_152), .d(s_28_15), .cin(t_6420), .o(t_6423), .co(t_6424), .cout(t_6425));
compressor_4_2 u2_2198(.a(t_171), .b(t_168), .c(t_165), .d(t_162), .cin(t_161), .o(t_6426), .co(t_6427), .cout(t_6428));
compressor_4_2 u2_2199(.a(t_172), .b(t_169), .c(t_166), .d(t_163), .cin(t_6425), .o(t_6429), .co(t_6430), .cout(t_6431));
compressor_4_2 u2_2200(.a(t_182), .b(t_179), .c(t_176), .d(t_173), .cin(t_6428), .o(t_6432), .co(t_6433), .cout(t_6434));
compressor_4_2 u2_2201(.a(t_183), .b(t_180), .c(t_177), .d(t_174), .cin(t_6431), .o(t_6435), .co(t_6436), .cout(t_6437));
compressor_4_2 u2_2202(.a(t_193), .b(t_190), .c(t_187), .d(t_184), .cin(t_6434), .o(t_6438), .co(t_6439), .cout(t_6440));
compressor_4_2 u2_2203(.a(t_194), .b(t_191), .c(t_188), .d(t_185), .cin(t_6437), .o(t_6441), .co(t_6442), .cout(t_6443));
compressor_4_2 u2_2204(.a(t_205), .b(t_202), .c(t_199), .d(t_196), .cin(t_6440), .o(t_6444), .co(t_6445), .cout(t_6446));
compressor_4_2 u2_2205(.a(t_206), .b(t_203), .c(t_200), .d(t_197), .cin(t_6443), .o(t_6447), .co(t_6448), .cout(t_6449));
compressor_4_2 u2_2206(.a(t_217), .b(t_214), .c(t_211), .d(t_208), .cin(t_6446), .o(t_6450), .co(t_6451), .cout(t_6452));
compressor_4_2 u2_2207(.a(t_215), .b(t_212), .c(t_209), .d(s_33_16), .cin(t_6449), .o(t_6453), .co(t_6454), .cout(t_6455));
compressor_4_2 u2_2208(.a(t_225), .b(t_222), .c(t_221), .d(t_218), .cin(t_6452), .o(t_6456), .co(t_6457), .cout(t_6458));
half_adder u0_2209(.a(t_231), .b(t_228), .o(t_6459), .cout(t_6460));
compressor_4_2 u2_2210(.a(t_232), .b(t_229), .c(t_226), .d(t_223), .cin(t_6455), .o(t_6461), .co(t_6462), .cout(t_6463));
compressor_4_2 u2_2211(.a(t_243), .b(t_240), .c(t_237), .d(t_234), .cin(t_6458), .o(t_6464), .co(t_6465), .cout(t_6466));
compressor_4_2 u2_2212(.a(t_244), .b(t_241), .c(t_238), .d(t_235), .cin(t_6463), .o(t_6467), .co(t_6468), .cout(t_6469));
compressor_4_2 u2_2213(.a(t_254), .b(t_251), .c(t_248), .d(t_247), .cin(t_6466), .o(t_6470), .co(t_6471), .cout(t_6472));
half_adder u0_2214(.a(t_260), .b(t_257), .o(t_6473), .cout(t_6474));
compressor_4_2 u2_2215(.a(t_255), .b(t_252), .c(t_249), .d(s_36_19), .cin(t_6469), .o(t_6475), .co(t_6476), .cout(t_6477));
compressor_4_2 u2_2216(.a(t_265), .b(t_262), .c(t_261), .d(t_258), .cin(t_6472), .o(t_6478), .co(t_6479), .cout(t_6480));
compressor_3_2 u1_2217(.a(t_274), .b(t_271), .cin(t_268), .o(t_6481), .cout(t_6482));
compressor_4_2 u2_2218(.a(t_272), .b(t_269), .c(t_266), .d(t_263), .cin(t_6477), .o(t_6483), .co(t_6484), .cout(t_6485));
compressor_4_2 u2_2219(.a(t_282), .b(t_279), .c(t_276), .d(t_275), .cin(t_6480), .o(t_6486), .co(t_6487), .cout(t_6488));
half_adder u0_2220(.a(t_288), .b(t_285), .o(t_6489), .cout(t_6490));
compressor_4_2 u2_2221(.a(t_286), .b(t_283), .c(t_280), .d(t_277), .cin(t_6485), .o(t_6491), .co(t_6492), .cout(t_6493));
compressor_4_2 u2_2222(.a(t_296), .b(t_293), .c(t_290), .d(t_289), .cin(t_6488), .o(t_6494), .co(t_6495), .cout(t_6496));
half_adder u0_2223(.a(t_302), .b(t_299), .o(t_6497), .cout(t_6498));
compressor_4_2 u2_2224(.a(t_300), .b(t_297), .c(t_294), .d(t_291), .cin(t_6493), .o(t_6499), .co(t_6500), .cout(t_6501));
compressor_4_2 u2_2225(.a(t_311), .b(t_308), .c(t_305), .d(t_303), .cin(t_6496), .o(t_6502), .co(t_6503), .cout(t_6504));
half_adder u0_2226(.a(t_317), .b(t_314), .o(t_6505), .cout(t_6506));
compressor_4_2 u2_2227(.a(t_315), .b(t_312), .c(t_309), .d(t_306), .cin(t_6501), .o(t_6507), .co(t_6508), .cout(t_6509));
compressor_4_2 u2_2228(.a(t_326), .b(t_323), .c(t_320), .d(t_318), .cin(t_6504), .o(t_6510), .co(t_6511), .cout(t_6512));
compressor_3_2 u1_2229(.a(t_335), .b(t_332), .cin(t_329), .o(t_6513), .cout(t_6514));
compressor_4_2 u2_2230(.a(t_327), .b(t_324), .c(t_321), .d(s_41_20), .cin(t_6509), .o(t_6515), .co(t_6516), .cout(t_6517));
compressor_4_2 u2_2231(.a(t_337), .b(t_336), .c(t_333), .d(t_330), .cin(t_6512), .o(t_6518), .co(t_6519), .cout(t_6520));
compressor_3_2 u1_2232(.a(t_346), .b(t_343), .cin(t_340), .o(t_6521), .cout(t_6522));
compressor_4_2 u2_2233(.a(t_347), .b(t_344), .c(t_341), .d(t_338), .cin(t_6517), .o(t_6523), .co(t_6524), .cout(t_6525));
compressor_4_2 u2_2234(.a(t_358), .b(t_355), .c(t_352), .d(t_350), .cin(t_6520), .o(t_6526), .co(t_6527), .cout(t_6528));
compressor_3_2 u1_2235(.a(t_367), .b(t_364), .cin(t_361), .o(t_6529), .cout(t_6530));
compressor_4_2 u2_2236(.a(t_362), .b(t_359), .c(t_356), .d(t_353), .cin(t_6525), .o(t_6531), .co(t_6532), .cout(t_6533));
compressor_4_2 u2_2237(.a(t_372), .b(t_369), .c(t_368), .d(t_365), .cin(t_6528), .o(t_6534), .co(t_6535), .cout(t_6536));
compressor_3_2 u1_2238(.a(t_381), .b(t_378), .cin(t_375), .o(t_6537), .cout(t_6538));
compressor_4_2 u2_2239(.a(t_376), .b(t_373), .c(t_370), .d(s_44_23), .cin(t_6533), .o(t_6539), .co(t_6540), .cout(t_6541));
compressor_4_2 u2_2240(.a(t_386), .b(t_385), .c(t_382), .d(t_379), .cin(t_6536), .o(t_6542), .co(t_6543), .cout(t_6544));
compressor_4_2 u2_2241(.a(t_401), .b(t_398), .c(t_395), .d(t_392), .cin(t_389), .o(t_6545), .co(t_6546), .cout(t_6547));
compressor_4_2 u2_2242(.a(t_396), .b(t_393), .c(t_390), .d(t_387), .cin(t_6541), .o(t_6548), .co(t_6549), .cout(t_6550));
compressor_4_2 u2_2243(.a(t_406), .b(t_403), .c(t_402), .d(t_399), .cin(t_6544), .o(t_6551), .co(t_6552), .cout(t_6553));
compressor_4_2 u2_2244(.a(t_418), .b(t_415), .c(t_412), .d(t_409), .cin(t_6547), .o(t_6554), .co(t_6555), .cout(t_6556));
compressor_4_2 u2_2245(.a(t_413), .b(t_410), .c(t_407), .d(t_404), .cin(t_6550), .o(t_6557), .co(t_6558), .cout(t_6559));
compressor_4_2 u2_2246(.a(t_423), .b(t_420), .c(t_419), .d(t_416), .cin(t_6553), .o(t_6560), .co(t_6561), .cout(t_6562));
compressor_4_2 u2_2247(.a(t_435), .b(t_432), .c(t_429), .d(t_426), .cin(t_6556), .o(t_6563), .co(t_6564), .cout(t_6565));
compressor_4_2 u2_2248(.a(t_430), .b(t_427), .c(t_424), .d(t_421), .cin(t_6559), .o(t_6566), .co(t_6567), .cout(t_6568));
compressor_4_2 u2_2249(.a(t_441), .b(t_438), .c(t_436), .d(t_433), .cin(t_6562), .o(t_6569), .co(t_6570), .cout(t_6571));
compressor_4_2 u2_2250(.a(t_453), .b(t_450), .c(t_447), .d(t_444), .cin(t_6565), .o(t_6572), .co(t_6573), .cout(t_6574));
compressor_4_2 u2_2251(.a(t_448), .b(t_445), .c(t_442), .d(t_439), .cin(t_6568), .o(t_6575), .co(t_6576), .cout(t_6577));
compressor_4_2 u2_2252(.a(t_459), .b(t_456), .c(t_454), .d(t_451), .cin(t_6571), .o(t_6578), .co(t_6579), .cout(t_6580));
compressor_4_2 u2_2253(.a(t_471), .b(t_468), .c(t_465), .d(t_462), .cin(t_6574), .o(t_6581), .co(t_6582), .cout(t_6583));
compressor_4_2 u2_2254(.a(t_463), .b(t_460), .c(t_457), .d(s_49_24), .cin(t_6577), .o(t_6584), .co(t_6585), .cout(t_6586));
compressor_4_2 u2_2255(.a(t_475), .b(t_472), .c(t_469), .d(t_466), .cin(t_6580), .o(t_6587), .co(t_6588), .cout(t_6589));
compressor_4_2 u2_2256(.a(t_485), .b(t_482), .c(t_479), .d(t_476), .cin(t_6583), .o(t_6590), .co(t_6591), .cout(t_6592));
half_adder u0_2257(.a(t_491), .b(t_488), .o(t_6593), .cout(t_6594));
compressor_4_2 u2_2258(.a(t_486), .b(t_483), .c(t_480), .d(t_477), .cin(t_6586), .o(t_6595), .co(t_6596), .cout(t_6597));
compressor_4_2 u2_2259(.a(t_497), .b(t_494), .c(t_492), .d(t_489), .cin(t_6589), .o(t_6598), .co(t_6599), .cout(t_6600));
compressor_4_2 u2_2260(.a(t_509), .b(t_506), .c(t_503), .d(t_500), .cin(t_6592), .o(t_6601), .co(t_6602), .cout(t_6603));
compressor_4_2 u2_2261(.a(t_504), .b(t_501), .c(t_498), .d(t_495), .cin(t_6597), .o(t_6604), .co(t_6605), .cout(t_6606));
compressor_4_2 u2_2262(.a(t_514), .b(t_513), .c(t_510), .d(t_507), .cin(t_6600), .o(t_6607), .co(t_6608), .cout(t_6609));
compressor_4_2 u2_2263(.a(t_526), .b(t_523), .c(t_520), .d(t_517), .cin(t_6603), .o(t_6610), .co(t_6611), .cout(t_6612));
half_adder u0_2264(.a(t_532), .b(t_529), .o(t_6613), .cout(t_6614));
compressor_4_2 u2_2265(.a(t_521), .b(t_518), .c(t_515), .d(s_52_27), .cin(t_6606), .o(t_6615), .co(t_6616), .cout(t_6617));
compressor_4_2 u2_2266(.a(t_533), .b(t_530), .c(t_527), .d(t_524), .cin(t_6609), .o(t_6618), .co(t_6619), .cout(t_6620));
compressor_4_2 u2_2267(.a(t_543), .b(t_540), .c(t_537), .d(t_534), .cin(t_6612), .o(t_6621), .co(t_6622), .cout(t_6623));
compressor_3_2 u1_2268(.a(t_552), .b(t_549), .cin(t_546), .o(t_6624), .cout(t_6625));
compressor_4_2 u2_2269(.a(t_544), .b(t_541), .c(t_538), .d(t_535), .cin(t_6617), .o(t_6626), .co(t_6627), .cout(t_6628));
compressor_4_2 u2_2270(.a(t_554), .b(t_553), .c(t_550), .d(t_547), .cin(t_6620), .o(t_6629), .co(t_6630), .cout(t_6631));
compressor_4_2 u2_2271(.a(t_566), .b(t_563), .c(t_560), .d(t_557), .cin(t_6623), .o(t_6632), .co(t_6633), .cout(t_6634));
half_adder u0_2272(.a(t_572), .b(t_569), .o(t_6635), .cout(t_6636));
compressor_4_2 u2_2273(.a(t_564), .b(t_561), .c(t_558), .d(t_555), .cin(t_6628), .o(t_6637), .co(t_6638), .cout(t_6639));
compressor_4_2 u2_2274(.a(t_574), .b(t_573), .c(t_570), .d(t_567), .cin(t_6631), .o(t_6640), .co(t_6641), .cout(t_6642));
compressor_4_2 u2_2275(.a(t_586), .b(t_583), .c(t_580), .d(t_577), .cin(t_6634), .o(t_6643), .co(t_6644), .cout(t_6645));
half_adder u0_2276(.a(t_592), .b(t_589), .o(t_6646), .cout(t_6647));
compressor_4_2 u2_2277(.a(t_584), .b(t_581), .c(t_578), .d(t_575), .cin(t_6639), .o(t_6648), .co(t_6649), .cout(t_6650));
compressor_4_2 u2_2278(.a(t_595), .b(t_593), .c(t_590), .d(t_587), .cin(t_6642), .o(t_6651), .co(t_6652), .cout(t_6653));
compressor_4_2 u2_2279(.a(t_607), .b(t_604), .c(t_601), .d(t_598), .cin(t_6645), .o(t_6654), .co(t_6655), .cout(t_6656));
half_adder u0_2280(.a(t_613), .b(t_610), .o(t_6657), .cout(t_6658));
compressor_4_2 u2_2281(.a(t_605), .b(t_602), .c(t_599), .d(t_596), .cin(t_6650), .o(t_6659), .co(t_6660), .cout(t_6661));
compressor_4_2 u2_2282(.a(t_616), .b(t_614), .c(t_611), .d(t_608), .cin(t_6653), .o(t_6662), .co(t_6663), .cout(t_6664));
compressor_4_2 u2_2283(.a(t_628), .b(t_625), .c(t_622), .d(t_619), .cin(t_6656), .o(t_6665), .co(t_6666), .cout(t_6667));
compressor_3_2 u1_2284(.a(t_637), .b(t_634), .cin(t_631), .o(t_6668), .cout(t_6669));
compressor_4_2 u2_2285(.a(t_623), .b(t_620), .c(t_617), .d(s_57_28), .cin(t_6661), .o(t_6670), .co(t_6671), .cout(t_6672));
compressor_4_2 u2_2286(.a(t_635), .b(t_632), .c(t_629), .d(t_626), .cin(t_6664), .o(t_6673), .co(t_6674), .cout(t_6675));
compressor_4_2 u2_2287(.a(t_645), .b(t_642), .c(t_639), .d(t_638), .cin(t_6667), .o(t_6676), .co(t_6677), .cout(t_6678));
compressor_3_2 u1_2288(.a(t_654), .b(t_651), .cin(t_648), .o(t_6679), .cout(t_6680));
compressor_4_2 u2_2289(.a(t_649), .b(t_646), .c(t_643), .d(t_640), .cin(t_6672), .o(t_6681), .co(t_6682), .cout(t_6683));
compressor_4_2 u2_2290(.a(t_660), .b(t_658), .c(t_655), .d(t_652), .cin(t_6675), .o(t_6684), .co(t_6685), .cout(t_6686));
compressor_4_2 u2_2291(.a(t_672), .b(t_669), .c(t_666), .d(t_663), .cin(t_6678), .o(t_6687), .co(t_6688), .cout(t_6689));
compressor_3_2 u1_2292(.a(t_681), .b(t_678), .cin(t_675), .o(t_6690), .cout(t_6691));
compressor_4_2 u2_2293(.a(t_670), .b(t_667), .c(t_664), .d(t_661), .cin(t_6683), .o(t_6692), .co(t_6693), .cout(t_6694));
compressor_4_2 u2_2294(.a(t_682), .b(t_679), .c(t_676), .d(t_673), .cin(t_6686), .o(t_6695), .co(t_6696), .cout(t_6697));
compressor_4_2 u2_2295(.a(t_692), .b(t_689), .c(t_686), .d(t_683), .cin(t_6689), .o(t_6698), .co(t_6699), .cout(t_6700));
compressor_3_2 u1_2296(.a(t_701), .b(t_698), .cin(t_695), .o(t_6701), .cout(t_6702));
compressor_4_2 u2_2297(.a(t_690), .b(t_687), .c(t_684), .d(s_60_31), .cin(t_6694), .o(t_6703), .co(t_6704), .cout(t_6705));
compressor_4_2 u2_2298(.a(t_702), .b(t_699), .c(t_696), .d(t_693), .cin(t_6697), .o(t_6706), .co(t_6707), .cout(t_6708));
compressor_4_2 u2_2299(.a(t_712), .b(t_709), .c(t_706), .d(t_705), .cin(t_6700), .o(t_6709), .co(t_6710), .cout(t_6711));
compressor_4_2 u2_2300(.a(t_727), .b(t_724), .c(t_721), .d(t_718), .cin(t_715), .o(t_6712), .co(t_6713), .cout(t_6714));
compressor_4_2 u2_2301(.a(t_716), .b(t_713), .c(t_710), .d(t_707), .cin(t_6705), .o(t_6715), .co(t_6716), .cout(t_6717));
compressor_4_2 u2_2302(.a(t_728), .b(t_725), .c(t_722), .d(t_719), .cin(t_6708), .o(t_6718), .co(t_6719), .cout(t_6720));
compressor_4_2 u2_2303(.a(t_738), .b(t_735), .c(t_732), .d(t_729), .cin(t_6711), .o(t_6721), .co(t_6722), .cout(t_6723));
compressor_4_2 u2_2304(.a(t_750), .b(t_747), .c(t_744), .d(t_741), .cin(t_6714), .o(t_6724), .co(t_6725), .cout(t_6726));
compressor_4_2 u2_2305(.a(t_739), .b(t_736), .c(t_733), .d(t_730), .cin(t_6717), .o(t_6727), .co(t_6728), .cout(t_6729));
compressor_4_2 u2_2306(.a(t_751), .b(t_748), .c(t_745), .d(t_742), .cin(t_6720), .o(t_6730), .co(t_6731), .cout(t_6732));
compressor_4_2 u2_2307(.a(t_761), .b(t_758), .c(t_755), .d(t_752), .cin(t_6723), .o(t_6733), .co(t_6734), .cout(t_6735));
compressor_4_2 u2_2308(.a(t_773), .b(t_770), .c(t_767), .d(t_764), .cin(t_6726), .o(t_6736), .co(t_6737), .cout(t_6738));
compressor_4_2 u2_2309(.a(t_762), .b(t_759), .c(t_756), .d(t_753), .cin(t_6729), .o(t_6739), .co(t_6740), .cout(t_6741));
compressor_4_2 u2_2310(.a(t_774), .b(t_771), .c(t_768), .d(t_765), .cin(t_6732), .o(t_6742), .co(t_6743), .cout(t_6744));
compressor_4_2 u2_2311(.a(t_785), .b(t_782), .c(t_779), .d(t_776), .cin(t_6735), .o(t_6745), .co(t_6746), .cout(t_6747));
compressor_4_2 u2_2312(.a(t_797), .b(t_794), .c(t_791), .d(t_788), .cin(t_6738), .o(t_6748), .co(t_6749), .cout(t_6750));
compressor_4_2 u2_2313(.a(t_786), .b(t_783), .c(t_780), .d(t_777), .cin(t_6741), .o(t_6751), .co(t_6752), .cout(t_6753));
compressor_4_2 u2_2314(.a(t_798), .b(t_795), .c(t_792), .d(t_789), .cin(t_6744), .o(t_6754), .co(t_6755), .cout(t_6756));
compressor_4_2 u2_2315(.a(t_809), .b(t_806), .c(t_803), .d(t_800), .cin(t_6747), .o(t_6757), .co(t_6758), .cout(t_6759));
compressor_4_2 u2_2316(.a(t_821), .b(t_818), .c(t_815), .d(t_812), .cin(t_6750), .o(t_6760), .co(t_6761), .cout(t_6762));
compressor_4_2 u2_2317(.a(t_807), .b(t_804), .c(t_801), .d(s_65_32), .cin(t_6753), .o(t_6763), .co(t_6764), .cout(t_6765));
compressor_4_2 u2_2318(.a(t_819), .b(t_816), .c(t_813), .d(t_810), .cin(t_6756), .o(t_6766), .co(t_6767), .cout(t_6768));
compressor_4_2 u2_2319(.a(t_829), .b(t_826), .c(t_825), .d(t_822), .cin(t_6759), .o(t_6769), .co(t_6770), .cout(t_6771));
compressor_4_2 u2_2320(.a(t_841), .b(t_838), .c(t_835), .d(t_832), .cin(t_6762), .o(t_6772), .co(t_6773), .cout(t_6774));
half_adder u0_2321(.a(t_847), .b(t_844), .o(t_6775), .cout(t_6776));
compressor_4_2 u2_2322(.a(t_836), .b(t_833), .c(t_830), .d(t_827), .cin(t_6765), .o(t_6777), .co(t_6778), .cout(t_6779));
compressor_4_2 u2_2323(.a(t_848), .b(t_845), .c(t_842), .d(t_839), .cin(t_6768), .o(t_6780), .co(t_6781), .cout(t_6782));
compressor_4_2 u2_2324(.a(t_859), .b(t_856), .c(t_853), .d(t_850), .cin(t_6771), .o(t_6783), .co(t_6784), .cout(t_6785));
compressor_4_2 u2_2325(.a(t_871), .b(t_868), .c(t_865), .d(t_862), .cin(t_6774), .o(t_6786), .co(t_6787), .cout(t_6788));
compressor_4_2 u2_2326(.a(t_860), .b(t_857), .c(t_854), .d(t_851), .cin(t_6779), .o(t_6789), .co(t_6790), .cout(t_6791));
compressor_4_2 u2_2327(.a(t_872), .b(t_869), .c(t_866), .d(t_863), .cin(t_6782), .o(t_6792), .co(t_6793), .cout(t_6794));
compressor_4_2 u2_2328(.a(t_882), .b(t_879), .c(t_876), .d(t_875), .cin(t_6785), .o(t_6795), .co(t_6796), .cout(t_6797));
compressor_4_2 u2_2329(.a(t_894), .b(t_891), .c(t_888), .d(t_885), .cin(t_6788), .o(t_6798), .co(t_6799), .cout(t_6800));
half_adder u0_2330(.a(t_900), .b(t_897), .o(t_6801), .cout(t_6802));
compressor_4_2 u2_2331(.a(t_883), .b(t_880), .c(t_877), .d(s_68_35), .cin(t_6791), .o(t_6803), .co(t_6804), .cout(t_6805));
compressor_4_2 u2_2332(.a(t_895), .b(t_892), .c(t_889), .d(t_886), .cin(t_6794), .o(t_6806), .co(t_6807), .cout(t_6808));
compressor_4_2 u2_2333(.a(t_905), .b(t_902), .c(t_901), .d(t_898), .cin(t_6797), .o(t_6809), .co(t_6810), .cout(t_6811));
compressor_4_2 u2_2334(.a(t_917), .b(t_914), .c(t_911), .d(t_908), .cin(t_6800), .o(t_6812), .co(t_6813), .cout(t_6814));
compressor_3_2 u1_2335(.a(t_926), .b(t_923), .cin(t_920), .o(t_6815), .cout(t_6816));
compressor_4_2 u2_2336(.a(t_912), .b(t_909), .c(t_906), .d(t_903), .cin(t_6805), .o(t_6817), .co(t_6818), .cout(t_6819));
compressor_4_2 u2_2337(.a(t_924), .b(t_921), .c(t_918), .d(t_915), .cin(t_6808), .o(t_6820), .co(t_6821), .cout(t_6822));
compressor_4_2 u2_2338(.a(t_934), .b(t_931), .c(t_928), .d(t_927), .cin(t_6811), .o(t_6823), .co(t_6824), .cout(t_6825));
compressor_4_2 u2_2339(.a(t_946), .b(t_943), .c(t_940), .d(t_937), .cin(t_6814), .o(t_6826), .co(t_6827), .cout(t_6828));
half_adder u0_2340(.a(t_952), .b(t_949), .o(t_6829), .cout(t_6830));
compressor_4_2 u2_2341(.a(t_938), .b(t_935), .c(t_932), .d(t_929), .cin(t_6819), .o(t_6831), .co(t_6832), .cout(t_6833));
compressor_4_2 u2_2342(.a(t_950), .b(t_947), .c(t_944), .d(t_941), .cin(t_6822), .o(t_6834), .co(t_6835), .cout(t_6836));
compressor_4_2 u2_2343(.a(t_960), .b(t_957), .c(t_954), .d(t_953), .cin(t_6825), .o(t_6837), .co(t_6838), .cout(t_6839));
compressor_4_2 u2_2344(.a(t_972), .b(t_969), .c(t_966), .d(t_963), .cin(t_6828), .o(t_6840), .co(t_6841), .cout(t_6842));
half_adder u0_2345(.a(t_978), .b(t_975), .o(t_6843), .cout(t_6844));
compressor_4_2 u2_2346(.a(t_964), .b(t_961), .c(t_958), .d(t_955), .cin(t_6833), .o(t_6845), .co(t_6846), .cout(t_6847));
compressor_4_2 u2_2347(.a(t_976), .b(t_973), .c(t_970), .d(t_967), .cin(t_6836), .o(t_6848), .co(t_6849), .cout(t_6850));
compressor_4_2 u2_2348(.a(t_987), .b(t_984), .c(t_981), .d(t_979), .cin(t_6839), .o(t_6851), .co(t_6852), .cout(t_6853));
compressor_4_2 u2_2349(.a(t_999), .b(t_996), .c(t_993), .d(t_990), .cin(t_6842), .o(t_6854), .co(t_6855), .cout(t_6856));
half_adder u0_2350(.a(t_1005), .b(t_1002), .o(t_6857), .cout(t_6858));
compressor_4_2 u2_2351(.a(t_991), .b(t_988), .c(t_985), .d(t_982), .cin(t_6847), .o(t_6859), .co(t_6860), .cout(t_6861));
compressor_4_2 u2_2352(.a(t_1003), .b(t_1000), .c(t_997), .d(t_994), .cin(t_6850), .o(t_6862), .co(t_6863), .cout(t_6864));
compressor_4_2 u2_2353(.a(t_1014), .b(t_1011), .c(t_1008), .d(t_1006), .cin(t_6853), .o(t_6865), .co(t_6866), .cout(t_6867));
compressor_4_2 u2_2354(.a(t_1026), .b(t_1023), .c(t_1020), .d(t_1017), .cin(t_6856), .o(t_6868), .co(t_6869), .cout(t_6870));
compressor_3_2 u1_2355(.a(t_1035), .b(t_1032), .cin(t_1029), .o(t_6871), .cout(t_6872));
compressor_4_2 u2_2356(.a(t_1015), .b(t_1012), .c(t_1009), .d(s_73_36), .cin(t_6861), .o(t_6873), .co(t_6874), .cout(t_6875));
compressor_4_2 u2_2357(.a(t_1027), .b(t_1024), .c(t_1021), .d(t_1018), .cin(t_6864), .o(t_6876), .co(t_6877), .cout(t_6878));
compressor_4_2 u2_2358(.a(t_1037), .b(t_1036), .c(t_1033), .d(t_1030), .cin(t_6867), .o(t_6879), .co(t_6880), .cout(t_6881));
compressor_4_2 u2_2359(.a(t_1049), .b(t_1046), .c(t_1043), .d(t_1040), .cin(t_6870), .o(t_6882), .co(t_6883), .cout(t_6884));
compressor_3_2 u1_2360(.a(t_1058), .b(t_1055), .cin(t_1052), .o(t_6885), .cout(t_6886));
compressor_4_2 u2_2361(.a(t_1047), .b(t_1044), .c(t_1041), .d(t_1038), .cin(t_6875), .o(t_6887), .co(t_6888), .cout(t_6889));
compressor_4_2 u2_2362(.a(t_1059), .b(t_1056), .c(t_1053), .d(t_1050), .cin(t_6878), .o(t_6890), .co(t_6891), .cout(t_6892));
compressor_4_2 u2_2363(.a(t_1070), .b(t_1067), .c(t_1064), .d(t_1062), .cin(t_6881), .o(t_6893), .co(t_6894), .cout(t_6895));
compressor_4_2 u2_2364(.a(t_1082), .b(t_1079), .c(t_1076), .d(t_1073), .cin(t_6884), .o(t_6896), .co(t_6897), .cout(t_6898));
compressor_3_2 u1_2365(.a(t_1091), .b(t_1088), .cin(t_1085), .o(t_6899), .cout(t_6900));
compressor_4_2 u2_2366(.a(t_1074), .b(t_1071), .c(t_1068), .d(t_1065), .cin(t_6889), .o(t_6901), .co(t_6902), .cout(t_6903));
compressor_4_2 u2_2367(.a(t_1086), .b(t_1083), .c(t_1080), .d(t_1077), .cin(t_6892), .o(t_6904), .co(t_6905), .cout(t_6906));
compressor_4_2 u2_2368(.a(t_1096), .b(t_1093), .c(t_1092), .d(t_1089), .cin(t_6895), .o(t_6907), .co(t_6908), .cout(t_6909));
compressor_4_2 u2_2369(.a(t_1108), .b(t_1105), .c(t_1102), .d(t_1099), .cin(t_6898), .o(t_6910), .co(t_6911), .cout(t_6912));
compressor_3_2 u1_2370(.a(t_1117), .b(t_1114), .cin(t_1111), .o(t_6913), .cout(t_6914));
compressor_4_2 u2_2371(.a(t_1100), .b(t_1097), .c(t_1094), .d(s_76_39), .cin(t_6903), .o(t_6915), .co(t_6916), .cout(t_6917));
compressor_4_2 u2_2372(.a(t_1112), .b(t_1109), .c(t_1106), .d(t_1103), .cin(t_6906), .o(t_6918), .co(t_6919), .cout(t_6920));
compressor_4_2 u2_2373(.a(t_1122), .b(t_1121), .c(t_1118), .d(t_1115), .cin(t_6909), .o(t_6921), .co(t_6922), .cout(t_6923));
compressor_4_2 u2_2374(.a(t_1134), .b(t_1131), .c(t_1128), .d(t_1125), .cin(t_6912), .o(t_6924), .co(t_6925), .cout(t_6926));
compressor_4_2 u2_2375(.a(t_1149), .b(t_1146), .c(t_1143), .d(t_1140), .cin(t_1137), .o(t_6927), .co(t_6928), .cout(t_6929));
compressor_4_2 u2_2376(.a(t_1132), .b(t_1129), .c(t_1126), .d(t_1123), .cin(t_6917), .o(t_6930), .co(t_6931), .cout(t_6932));
compressor_4_2 u2_2377(.a(t_1144), .b(t_1141), .c(t_1138), .d(t_1135), .cin(t_6920), .o(t_6933), .co(t_6934), .cout(t_6935));
compressor_4_2 u2_2378(.a(t_1154), .b(t_1151), .c(t_1150), .d(t_1147), .cin(t_6923), .o(t_6936), .co(t_6937), .cout(t_6938));
compressor_4_2 u2_2379(.a(t_1166), .b(t_1163), .c(t_1160), .d(t_1157), .cin(t_6926), .o(t_6939), .co(t_6940), .cout(t_6941));
compressor_4_2 u2_2380(.a(t_1178), .b(t_1175), .c(t_1172), .d(t_1169), .cin(t_6929), .o(t_6942), .co(t_6943), .cout(t_6944));
compressor_4_2 u2_2381(.a(t_1161), .b(t_1158), .c(t_1155), .d(t_1152), .cin(t_6932), .o(t_6945), .co(t_6946), .cout(t_6947));
compressor_4_2 u2_2382(.a(t_1173), .b(t_1170), .c(t_1167), .d(t_1164), .cin(t_6935), .o(t_6948), .co(t_6949), .cout(t_6950));
compressor_4_2 u2_2383(.a(t_1183), .b(t_1180), .c(t_1179), .d(t_1176), .cin(t_6938), .o(t_6951), .co(t_6952), .cout(t_6953));
compressor_4_2 u2_2384(.a(t_1195), .b(t_1192), .c(t_1189), .d(t_1186), .cin(t_6941), .o(t_6954), .co(t_6955), .cout(t_6956));
compressor_4_2 u2_2385(.a(t_1207), .b(t_1204), .c(t_1201), .d(t_1198), .cin(t_6944), .o(t_6957), .co(t_6958), .cout(t_6959));
compressor_4_2 u2_2386(.a(t_1190), .b(t_1187), .c(t_1184), .d(t_1181), .cin(t_6947), .o(t_6960), .co(t_6961), .cout(t_6962));
compressor_4_2 u2_2387(.a(t_1202), .b(t_1199), .c(t_1196), .d(t_1193), .cin(t_6950), .o(t_6963), .co(t_6964), .cout(t_6965));
compressor_4_2 u2_2388(.a(t_1213), .b(t_1210), .c(t_1208), .d(t_1205), .cin(t_6953), .o(t_6966), .co(t_6967), .cout(t_6968));
compressor_4_2 u2_2389(.a(t_1225), .b(t_1222), .c(t_1219), .d(t_1216), .cin(t_6956), .o(t_6969), .co(t_6970), .cout(t_6971));
compressor_4_2 u2_2390(.a(t_1237), .b(t_1234), .c(t_1231), .d(t_1228), .cin(t_6959), .o(t_6972), .co(t_6973), .cout(t_6974));
compressor_4_2 u2_2391(.a(t_1220), .b(t_1217), .c(t_1214), .d(t_1211), .cin(t_6962), .o(t_6975), .co(t_6976), .cout(t_6977));
compressor_4_2 u2_2392(.a(t_1232), .b(t_1229), .c(t_1226), .d(t_1223), .cin(t_6965), .o(t_6978), .co(t_6979), .cout(t_6980));
compressor_4_2 u2_2393(.a(t_1243), .b(t_1240), .c(t_1238), .d(t_1235), .cin(t_6968), .o(t_6981), .co(t_6982), .cout(t_6983));
compressor_4_2 u2_2394(.a(t_1255), .b(t_1252), .c(t_1249), .d(t_1246), .cin(t_6971), .o(t_6984), .co(t_6985), .cout(t_6986));
compressor_4_2 u2_2395(.a(t_1267), .b(t_1264), .c(t_1261), .d(t_1258), .cin(t_6974), .o(t_6987), .co(t_6988), .cout(t_6989));
compressor_4_2 u2_2396(.a(t_1247), .b(t_1244), .c(t_1241), .d(s_81_40), .cin(t_6977), .o(t_6990), .co(t_6991), .cout(t_6992));
compressor_4_2 u2_2397(.a(t_1259), .b(t_1256), .c(t_1253), .d(t_1250), .cin(t_6980), .o(t_6993), .co(t_6994), .cout(t_6995));
compressor_4_2 u2_2398(.a(t_1271), .b(t_1268), .c(t_1265), .d(t_1262), .cin(t_6983), .o(t_6996), .co(t_6997), .cout(t_6998));
compressor_4_2 u2_2399(.a(t_1281), .b(t_1278), .c(t_1275), .d(t_1272), .cin(t_6986), .o(t_6999), .co(t_7000), .cout(t_7001));
compressor_4_2 u2_2400(.a(t_1293), .b(t_1290), .c(t_1287), .d(t_1284), .cin(t_6989), .o(t_7002), .co(t_7003), .cout(t_7004));
half_adder u0_2401(.a(t_1299), .b(t_1296), .o(t_7005), .cout(t_7006));
compressor_4_2 u2_2402(.a(t_1282), .b(t_1279), .c(t_1276), .d(t_1273), .cin(t_6992), .o(t_7007), .co(t_7008), .cout(t_7009));
compressor_4_2 u2_2403(.a(t_1294), .b(t_1291), .c(t_1288), .d(t_1285), .cin(t_6995), .o(t_7010), .co(t_7011), .cout(t_7012));
compressor_4_2 u2_2404(.a(t_1305), .b(t_1302), .c(t_1300), .d(t_1297), .cin(t_6998), .o(t_7013), .co(t_7014), .cout(t_7015));
compressor_4_2 u2_2405(.a(t_1317), .b(t_1314), .c(t_1311), .d(t_1308), .cin(t_7001), .o(t_7016), .co(t_7017), .cout(t_7018));
compressor_4_2 u2_2406(.a(t_1329), .b(t_1326), .c(t_1323), .d(t_1320), .cin(t_7004), .o(t_7019), .co(t_7020), .cout(t_7021));
compressor_4_2 u2_2407(.a(t_1312), .b(t_1309), .c(t_1306), .d(t_1303), .cin(t_7009), .o(t_7022), .co(t_7023), .cout(t_7024));
compressor_4_2 u2_2408(.a(t_1324), .b(t_1321), .c(t_1318), .d(t_1315), .cin(t_7012), .o(t_7025), .co(t_7026), .cout(t_7027));
compressor_4_2 u2_2409(.a(t_1334), .b(t_1333), .c(t_1330), .d(t_1327), .cin(t_7015), .o(t_7028), .co(t_7029), .cout(t_7030));
compressor_4_2 u2_2410(.a(t_1346), .b(t_1343), .c(t_1340), .d(t_1337), .cin(t_7018), .o(t_7031), .co(t_7032), .cout(t_7033));
compressor_4_2 u2_2411(.a(t_1358), .b(t_1355), .c(t_1352), .d(t_1349), .cin(t_7021), .o(t_7034), .co(t_7035), .cout(t_7036));
half_adder u0_2412(.a(t_1364), .b(t_1361), .o(t_7037), .cout(t_7038));
compressor_4_2 u2_2413(.a(t_1341), .b(t_1338), .c(t_1335), .d(s_84_43), .cin(t_7024), .o(t_7039), .co(t_7040), .cout(t_7041));
compressor_4_2 u2_2414(.a(t_1353), .b(t_1350), .c(t_1347), .d(t_1344), .cin(t_7027), .o(t_7042), .co(t_7043), .cout(t_7044));
compressor_4_2 u2_2415(.a(t_1365), .b(t_1362), .c(t_1359), .d(t_1356), .cin(t_7030), .o(t_7045), .co(t_7046), .cout(t_7047));
compressor_4_2 u2_2416(.a(t_1375), .b(t_1372), .c(t_1369), .d(t_1366), .cin(t_7033), .o(t_7048), .co(t_7049), .cout(t_7050));
compressor_4_2 u2_2417(.a(t_1387), .b(t_1384), .c(t_1381), .d(t_1378), .cin(t_7036), .o(t_7051), .co(t_7052), .cout(t_7053));
compressor_3_2 u1_2418(.a(t_1396), .b(t_1393), .cin(t_1390), .o(t_7054), .cout(t_7055));
compressor_4_2 u2_2419(.a(t_1376), .b(t_1373), .c(t_1370), .d(t_1367), .cin(t_7041), .o(t_7056), .co(t_7057), .cout(t_7058));
compressor_4_2 u2_2420(.a(t_1388), .b(t_1385), .c(t_1382), .d(t_1379), .cin(t_7044), .o(t_7059), .co(t_7060), .cout(t_7061));
compressor_4_2 u2_2421(.a(t_1398), .b(t_1397), .c(t_1394), .d(t_1391), .cin(t_7047), .o(t_7062), .co(t_7063), .cout(t_7064));
compressor_4_2 u2_2422(.a(t_1410), .b(t_1407), .c(t_1404), .d(t_1401), .cin(t_7050), .o(t_7065), .co(t_7066), .cout(t_7067));
compressor_4_2 u2_2423(.a(t_1422), .b(t_1419), .c(t_1416), .d(t_1413), .cin(t_7053), .o(t_7068), .co(t_7069), .cout(t_7070));
half_adder u0_2424(.a(t_1428), .b(t_1425), .o(t_7071), .cout(t_7072));
compressor_4_2 u2_2425(.a(t_1408), .b(t_1405), .c(t_1402), .d(t_1399), .cin(t_7058), .o(t_7073), .co(t_7074), .cout(t_7075));
compressor_4_2 u2_2426(.a(t_1420), .b(t_1417), .c(t_1414), .d(t_1411), .cin(t_7061), .o(t_7076), .co(t_7077), .cout(t_7078));
compressor_4_2 u2_2427(.a(t_1430), .b(t_1429), .c(t_1426), .d(t_1423), .cin(t_7064), .o(t_7079), .co(t_7080), .cout(t_7081));
compressor_4_2 u2_2428(.a(t_1442), .b(t_1439), .c(t_1436), .d(t_1433), .cin(t_7067), .o(t_7082), .co(t_7083), .cout(t_7084));
compressor_4_2 u2_2429(.a(t_1454), .b(t_1451), .c(t_1448), .d(t_1445), .cin(t_7070), .o(t_7085), .co(t_7086), .cout(t_7087));
half_adder u0_2430(.a(t_1460), .b(t_1457), .o(t_7088), .cout(t_7089));
compressor_4_2 u2_2431(.a(t_1440), .b(t_1437), .c(t_1434), .d(t_1431), .cin(t_7075), .o(t_7090), .co(t_7091), .cout(t_7092));
compressor_4_2 u2_2432(.a(t_1452), .b(t_1449), .c(t_1446), .d(t_1443), .cin(t_7078), .o(t_7093), .co(t_7094), .cout(t_7095));
compressor_4_2 u2_2433(.a(t_1463), .b(t_1461), .c(t_1458), .d(t_1455), .cin(t_7081), .o(t_7096), .co(t_7097), .cout(t_7098));
compressor_4_2 u2_2434(.a(t_1475), .b(t_1472), .c(t_1469), .d(t_1466), .cin(t_7084), .o(t_7099), .co(t_7100), .cout(t_7101));
compressor_4_2 u2_2435(.a(t_1487), .b(t_1484), .c(t_1481), .d(t_1478), .cin(t_7087), .o(t_7102), .co(t_7103), .cout(t_7104));
half_adder u0_2436(.a(t_1493), .b(t_1490), .o(t_7105), .cout(t_7106));
compressor_4_2 u2_2437(.a(t_1473), .b(t_1470), .c(t_1467), .d(t_1464), .cin(t_7092), .o(t_7107), .co(t_7108), .cout(t_7109));
compressor_4_2 u2_2438(.a(t_1485), .b(t_1482), .c(t_1479), .d(t_1476), .cin(t_7095), .o(t_7110), .co(t_7111), .cout(t_7112));
compressor_4_2 u2_2439(.a(t_1496), .b(t_1494), .c(t_1491), .d(t_1488), .cin(t_7098), .o(t_7113), .co(t_7114), .cout(t_7115));
compressor_4_2 u2_2440(.a(t_1508), .b(t_1505), .c(t_1502), .d(t_1499), .cin(t_7101), .o(t_7116), .co(t_7117), .cout(t_7118));
compressor_4_2 u2_2441(.a(t_1520), .b(t_1517), .c(t_1514), .d(t_1511), .cin(t_7104), .o(t_7119), .co(t_7120), .cout(t_7121));
compressor_3_2 u1_2442(.a(t_1529), .b(t_1526), .cin(t_1523), .o(t_7122), .cout(t_7123));
compressor_4_2 u2_2443(.a(t_1503), .b(t_1500), .c(t_1497), .d(s_89_44), .cin(t_7109), .o(t_7124), .co(t_7125), .cout(t_7126));
compressor_4_2 u2_2444(.a(t_1515), .b(t_1512), .c(t_1509), .d(t_1506), .cin(t_7112), .o(t_7127), .co(t_7128), .cout(t_7129));
compressor_4_2 u2_2445(.a(t_1527), .b(t_1524), .c(t_1521), .d(t_1518), .cin(t_7115), .o(t_7130), .co(t_7131), .cout(t_7132));
compressor_4_2 u2_2446(.a(t_1537), .b(t_1534), .c(t_1531), .d(t_1530), .cin(t_7118), .o(t_7133), .co(t_7134), .cout(t_7135));
compressor_4_2 u2_2447(.a(t_1549), .b(t_1546), .c(t_1543), .d(t_1540), .cin(t_7121), .o(t_7136), .co(t_7137), .cout(t_7138));
compressor_3_2 u1_2448(.a(t_1558), .b(t_1555), .cin(t_1552), .o(t_7139), .cout(t_7140));
compressor_4_2 u2_2449(.a(t_1541), .b(t_1538), .c(t_1535), .d(t_1532), .cin(t_7126), .o(t_7141), .co(t_7142), .cout(t_7143));
compressor_4_2 u2_2450(.a(t_1553), .b(t_1550), .c(t_1547), .d(t_1544), .cin(t_7129), .o(t_7144), .co(t_7145), .cout(t_7146));
compressor_4_2 u2_2451(.a(t_1564), .b(t_1562), .c(t_1559), .d(t_1556), .cin(t_7132), .o(t_7147), .co(t_7148), .cout(t_7149));
compressor_4_2 u2_2452(.a(t_1576), .b(t_1573), .c(t_1570), .d(t_1567), .cin(t_7135), .o(t_7150), .co(t_7151), .cout(t_7152));
compressor_4_2 u2_2453(.a(t_1588), .b(t_1585), .c(t_1582), .d(t_1579), .cin(t_7138), .o(t_7153), .co(t_7154), .cout(t_7155));
compressor_3_2 u1_2454(.a(t_1597), .b(t_1594), .cin(t_1591), .o(t_7156), .cout(t_7157));
compressor_4_2 u2_2455(.a(t_1574), .b(t_1571), .c(t_1568), .d(t_1565), .cin(t_7143), .o(t_7158), .co(t_7159), .cout(t_7160));
compressor_4_2 u2_2456(.a(t_1586), .b(t_1583), .c(t_1580), .d(t_1577), .cin(t_7146), .o(t_7161), .co(t_7162), .cout(t_7163));
compressor_4_2 u2_2457(.a(t_1598), .b(t_1595), .c(t_1592), .d(t_1589), .cin(t_7149), .o(t_7164), .co(t_7165), .cout(t_7166));
compressor_4_2 u2_2458(.a(t_1608), .b(t_1605), .c(t_1602), .d(t_1599), .cin(t_7152), .o(t_7167), .co(t_7168), .cout(t_7169));
compressor_4_2 u2_2459(.a(t_1620), .b(t_1617), .c(t_1614), .d(t_1611), .cin(t_7155), .o(t_7170), .co(t_7171), .cout(t_7172));
compressor_3_2 u1_2460(.a(t_1629), .b(t_1626), .cin(t_1623), .o(t_7173), .cout(t_7174));
compressor_4_2 u2_2461(.a(t_1606), .b(t_1603), .c(t_1600), .d(s_92_47), .cin(t_7160), .o(t_7175), .co(t_7176), .cout(t_7177));
compressor_4_2 u2_2462(.a(t_1618), .b(t_1615), .c(t_1612), .d(t_1609), .cin(t_7163), .o(t_7178), .co(t_7179), .cout(t_7180));
compressor_4_2 u2_2463(.a(t_1630), .b(t_1627), .c(t_1624), .d(t_1621), .cin(t_7166), .o(t_7181), .co(t_7182), .cout(t_7183));
compressor_4_2 u2_2464(.a(t_1640), .b(t_1637), .c(t_1634), .d(t_1633), .cin(t_7169), .o(t_7184), .co(t_7185), .cout(t_7186));
compressor_4_2 u2_2465(.a(t_1652), .b(t_1649), .c(t_1646), .d(t_1643), .cin(t_7172), .o(t_7187), .co(t_7188), .cout(t_7189));
compressor_4_2 u2_2466(.a(t_1667), .b(t_1664), .c(t_1661), .d(t_1658), .cin(t_1655), .o(t_7190), .co(t_7191), .cout(t_7192));
compressor_4_2 u2_2467(.a(t_1644), .b(t_1641), .c(t_1638), .d(t_1635), .cin(t_7177), .o(t_7193), .co(t_7194), .cout(t_7195));
compressor_4_2 u2_2468(.a(t_1656), .b(t_1653), .c(t_1650), .d(t_1647), .cin(t_7180), .o(t_7196), .co(t_7197), .cout(t_7198));
compressor_4_2 u2_2469(.a(t_1668), .b(t_1665), .c(t_1662), .d(t_1659), .cin(t_7183), .o(t_7199), .co(t_7200), .cout(t_7201));
compressor_4_2 u2_2470(.a(t_1678), .b(t_1675), .c(t_1672), .d(t_1669), .cin(t_7186), .o(t_7202), .co(t_7203), .cout(t_7204));
compressor_4_2 u2_2471(.a(t_1690), .b(t_1687), .c(t_1684), .d(t_1681), .cin(t_7189), .o(t_7205), .co(t_7206), .cout(t_7207));
compressor_4_2 u2_2472(.a(t_1702), .b(t_1699), .c(t_1696), .d(t_1693), .cin(t_7192), .o(t_7208), .co(t_7209), .cout(t_7210));
compressor_4_2 u2_2473(.a(t_1679), .b(t_1676), .c(t_1673), .d(t_1670), .cin(t_7195), .o(t_7211), .co(t_7212), .cout(t_7213));
compressor_4_2 u2_2474(.a(t_1691), .b(t_1688), .c(t_1685), .d(t_1682), .cin(t_7198), .o(t_7214), .co(t_7215), .cout(t_7216));
compressor_4_2 u2_2475(.a(t_1703), .b(t_1700), .c(t_1697), .d(t_1694), .cin(t_7201), .o(t_7217), .co(t_7218), .cout(t_7219));
compressor_4_2 u2_2476(.a(t_1713), .b(t_1710), .c(t_1707), .d(t_1704), .cin(t_7204), .o(t_7220), .co(t_7221), .cout(t_7222));
compressor_4_2 u2_2477(.a(t_1725), .b(t_1722), .c(t_1719), .d(t_1716), .cin(t_7207), .o(t_7223), .co(t_7224), .cout(t_7225));
compressor_4_2 u2_2478(.a(t_1737), .b(t_1734), .c(t_1731), .d(t_1728), .cin(t_7210), .o(t_7226), .co(t_7227), .cout(t_7228));
compressor_4_2 u2_2479(.a(t_1714), .b(t_1711), .c(t_1708), .d(t_1705), .cin(t_7213), .o(t_7229), .co(t_7230), .cout(t_7231));
compressor_4_2 u2_2480(.a(t_1726), .b(t_1723), .c(t_1720), .d(t_1717), .cin(t_7216), .o(t_7232), .co(t_7233), .cout(t_7234));
compressor_4_2 u2_2481(.a(t_1738), .b(t_1735), .c(t_1732), .d(t_1729), .cin(t_7219), .o(t_7235), .co(t_7236), .cout(t_7237));
compressor_4_2 u2_2482(.a(t_1749), .b(t_1746), .c(t_1743), .d(t_1740), .cin(t_7222), .o(t_7238), .co(t_7239), .cout(t_7240));
compressor_4_2 u2_2483(.a(t_1761), .b(t_1758), .c(t_1755), .d(t_1752), .cin(t_7225), .o(t_7241), .co(t_7242), .cout(t_7243));
compressor_4_2 u2_2484(.a(t_1773), .b(t_1770), .c(t_1767), .d(t_1764), .cin(t_7228), .o(t_7244), .co(t_7245), .cout(t_7246));
compressor_4_2 u2_2485(.a(t_1750), .b(t_1747), .c(t_1744), .d(t_1741), .cin(t_7231), .o(t_7247), .co(t_7248), .cout(t_7249));
compressor_4_2 u2_2486(.a(t_1762), .b(t_1759), .c(t_1756), .d(t_1753), .cin(t_7234), .o(t_7250), .co(t_7251), .cout(t_7252));
compressor_4_2 u2_2487(.a(t_1774), .b(t_1771), .c(t_1768), .d(t_1765), .cin(t_7237), .o(t_7253), .co(t_7254), .cout(t_7255));
compressor_4_2 u2_2488(.a(t_1785), .b(t_1782), .c(t_1779), .d(t_1776), .cin(t_7240), .o(t_7256), .co(t_7257), .cout(t_7258));
compressor_4_2 u2_2489(.a(t_1797), .b(t_1794), .c(t_1791), .d(t_1788), .cin(t_7243), .o(t_7259), .co(t_7260), .cout(t_7261));
compressor_4_2 u2_2490(.a(t_1809), .b(t_1806), .c(t_1803), .d(t_1800), .cin(t_7246), .o(t_7262), .co(t_7263), .cout(t_7264));
compressor_4_2 u2_2491(.a(t_1783), .b(t_1780), .c(t_1777), .d(s_97_48), .cin(t_7249), .o(t_7265), .co(t_7266), .cout(t_7267));
compressor_4_2 u2_2492(.a(t_1795), .b(t_1792), .c(t_1789), .d(t_1786), .cin(t_7252), .o(t_7268), .co(t_7269), .cout(t_7270));
compressor_4_2 u2_2493(.a(t_1807), .b(t_1804), .c(t_1801), .d(t_1798), .cin(t_7255), .o(t_7271), .co(t_7272), .cout(t_7273));
compressor_4_2 u2_2494(.a(t_1817), .b(t_1814), .c(t_1813), .d(t_1810), .cin(t_7258), .o(t_7274), .co(t_7275), .cout(t_7276));
compressor_4_2 u2_2495(.a(t_1829), .b(t_1826), .c(t_1823), .d(t_1820), .cin(t_7261), .o(t_7277), .co(t_7278), .cout(t_7279));
compressor_4_2 u2_2496(.a(t_1841), .b(t_1838), .c(t_1835), .d(t_1832), .cin(t_7264), .o(t_7280), .co(t_7281), .cout(t_7282));
half_adder u0_2497(.a(t_1847), .b(t_1844), .o(t_7283), .cout(t_7284));
compressor_4_2 u2_2498(.a(t_1824), .b(t_1821), .c(t_1818), .d(t_1815), .cin(t_7267), .o(t_7285), .co(t_7286), .cout(t_7287));
compressor_4_2 u2_2499(.a(t_1836), .b(t_1833), .c(t_1830), .d(t_1827), .cin(t_7270), .o(t_7288), .co(t_7289), .cout(t_7290));
compressor_4_2 u2_2500(.a(t_1848), .b(t_1845), .c(t_1842), .d(t_1839), .cin(t_7273), .o(t_7291), .co(t_7292), .cout(t_7293));
compressor_4_2 u2_2501(.a(t_1859), .b(t_1856), .c(t_1853), .d(t_1850), .cin(t_7276), .o(t_7294), .co(t_7295), .cout(t_7296));
compressor_4_2 u2_2502(.a(t_1871), .b(t_1868), .c(t_1865), .d(t_1862), .cin(t_7279), .o(t_7297), .co(t_7298), .cout(t_7299));
compressor_4_2 u2_2503(.a(t_1883), .b(t_1880), .c(t_1877), .d(t_1874), .cin(t_7282), .o(t_7300), .co(t_7301), .cout(t_7302));
compressor_4_2 u2_2504(.a(t_1860), .b(t_1857), .c(t_1854), .d(t_1851), .cin(t_7287), .o(t_7303), .co(t_7304), .cout(t_7305));
compressor_4_2 u2_2505(.a(t_1872), .b(t_1869), .c(t_1866), .d(t_1863), .cin(t_7290), .o(t_7306), .co(t_7307), .cout(t_7308));
compressor_4_2 u2_2506(.a(t_1884), .b(t_1881), .c(t_1878), .d(t_1875), .cin(t_7293), .o(t_7309), .co(t_7310), .cout(t_7311));
compressor_4_2 u2_2507(.a(t_1894), .b(t_1891), .c(t_1888), .d(t_1887), .cin(t_7296), .o(t_7312), .co(t_7313), .cout(t_7314));
compressor_4_2 u2_2508(.a(t_1906), .b(t_1903), .c(t_1900), .d(t_1897), .cin(t_7299), .o(t_7315), .co(t_7316), .cout(t_7317));
compressor_4_2 u2_2509(.a(t_1918), .b(t_1915), .c(t_1912), .d(t_1909), .cin(t_7302), .o(t_7318), .co(t_7319), .cout(t_7320));
half_adder u0_2510(.a(t_1924), .b(t_1921), .o(t_7321), .cout(t_7322));
compressor_4_2 u2_2511(.a(t_1895), .b(t_1892), .c(t_1889), .d(s_100_51), .cin(t_7305), .o(t_7323), .co(t_7324), .cout(t_7325));
compressor_4_2 u2_2512(.a(t_1907), .b(t_1904), .c(t_1901), .d(t_1898), .cin(t_7308), .o(t_7326), .co(t_7327), .cout(t_7328));
compressor_4_2 u2_2513(.a(t_1919), .b(t_1916), .c(t_1913), .d(t_1910), .cin(t_7311), .o(t_7329), .co(t_7330), .cout(t_7331));
compressor_4_2 u2_2514(.a(t_1929), .b(t_1926), .c(t_1925), .d(t_1922), .cin(t_7314), .o(t_7332), .co(t_7333), .cout(t_7334));
compressor_4_2 u2_2515(.a(t_1941), .b(t_1938), .c(t_1935), .d(t_1932), .cin(t_7317), .o(t_7335), .co(t_7336), .cout(t_7337));
compressor_4_2 u2_2516(.a(t_1953), .b(t_1950), .c(t_1947), .d(t_1944), .cin(t_7320), .o(t_7338), .co(t_7339), .cout(t_7340));
compressor_3_2 u1_2517(.a(t_1962), .b(t_1959), .cin(t_1956), .o(t_7341), .cout(t_7342));
compressor_4_2 u2_2518(.a(t_1936), .b(t_1933), .c(t_1930), .d(t_1927), .cin(t_7325), .o(t_7343), .co(t_7344), .cout(t_7345));
compressor_4_2 u2_2519(.a(t_1948), .b(t_1945), .c(t_1942), .d(t_1939), .cin(t_7328), .o(t_7346), .co(t_7347), .cout(t_7348));
compressor_4_2 u2_2520(.a(t_1960), .b(t_1957), .c(t_1954), .d(t_1951), .cin(t_7331), .o(t_7349), .co(t_7350), .cout(t_7351));
compressor_4_2 u2_2521(.a(t_1970), .b(t_1967), .c(t_1964), .d(t_1963), .cin(t_7334), .o(t_7352), .co(t_7353), .cout(t_7354));
compressor_4_2 u2_2522(.a(t_1982), .b(t_1979), .c(t_1976), .d(t_1973), .cin(t_7337), .o(t_7355), .co(t_7356), .cout(t_7357));
compressor_4_2 u2_2523(.a(t_1994), .b(t_1991), .c(t_1988), .d(t_1985), .cin(t_7340), .o(t_7358), .co(t_7359), .cout(t_7360));
half_adder u0_2524(.a(t_2000), .b(t_1997), .o(t_7361), .cout(t_7362));
compressor_4_2 u2_2525(.a(t_1974), .b(t_1971), .c(t_1968), .d(t_1965), .cin(t_7345), .o(t_7363), .co(t_7364), .cout(t_7365));
compressor_4_2 u2_2526(.a(t_1986), .b(t_1983), .c(t_1980), .d(t_1977), .cin(t_7348), .o(t_7366), .co(t_7367), .cout(t_7368));
compressor_4_2 u2_2527(.a(t_1998), .b(t_1995), .c(t_1992), .d(t_1989), .cin(t_7351), .o(t_7369), .co(t_7370), .cout(t_7371));
compressor_4_2 u2_2528(.a(t_2008), .b(t_2005), .c(t_2002), .d(t_2001), .cin(t_7354), .o(t_7372), .co(t_7373), .cout(t_7374));
compressor_4_2 u2_2529(.a(t_2020), .b(t_2017), .c(t_2014), .d(t_2011), .cin(t_7357), .o(t_7375), .co(t_7376), .cout(t_7377));
compressor_4_2 u2_2530(.a(t_2032), .b(t_2029), .c(t_2026), .d(t_2023), .cin(t_7360), .o(t_7378), .co(t_7379), .cout(t_7380));
half_adder u0_2531(.a(t_2038), .b(t_2035), .o(t_7381), .cout(t_7382));
compressor_4_2 u2_2532(.a(t_2012), .b(t_2009), .c(t_2006), .d(t_2003), .cin(t_7365), .o(t_7383), .co(t_7384), .cout(t_7385));
compressor_4_2 u2_2533(.a(t_2024), .b(t_2021), .c(t_2018), .d(t_2015), .cin(t_7368), .o(t_7386), .co(t_7387), .cout(t_7388));
compressor_4_2 u2_2534(.a(t_2036), .b(t_2033), .c(t_2030), .d(t_2027), .cin(t_7371), .o(t_7389), .co(t_7390), .cout(t_7391));
compressor_4_2 u2_2535(.a(t_2047), .b(t_2044), .c(t_2041), .d(t_2039), .cin(t_7374), .o(t_7392), .co(t_7393), .cout(t_7394));
compressor_4_2 u2_2536(.a(t_2059), .b(t_2056), .c(t_2053), .d(t_2050), .cin(t_7377), .o(t_7395), .co(t_7396), .cout(t_7397));
compressor_4_2 u2_2537(.a(t_2071), .b(t_2068), .c(t_2065), .d(t_2062), .cin(t_7380), .o(t_7398), .co(t_7399), .cout(t_7400));
half_adder u0_2538(.a(t_2077), .b(t_2074), .o(t_7401), .cout(t_7402));
compressor_4_2 u2_2539(.a(t_2051), .b(t_2048), .c(t_2045), .d(t_2042), .cin(t_7385), .o(t_7403), .co(t_7404), .cout(t_7405));
compressor_4_2 u2_2540(.a(t_2063), .b(t_2060), .c(t_2057), .d(t_2054), .cin(t_7388), .o(t_7406), .co(t_7407), .cout(t_7408));
compressor_4_2 u2_2541(.a(t_2075), .b(t_2072), .c(t_2069), .d(t_2066), .cin(t_7391), .o(t_7409), .co(t_7410), .cout(t_7411));
compressor_4_2 u2_2542(.a(t_2086), .b(t_2083), .c(t_2080), .d(t_2078), .cin(t_7394), .o(t_7412), .co(t_7413), .cout(t_7414));
compressor_4_2 u2_2543(.a(t_2098), .b(t_2095), .c(t_2092), .d(t_2089), .cin(t_7397), .o(t_7415), .co(t_7416), .cout(t_7417));
compressor_4_2 u2_2544(.a(t_2110), .b(t_2107), .c(t_2104), .d(t_2101), .cin(t_7400), .o(t_7418), .co(t_7419), .cout(t_7420));
compressor_3_2 u1_2545(.a(t_2119), .b(t_2116), .cin(t_2113), .o(t_7421), .cout(t_7422));
compressor_4_2 u2_2546(.a(t_2087), .b(t_2084), .c(t_2081), .d(s_105_52), .cin(t_7405), .o(t_7423), .co(t_7424), .cout(t_7425));
compressor_4_2 u2_2547(.a(t_2099), .b(t_2096), .c(t_2093), .d(t_2090), .cin(t_7408), .o(t_7426), .co(t_7427), .cout(t_7428));
compressor_4_2 u2_2548(.a(t_2111), .b(t_2108), .c(t_2105), .d(t_2102), .cin(t_7411), .o(t_7429), .co(t_7430), .cout(t_7431));
compressor_4_2 u2_2549(.a(t_2121), .b(t_2120), .c(t_2117), .d(t_2114), .cin(t_7414), .o(t_7432), .co(t_7433), .cout(t_7434));
compressor_4_2 u2_2550(.a(t_2133), .b(t_2130), .c(t_2127), .d(t_2124), .cin(t_7417), .o(t_7435), .co(t_7436), .cout(t_7437));
compressor_4_2 u2_2551(.a(t_2145), .b(t_2142), .c(t_2139), .d(t_2136), .cin(t_7420), .o(t_7438), .co(t_7439), .cout(t_7440));
compressor_3_2 u1_2552(.a(t_2154), .b(t_2151), .cin(t_2148), .o(t_7441), .cout(t_7442));
compressor_4_2 u2_2553(.a(t_2131), .b(t_2128), .c(t_2125), .d(t_2122), .cin(t_7425), .o(t_7443), .co(t_7444), .cout(t_7445));
compressor_4_2 u2_2554(.a(t_2143), .b(t_2140), .c(t_2137), .d(t_2134), .cin(t_7428), .o(t_7446), .co(t_7447), .cout(t_7448));
compressor_4_2 u2_2555(.a(t_2155), .b(t_2152), .c(t_2149), .d(t_2146), .cin(t_7431), .o(t_7449), .co(t_7450), .cout(t_7451));
compressor_4_2 u2_2556(.a(t_2166), .b(t_2163), .c(t_2160), .d(t_2158), .cin(t_7434), .o(t_7452), .co(t_7453), .cout(t_7454));
compressor_4_2 u2_2557(.a(t_2178), .b(t_2175), .c(t_2172), .d(t_2169), .cin(t_7437), .o(t_7455), .co(t_7456), .cout(t_7457));
compressor_4_2 u2_2558(.a(t_2190), .b(t_2187), .c(t_2184), .d(t_2181), .cin(t_7440), .o(t_7458), .co(t_7459), .cout(t_7460));
compressor_3_2 u1_2559(.a(t_2199), .b(t_2196), .cin(t_2193), .o(t_7461), .cout(t_7462));
compressor_4_2 u2_2560(.a(t_2170), .b(t_2167), .c(t_2164), .d(t_2161), .cin(t_7445), .o(t_7463), .co(t_7464), .cout(t_7465));
compressor_4_2 u2_2561(.a(t_2182), .b(t_2179), .c(t_2176), .d(t_2173), .cin(t_7448), .o(t_7466), .co(t_7467), .cout(t_7468));
compressor_4_2 u2_2562(.a(t_2194), .b(t_2191), .c(t_2188), .d(t_2185), .cin(t_7451), .o(t_7469), .co(t_7470), .cout(t_7471));
compressor_4_2 u2_2563(.a(t_2204), .b(t_2201), .c(t_2200), .d(t_2197), .cin(t_7454), .o(t_7472), .co(t_7473), .cout(t_7474));
compressor_4_2 u2_2564(.a(t_2216), .b(t_2213), .c(t_2210), .d(t_2207), .cin(t_7457), .o(t_7475), .co(t_7476), .cout(t_7477));
compressor_4_2 u2_2565(.a(t_2228), .b(t_2225), .c(t_2222), .d(t_2219), .cin(t_7460), .o(t_7478), .co(t_7479), .cout(t_7480));
compressor_3_2 u1_2566(.a(t_2237), .b(t_2234), .cin(t_2231), .o(t_7481), .cout(t_7482));
compressor_4_2 u2_2567(.a(t_2208), .b(t_2205), .c(t_2202), .d(s_108_55), .cin(t_7465), .o(t_7483), .co(t_7484), .cout(t_7485));
compressor_4_2 u2_2568(.a(t_2220), .b(t_2217), .c(t_2214), .d(t_2211), .cin(t_7468), .o(t_7486), .co(t_7487), .cout(t_7488));
compressor_4_2 u2_2569(.a(t_2232), .b(t_2229), .c(t_2226), .d(t_2223), .cin(t_7471), .o(t_7489), .co(t_7490), .cout(t_7491));
compressor_4_2 u2_2570(.a(t_2242), .b(t_2241), .c(t_2238), .d(t_2235), .cin(t_7474), .o(t_7492), .co(t_7493), .cout(t_7494));
compressor_4_2 u2_2571(.a(t_2254), .b(t_2251), .c(t_2248), .d(t_2245), .cin(t_7477), .o(t_7495), .co(t_7496), .cout(t_7497));
compressor_4_2 u2_2572(.a(t_2266), .b(t_2263), .c(t_2260), .d(t_2257), .cin(t_7480), .o(t_7498), .co(t_7499), .cout(t_7500));
compressor_4_2 u2_2573(.a(t_2281), .b(t_2278), .c(t_2275), .d(t_2272), .cin(t_2269), .o(t_7501), .co(t_7502), .cout(t_7503));
compressor_4_2 u2_2574(.a(t_2252), .b(t_2249), .c(t_2246), .d(t_2243), .cin(t_7485), .o(t_7504), .co(t_7505), .cout(t_7506));
compressor_4_2 u2_2575(.a(t_2264), .b(t_2261), .c(t_2258), .d(t_2255), .cin(t_7488), .o(t_7507), .co(t_7508), .cout(t_7509));
compressor_4_2 u2_2576(.a(t_2276), .b(t_2273), .c(t_2270), .d(t_2267), .cin(t_7491), .o(t_7510), .co(t_7511), .cout(t_7512));
compressor_4_2 u2_2577(.a(t_2286), .b(t_2283), .c(t_2282), .d(t_2279), .cin(t_7494), .o(t_7513), .co(t_7514), .cout(t_7515));
compressor_4_2 u2_2578(.a(t_2298), .b(t_2295), .c(t_2292), .d(t_2289), .cin(t_7497), .o(t_7516), .co(t_7517), .cout(t_7518));
compressor_4_2 u2_2579(.a(t_2310), .b(t_2307), .c(t_2304), .d(t_2301), .cin(t_7500), .o(t_7519), .co(t_7520), .cout(t_7521));
compressor_4_2 u2_2580(.a(t_2322), .b(t_2319), .c(t_2316), .d(t_2313), .cin(t_7503), .o(t_7522), .co(t_7523), .cout(t_7524));
compressor_4_2 u2_2581(.a(t_2293), .b(t_2290), .c(t_2287), .d(t_2284), .cin(t_7506), .o(t_7525), .co(t_7526), .cout(t_7527));
compressor_4_2 u2_2582(.a(t_2305), .b(t_2302), .c(t_2299), .d(t_2296), .cin(t_7509), .o(t_7528), .co(t_7529), .cout(t_7530));
compressor_4_2 u2_2583(.a(t_2317), .b(t_2314), .c(t_2311), .d(t_2308), .cin(t_7512), .o(t_7531), .co(t_7532), .cout(t_7533));
compressor_4_2 u2_2584(.a(t_2327), .b(t_2324), .c(t_2323), .d(t_2320), .cin(t_7515), .o(t_7534), .co(t_7535), .cout(t_7536));
compressor_4_2 u2_2585(.a(t_2339), .b(t_2336), .c(t_2333), .d(t_2330), .cin(t_7518), .o(t_7537), .co(t_7538), .cout(t_7539));
compressor_4_2 u2_2586(.a(t_2351), .b(t_2348), .c(t_2345), .d(t_2342), .cin(t_7521), .o(t_7540), .co(t_7541), .cout(t_7542));
compressor_4_2 u2_2587(.a(t_2363), .b(t_2360), .c(t_2357), .d(t_2354), .cin(t_7524), .o(t_7543), .co(t_7544), .cout(t_7545));
compressor_4_2 u2_2588(.a(t_2334), .b(t_2331), .c(t_2328), .d(t_2325), .cin(t_7527), .o(t_7546), .co(t_7547), .cout(t_7548));
compressor_4_2 u2_2589(.a(t_2346), .b(t_2343), .c(t_2340), .d(t_2337), .cin(t_7530), .o(t_7549), .co(t_7550), .cout(t_7551));
compressor_4_2 u2_2590(.a(t_2358), .b(t_2355), .c(t_2352), .d(t_2349), .cin(t_7533), .o(t_7552), .co(t_7553), .cout(t_7554));
compressor_4_2 u2_2591(.a(t_2369), .b(t_2366), .c(t_2364), .d(t_2361), .cin(t_7536), .o(t_7555), .co(t_7556), .cout(t_7557));
compressor_4_2 u2_2592(.a(t_2381), .b(t_2378), .c(t_2375), .d(t_2372), .cin(t_7539), .o(t_7558), .co(t_7559), .cout(t_7560));
compressor_4_2 u2_2593(.a(t_2393), .b(t_2390), .c(t_2387), .d(t_2384), .cin(t_7542), .o(t_7561), .co(t_7562), .cout(t_7563));
compressor_4_2 u2_2594(.a(t_2405), .b(t_2402), .c(t_2399), .d(t_2396), .cin(t_7545), .o(t_7564), .co(t_7565), .cout(t_7566));
compressor_4_2 u2_2595(.a(t_2376), .b(t_2373), .c(t_2370), .d(t_2367), .cin(t_7548), .o(t_7567), .co(t_7568), .cout(t_7569));
compressor_4_2 u2_2596(.a(t_2388), .b(t_2385), .c(t_2382), .d(t_2379), .cin(t_7551), .o(t_7570), .co(t_7571), .cout(t_7572));
compressor_4_2 u2_2597(.a(t_2400), .b(t_2397), .c(t_2394), .d(t_2391), .cin(t_7554), .o(t_7573), .co(t_7574), .cout(t_7575));
compressor_4_2 u2_2598(.a(t_2411), .b(t_2408), .c(t_2406), .d(t_2403), .cin(t_7557), .o(t_7576), .co(t_7577), .cout(t_7578));
compressor_4_2 u2_2599(.a(t_2423), .b(t_2420), .c(t_2417), .d(t_2414), .cin(t_7560), .o(t_7579), .co(t_7580), .cout(t_7581));
compressor_4_2 u2_2600(.a(t_2435), .b(t_2432), .c(t_2429), .d(t_2426), .cin(t_7563), .o(t_7582), .co(t_7583), .cout(t_7584));
compressor_4_2 u2_2601(.a(t_2447), .b(t_2444), .c(t_2441), .d(t_2438), .cin(t_7566), .o(t_7585), .co(t_7586), .cout(t_7587));
compressor_4_2 u2_2602(.a(t_2415), .b(t_2412), .c(t_2409), .d(s_113_56), .cin(t_7569), .o(t_7588), .co(t_7589), .cout(t_7590));
compressor_4_2 u2_2603(.a(t_2427), .b(t_2424), .c(t_2421), .d(t_2418), .cin(t_7572), .o(t_7591), .co(t_7592), .cout(t_7593));
compressor_4_2 u2_2604(.a(t_2439), .b(t_2436), .c(t_2433), .d(t_2430), .cin(t_7575), .o(t_7594), .co(t_7595), .cout(t_7596));
compressor_4_2 u2_2605(.a(t_2451), .b(t_2448), .c(t_2445), .d(t_2442), .cin(t_7578), .o(t_7597), .co(t_7598), .cout(t_7599));
compressor_4_2 u2_2606(.a(t_2461), .b(t_2458), .c(t_2455), .d(t_2452), .cin(t_7581), .o(t_7600), .co(t_7601), .cout(t_7602));
compressor_4_2 u2_2607(.a(t_2473), .b(t_2470), .c(t_2467), .d(t_2464), .cin(t_7584), .o(t_7603), .co(t_7604), .cout(t_7605));
compressor_4_2 u2_2608(.a(t_2485), .b(t_2482), .c(t_2479), .d(t_2476), .cin(t_7587), .o(t_7606), .co(t_7607), .cout(t_7608));
half_adder u0_2609(.a(t_2491), .b(t_2488), .o(t_7609), .cout(t_7610));
compressor_4_2 u2_2610(.a(t_2462), .b(t_2459), .c(t_2456), .d(t_2453), .cin(t_7590), .o(t_7611), .co(t_7612), .cout(t_7613));
compressor_4_2 u2_2611(.a(t_2474), .b(t_2471), .c(t_2468), .d(t_2465), .cin(t_7593), .o(t_7614), .co(t_7615), .cout(t_7616));
compressor_4_2 u2_2612(.a(t_2486), .b(t_2483), .c(t_2480), .d(t_2477), .cin(t_7596), .o(t_7617), .co(t_7618), .cout(t_7619));
compressor_4_2 u2_2613(.a(t_2497), .b(t_2494), .c(t_2492), .d(t_2489), .cin(t_7599), .o(t_7620), .co(t_7621), .cout(t_7622));
compressor_4_2 u2_2614(.a(t_2509), .b(t_2506), .c(t_2503), .d(t_2500), .cin(t_7602), .o(t_7623), .co(t_7624), .cout(t_7625));
compressor_4_2 u2_2615(.a(t_2521), .b(t_2518), .c(t_2515), .d(t_2512), .cin(t_7605), .o(t_7626), .co(t_7627), .cout(t_7628));
compressor_4_2 u2_2616(.a(t_2533), .b(t_2530), .c(t_2527), .d(t_2524), .cin(t_7608), .o(t_7629), .co(t_7630), .cout(t_7631));
compressor_4_2 u2_2617(.a(t_2504), .b(t_2501), .c(t_2498), .d(t_2495), .cin(t_7613), .o(t_7632), .co(t_7633), .cout(t_7634));
compressor_4_2 u2_2618(.a(t_2516), .b(t_2513), .c(t_2510), .d(t_2507), .cin(t_7616), .o(t_7635), .co(t_7636), .cout(t_7637));
compressor_4_2 u2_2619(.a(t_2528), .b(t_2525), .c(t_2522), .d(t_2519), .cin(t_7619), .o(t_7638), .co(t_7639), .cout(t_7640));
compressor_4_2 u2_2620(.a(t_2538), .b(t_2537), .c(t_2534), .d(t_2531), .cin(t_7622), .o(t_7641), .co(t_7642), .cout(t_7643));
compressor_4_2 u2_2621(.a(t_2550), .b(t_2547), .c(t_2544), .d(t_2541), .cin(t_7625), .o(t_7644), .co(t_7645), .cout(t_7646));
compressor_4_2 u2_2622(.a(t_2562), .b(t_2559), .c(t_2556), .d(t_2553), .cin(t_7628), .o(t_7647), .co(t_7648), .cout(t_7649));
compressor_4_2 u2_2623(.a(t_2574), .b(t_2571), .c(t_2568), .d(t_2565), .cin(t_7631), .o(t_7650), .co(t_7651), .cout(t_7652));
half_adder u0_2624(.a(t_2580), .b(t_2577), .o(t_7653), .cout(t_7654));
compressor_4_2 u2_2625(.a(t_2545), .b(t_2542), .c(t_2539), .d(s_116_59), .cin(t_7634), .o(t_7655), .co(t_7656), .cout(t_7657));
compressor_4_2 u2_2626(.a(t_2557), .b(t_2554), .c(t_2551), .d(t_2548), .cin(t_7637), .o(t_7658), .co(t_7659), .cout(t_7660));
compressor_4_2 u2_2627(.a(t_2569), .b(t_2566), .c(t_2563), .d(t_2560), .cin(t_7640), .o(t_7661), .co(t_7662), .cout(t_7663));
compressor_4_2 u2_2628(.a(t_2581), .b(t_2578), .c(t_2575), .d(t_2572), .cin(t_7643), .o(t_7664), .co(t_7665), .cout(t_7666));
compressor_4_2 u2_2629(.a(t_2591), .b(t_2588), .c(t_2585), .d(t_2582), .cin(t_7646), .o(t_7667), .co(t_7668), .cout(t_7669));
compressor_4_2 u2_2630(.a(t_2603), .b(t_2600), .c(t_2597), .d(t_2594), .cin(t_7649), .o(t_7670), .co(t_7671), .cout(t_7672));
compressor_4_2 u2_2631(.a(t_2615), .b(t_2612), .c(t_2609), .d(t_2606), .cin(t_7652), .o(t_7673), .co(t_7674), .cout(t_7675));
compressor_3_2 u1_2632(.a(t_2624), .b(t_2621), .cin(t_2618), .o(t_7676), .cout(t_7677));
compressor_4_2 u2_2633(.a(t_2592), .b(t_2589), .c(t_2586), .d(t_2583), .cin(t_7657), .o(t_7678), .co(t_7679), .cout(t_7680));
compressor_4_2 u2_2634(.a(t_2604), .b(t_2601), .c(t_2598), .d(t_2595), .cin(t_7660), .o(t_7681), .co(t_7682), .cout(t_7683));
compressor_4_2 u2_2635(.a(t_2616), .b(t_2613), .c(t_2610), .d(t_2607), .cin(t_7663), .o(t_7684), .co(t_7685), .cout(t_7686));
compressor_4_2 u2_2636(.a(t_2626), .b(t_2625), .c(t_2622), .d(t_2619), .cin(t_7666), .o(t_7687), .co(t_7688), .cout(t_7689));
compressor_4_2 u2_2637(.a(t_2638), .b(t_2635), .c(t_2632), .d(t_2629), .cin(t_7669), .o(t_7690), .co(t_7691), .cout(t_7692));
compressor_4_2 u2_2638(.a(t_2650), .b(t_2647), .c(t_2644), .d(t_2641), .cin(t_7672), .o(t_7693), .co(t_7694), .cout(t_7695));
compressor_4_2 u2_2639(.a(t_2662), .b(t_2659), .c(t_2656), .d(t_2653), .cin(t_7675), .o(t_7696), .co(t_7697), .cout(t_7698));
half_adder u0_2640(.a(t_2668), .b(t_2665), .o(t_7699), .cout(t_7700));
compressor_4_2 u2_2641(.a(t_2636), .b(t_2633), .c(t_2630), .d(t_2627), .cin(t_7680), .o(t_7701), .co(t_7702), .cout(t_7703));
compressor_4_2 u2_2642(.a(t_2648), .b(t_2645), .c(t_2642), .d(t_2639), .cin(t_7683), .o(t_7704), .co(t_7705), .cout(t_7706));
compressor_4_2 u2_2643(.a(t_2660), .b(t_2657), .c(t_2654), .d(t_2651), .cin(t_7686), .o(t_7707), .co(t_7708), .cout(t_7709));
compressor_4_2 u2_2644(.a(t_2670), .b(t_2669), .c(t_2666), .d(t_2663), .cin(t_7689), .o(t_7710), .co(t_7711), .cout(t_7712));
compressor_4_2 u2_2645(.a(t_2682), .b(t_2679), .c(t_2676), .d(t_2673), .cin(t_7692), .o(t_7713), .co(t_7714), .cout(t_7715));
compressor_4_2 u2_2646(.a(t_2694), .b(t_2691), .c(t_2688), .d(t_2685), .cin(t_7695), .o(t_7716), .co(t_7717), .cout(t_7718));
compressor_4_2 u2_2647(.a(t_2706), .b(t_2703), .c(t_2700), .d(t_2697), .cin(t_7698), .o(t_7719), .co(t_7720), .cout(t_7721));
half_adder u0_2648(.a(t_2712), .b(t_2709), .o(t_7722), .cout(t_7723));
compressor_4_2 u2_2649(.a(t_2680), .b(t_2677), .c(t_2674), .d(t_2671), .cin(t_7703), .o(t_7724), .co(t_7725), .cout(t_7726));
compressor_4_2 u2_2650(.a(t_2692), .b(t_2689), .c(t_2686), .d(t_2683), .cin(t_7706), .o(t_7727), .co(t_7728), .cout(t_7729));
compressor_4_2 u2_2651(.a(t_2704), .b(t_2701), .c(t_2698), .d(t_2695), .cin(t_7709), .o(t_7730), .co(t_7731), .cout(t_7732));
compressor_4_2 u2_2652(.a(t_2715), .b(t_2713), .c(t_2710), .d(t_2707), .cin(t_7712), .o(t_7733), .co(t_7734), .cout(t_7735));
compressor_4_2 u2_2653(.a(t_2727), .b(t_2724), .c(t_2721), .d(t_2718), .cin(t_7715), .o(t_7736), .co(t_7737), .cout(t_7738));
compressor_4_2 u2_2654(.a(t_2739), .b(t_2736), .c(t_2733), .d(t_2730), .cin(t_7718), .o(t_7739), .co(t_7740), .cout(t_7741));
compressor_4_2 u2_2655(.a(t_2751), .b(t_2748), .c(t_2745), .d(t_2742), .cin(t_7721), .o(t_7742), .co(t_7743), .cout(t_7744));
half_adder u0_2656(.a(t_2757), .b(t_2754), .o(t_7745), .cout(t_7746));
compressor_4_2 u2_2657(.a(t_2725), .b(t_2722), .c(t_2719), .d(t_2716), .cin(t_7726), .o(t_7747), .co(t_7748), .cout(t_7749));
compressor_4_2 u2_2658(.a(t_2737), .b(t_2734), .c(t_2731), .d(t_2728), .cin(t_7729), .o(t_7750), .co(t_7751), .cout(t_7752));
compressor_4_2 u2_2659(.a(t_2749), .b(t_2746), .c(t_2743), .d(t_2740), .cin(t_7732), .o(t_7753), .co(t_7754), .cout(t_7755));
compressor_4_2 u2_2660(.a(t_2760), .b(t_2758), .c(t_2755), .d(t_2752), .cin(t_7735), .o(t_7756), .co(t_7757), .cout(t_7758));
compressor_4_2 u2_2661(.a(t_2772), .b(t_2769), .c(t_2766), .d(t_2763), .cin(t_7738), .o(t_7759), .co(t_7760), .cout(t_7761));
compressor_4_2 u2_2662(.a(t_2784), .b(t_2781), .c(t_2778), .d(t_2775), .cin(t_7741), .o(t_7762), .co(t_7763), .cout(t_7764));
compressor_4_2 u2_2663(.a(t_2796), .b(t_2793), .c(t_2790), .d(t_2787), .cin(t_7744), .o(t_7765), .co(t_7766), .cout(t_7767));
compressor_3_2 u1_2664(.a(t_2805), .b(t_2802), .cin(t_2799), .o(t_7768), .cout(t_7769));
compressor_4_2 u2_2665(.a(t_2767), .b(t_2764), .c(t_2761), .d(s_121_60), .cin(t_7749), .o(t_7770), .co(t_7771), .cout(t_7772));
compressor_4_2 u2_2666(.a(t_2779), .b(t_2776), .c(t_2773), .d(t_2770), .cin(t_7752), .o(t_7773), .co(t_7774), .cout(t_7775));
compressor_4_2 u2_2667(.a(t_2791), .b(t_2788), .c(t_2785), .d(t_2782), .cin(t_7755), .o(t_7776), .co(t_7777), .cout(t_7778));
compressor_4_2 u2_2668(.a(t_2803), .b(t_2800), .c(t_2797), .d(t_2794), .cin(t_7758), .o(t_7779), .co(t_7780), .cout(t_7781));
compressor_4_2 u2_2669(.a(t_2813), .b(t_2810), .c(t_2807), .d(t_2806), .cin(t_7761), .o(t_7782), .co(t_7783), .cout(t_7784));
compressor_4_2 u2_2670(.a(t_2825), .b(t_2822), .c(t_2819), .d(t_2816), .cin(t_7764), .o(t_7785), .co(t_7786), .cout(t_7787));
compressor_4_2 u2_2671(.a(t_2837), .b(t_2834), .c(t_2831), .d(t_2828), .cin(t_7767), .o(t_7788), .co(t_7789), .cout(t_7790));
compressor_3_2 u1_2672(.a(t_2846), .b(t_2843), .cin(t_2840), .o(t_7791), .cout(t_7792));
compressor_4_2 u2_2673(.a(t_2817), .b(t_2814), .c(t_2811), .d(t_2808), .cin(t_7772), .o(t_7793), .co(t_7794), .cout(t_7795));
compressor_4_2 u2_2674(.a(t_2829), .b(t_2826), .c(t_2823), .d(t_2820), .cin(t_7775), .o(t_7796), .co(t_7797), .cout(t_7798));
compressor_4_2 u2_2675(.a(t_2841), .b(t_2838), .c(t_2835), .d(t_2832), .cin(t_7778), .o(t_7799), .co(t_7800), .cout(t_7801));
compressor_4_2 u2_2676(.a(t_2852), .b(t_2850), .c(t_2847), .d(t_2844), .cin(t_7781), .o(t_7802), .co(t_7803), .cout(t_7804));
compressor_4_2 u2_2677(.a(t_2864), .b(t_2861), .c(t_2858), .d(t_2855), .cin(t_7784), .o(t_7805), .co(t_7806), .cout(t_7807));
compressor_4_2 u2_2678(.a(t_2876), .b(t_2873), .c(t_2870), .d(t_2867), .cin(t_7787), .o(t_7808), .co(t_7809), .cout(t_7810));
compressor_4_2 u2_2679(.a(t_2888), .b(t_2885), .c(t_2882), .d(t_2879), .cin(t_7790), .o(t_7811), .co(t_7812), .cout(t_7813));
compressor_3_2 u1_2680(.a(t_2897), .b(t_2894), .cin(t_2891), .o(t_7814), .cout(t_7815));
compressor_4_2 u2_2681(.a(t_2862), .b(t_2859), .c(t_2856), .d(t_2853), .cin(t_7795), .o(t_7816), .co(t_7817), .cout(t_7818));
compressor_4_2 u2_2682(.a(t_2874), .b(t_2871), .c(t_2868), .d(t_2865), .cin(t_7798), .o(t_7819), .co(t_7820), .cout(t_7821));
compressor_4_2 u2_2683(.a(t_2886), .b(t_2883), .c(t_2880), .d(t_2877), .cin(t_7801), .o(t_7822), .co(t_7823), .cout(t_7824));
compressor_4_2 u2_2684(.a(t_2898), .b(t_2895), .c(t_2892), .d(t_2889), .cin(t_7804), .o(t_7825), .co(t_7826), .cout(t_7827));
compressor_4_2 u2_2685(.a(t_2908), .b(t_2905), .c(t_2902), .d(t_2899), .cin(t_7807), .o(t_7828), .co(t_7829), .cout(t_7830));
compressor_4_2 u2_2686(.a(t_2920), .b(t_2917), .c(t_2914), .d(t_2911), .cin(t_7810), .o(t_7831), .co(t_7832), .cout(t_7833));
compressor_4_2 u2_2687(.a(t_2932), .b(t_2929), .c(t_2926), .d(t_2923), .cin(t_7813), .o(t_7834), .co(t_7835), .cout(t_7836));
compressor_3_2 u1_2688(.a(t_2941), .b(t_2938), .cin(t_2935), .o(t_7837), .cout(t_7838));
compressor_4_2 u2_2689(.a(t_2906), .b(t_2903), .c(t_2900), .d(s_124_63), .cin(t_7818), .o(t_7839), .co(t_7840), .cout(t_7841));
compressor_4_2 u2_2690(.a(t_2918), .b(t_2915), .c(t_2912), .d(t_2909), .cin(t_7821), .o(t_7842), .co(t_7843), .cout(t_7844));
compressor_4_2 u2_2691(.a(t_2930), .b(t_2927), .c(t_2924), .d(t_2921), .cin(t_7824), .o(t_7845), .co(t_7846), .cout(t_7847));
compressor_4_2 u2_2692(.a(t_2942), .b(t_2939), .c(t_2936), .d(t_2933), .cin(t_7827), .o(t_7848), .co(t_7849), .cout(t_7850));
compressor_4_2 u2_2693(.a(t_2952), .b(t_2949), .c(t_2946), .d(t_2945), .cin(t_7830), .o(t_7851), .co(t_7852), .cout(t_7853));
compressor_4_2 u2_2694(.a(t_2964), .b(t_2961), .c(t_2958), .d(t_2955), .cin(t_7833), .o(t_7854), .co(t_7855), .cout(t_7856));
compressor_4_2 u2_2695(.a(t_2976), .b(t_2973), .c(t_2970), .d(t_2967), .cin(t_7836), .o(t_7857), .co(t_7858), .cout(t_7859));
compressor_4_2 u2_2696(.a(t_2991), .b(t_2988), .c(t_2985), .d(t_2982), .cin(t_2979), .o(t_7860), .co(t_7861), .cout(t_7862));
compressor_4_2 u2_2697(.a(t_2956), .b(t_2953), .c(t_2950), .d(t_2947), .cin(t_7841), .o(t_7863), .co(t_7864), .cout(t_7865));
compressor_4_2 u2_2698(.a(t_2968), .b(t_2965), .c(t_2962), .d(t_2959), .cin(t_7844), .o(t_7866), .co(t_7867), .cout(t_7868));
compressor_4_2 u2_2699(.a(t_2980), .b(t_2977), .c(t_2974), .d(t_2971), .cin(t_7847), .o(t_7869), .co(t_7870), .cout(t_7871));
compressor_4_2 u2_2700(.a(t_2992), .b(t_2989), .c(t_2986), .d(t_2983), .cin(t_7850), .o(t_7872), .co(t_7873), .cout(t_7874));
compressor_4_2 u2_2701(.a(t_3002), .b(t_2999), .c(t_2996), .d(t_2993), .cin(t_7853), .o(t_7875), .co(t_7876), .cout(t_7877));
compressor_4_2 u2_2702(.a(t_3014), .b(t_3011), .c(t_3008), .d(t_3005), .cin(t_7856), .o(t_7878), .co(t_7879), .cout(t_7880));
compressor_4_2 u2_2703(.a(t_3026), .b(t_3023), .c(t_3020), .d(t_3017), .cin(t_7859), .o(t_7881), .co(t_7882), .cout(t_7883));
compressor_4_2 u2_2704(.a(t_3038), .b(t_3035), .c(t_3032), .d(t_3029), .cin(t_7862), .o(t_7884), .co(t_7885), .cout(t_7886));
compressor_4_2 u2_2705(.a(t_3003), .b(t_3000), .c(t_2997), .d(t_2994), .cin(t_7865), .o(t_7887), .co(t_7888), .cout(t_7889));
compressor_4_2 u2_2706(.a(t_3015), .b(t_3012), .c(t_3009), .d(t_3006), .cin(t_7868), .o(t_7890), .co(t_7891), .cout(t_7892));
compressor_4_2 u2_2707(.a(t_3027), .b(t_3024), .c(t_3021), .d(t_3018), .cin(t_7871), .o(t_7893), .co(t_7894), .cout(t_7895));
compressor_4_2 u2_2708(.a(t_3039), .b(t_3036), .c(t_3033), .d(t_3030), .cin(t_7874), .o(t_7896), .co(t_7897), .cout(t_7898));
compressor_4_2 u2_2709(.a(t_3049), .b(t_3046), .c(t_3043), .d(t_3040), .cin(t_7877), .o(t_7899), .co(t_7900), .cout(t_7901));
compressor_4_2 u2_2710(.a(t_3061), .b(t_3058), .c(t_3055), .d(t_3052), .cin(t_7880), .o(t_7902), .co(t_7903), .cout(t_7904));
compressor_4_2 u2_2711(.a(t_3073), .b(t_3070), .c(t_3067), .d(t_3064), .cin(t_7883), .o(t_7905), .co(t_7906), .cout(t_7907));
compressor_4_2 u2_2712(.a(t_3085), .b(t_3082), .c(t_3079), .d(t_3076), .cin(t_7886), .o(t_7908), .co(t_7909), .cout(t_7910));
compressor_4_2 u2_2713(.a(t_3050), .b(t_3047), .c(t_3044), .d(t_3041), .cin(t_7889), .o(t_7911), .co(t_7912), .cout(t_7913));
compressor_4_2 u2_2714(.a(t_3062), .b(t_3059), .c(t_3056), .d(t_3053), .cin(t_7892), .o(t_7914), .co(t_7915), .cout(t_7916));
compressor_4_2 u2_2715(.a(t_3074), .b(t_3071), .c(t_3068), .d(t_3065), .cin(t_7895), .o(t_7917), .co(t_7918), .cout(t_7919));
compressor_4_2 u2_2716(.a(t_3086), .b(t_3083), .c(t_3080), .d(t_3077), .cin(t_7898), .o(t_7920), .co(t_7921), .cout(t_7922));
compressor_4_2 u2_2717(.a(t_3097), .b(t_3094), .c(t_3091), .d(t_3088), .cin(t_7901), .o(t_7923), .co(t_7924), .cout(t_7925));
compressor_4_2 u2_2718(.a(t_3109), .b(t_3106), .c(t_3103), .d(t_3100), .cin(t_7904), .o(t_7926), .co(t_7927), .cout(t_7928));
compressor_4_2 u2_2719(.a(t_3121), .b(t_3118), .c(t_3115), .d(t_3112), .cin(t_7907), .o(t_7929), .co(t_7930), .cout(t_7931));
compressor_4_2 u2_2720(.a(t_3133), .b(t_3130), .c(t_3127), .d(t_3124), .cin(t_7910), .o(t_7932), .co(t_7933), .cout(t_7934));
compressor_4_2 u2_2721(.a(t_3095), .b(t_3092), .c(t_3089), .d(s_128_64), .cin(t_7913), .o(t_7935), .co(t_7936), .cout(t_7937));
compressor_4_2 u2_2722(.a(t_3107), .b(t_3104), .c(t_3101), .d(t_3098), .cin(t_7916), .o(t_7938), .co(t_7939), .cout(t_7940));
compressor_4_2 u2_2723(.a(t_3119), .b(t_3116), .c(t_3113), .d(t_3110), .cin(t_7919), .o(t_7941), .co(t_7942), .cout(t_7943));
compressor_4_2 u2_2724(.a(t_3131), .b(t_3128), .c(t_3125), .d(t_3122), .cin(t_7922), .o(t_7944), .co(t_7945), .cout(t_7946));
compressor_4_2 u2_2725(.a(t_3142), .b(t_3139), .c(t_3136), .d(t_3134), .cin(t_7925), .o(t_7947), .co(t_7948), .cout(t_7949));
compressor_4_2 u2_2726(.a(t_3154), .b(t_3151), .c(t_3148), .d(t_3145), .cin(t_7928), .o(t_7950), .co(t_7951), .cout(t_7952));
compressor_4_2 u2_2727(.a(t_3166), .b(t_3163), .c(t_3160), .d(t_3157), .cin(t_7931), .o(t_7953), .co(t_7954), .cout(t_7955));
compressor_4_2 u2_2728(.a(t_3178), .b(t_3175), .c(t_3172), .d(t_3169), .cin(t_7934), .o(t_7956), .co(t_7957), .cout(t_7958));
compressor_4_2 u2_2729(.a(t_3143), .b(t_3140), .c(t_3137), .d(s_129_64), .cin(t_7937), .o(t_7959), .co(t_7960), .cout(t_7961));
compressor_4_2 u2_2730(.a(t_3155), .b(t_3152), .c(t_3149), .d(t_3146), .cin(t_7940), .o(t_7962), .co(t_7963), .cout(t_7964));
compressor_4_2 u2_2731(.a(t_3167), .b(t_3164), .c(t_3161), .d(t_3158), .cin(t_7943), .o(t_7965), .co(t_7966), .cout(t_7967));
compressor_4_2 u2_2732(.a(t_3179), .b(t_3176), .c(t_3173), .d(t_3170), .cin(t_7946), .o(t_7968), .co(t_7969), .cout(t_7970));
compressor_4_2 u2_2733(.a(t_3190), .b(t_3187), .c(t_3184), .d(t_3182), .cin(t_7949), .o(t_7971), .co(t_7972), .cout(t_7973));
compressor_4_2 u2_2734(.a(t_3202), .b(t_3199), .c(t_3196), .d(t_3193), .cin(t_7952), .o(t_7974), .co(t_7975), .cout(t_7976));
compressor_4_2 u2_2735(.a(t_3214), .b(t_3211), .c(t_3208), .d(t_3205), .cin(t_7955), .o(t_7977), .co(t_7978), .cout(t_7979));
compressor_4_2 u2_2736(.a(t_3226), .b(t_3223), .c(t_3220), .d(t_3217), .cin(t_7958), .o(t_7980), .co(t_7981), .cout(t_7982));
compressor_4_2 u2_2737(.a(t_3194), .b(t_3191), .c(t_3188), .d(t_3185), .cin(t_7961), .o(t_7983), .co(t_7984), .cout(t_7985));
compressor_4_2 u2_2738(.a(t_3206), .b(t_3203), .c(t_3200), .d(t_3197), .cin(t_7964), .o(t_7986), .co(t_7987), .cout(t_7988));
compressor_4_2 u2_2739(.a(t_3218), .b(t_3215), .c(t_3212), .d(t_3209), .cin(t_7967), .o(t_7989), .co(t_7990), .cout(t_7991));
compressor_4_2 u2_2740(.a(t_3230), .b(t_3227), .c(t_3224), .d(t_3221), .cin(t_7970), .o(t_7992), .co(t_7993), .cout(t_7994));
compressor_4_2 u2_2741(.a(t_3241), .b(t_3238), .c(t_3235), .d(t_3232), .cin(t_7973), .o(t_7995), .co(t_7996), .cout(t_7997));
compressor_4_2 u2_2742(.a(t_3253), .b(t_3250), .c(t_3247), .d(t_3244), .cin(t_7976), .o(t_7998), .co(t_7999), .cout(t_8000));
compressor_4_2 u2_2743(.a(t_3265), .b(t_3262), .c(t_3259), .d(t_3256), .cin(t_7979), .o(t_8001), .co(t_8002), .cout(t_8003));
compressor_4_2 u2_2744(.a(t_3277), .b(t_3274), .c(t_3271), .d(t_3268), .cin(t_7982), .o(t_8004), .co(t_8005), .cout(t_8006));
compressor_4_2 u2_2745(.a(t_3242), .b(t_3239), .c(t_3236), .d(t_3233), .cin(t_7985), .o(t_8007), .co(t_8008), .cout(t_8009));
compressor_4_2 u2_2746(.a(t_3254), .b(t_3251), .c(t_3248), .d(t_3245), .cin(t_7988), .o(t_8010), .co(t_8011), .cout(t_8012));
compressor_4_2 u2_2747(.a(t_3266), .b(t_3263), .c(t_3260), .d(t_3257), .cin(t_7991), .o(t_8013), .co(t_8014), .cout(t_8015));
compressor_4_2 u2_2748(.a(t_3278), .b(t_3275), .c(t_3272), .d(t_3269), .cin(t_7994), .o(t_8016), .co(t_8017), .cout(t_8018));
compressor_4_2 u2_2749(.a(t_3289), .b(t_3286), .c(t_3283), .d(t_3280), .cin(t_7997), .o(t_8019), .co(t_8020), .cout(t_8021));
compressor_4_2 u2_2750(.a(t_3301), .b(t_3298), .c(t_3295), .d(t_3292), .cin(t_8000), .o(t_8022), .co(t_8023), .cout(t_8024));
compressor_4_2 u2_2751(.a(t_3313), .b(t_3310), .c(t_3307), .d(t_3304), .cin(t_8003), .o(t_8025), .co(t_8026), .cout(t_8027));
compressor_4_2 u2_2752(.a(t_3325), .b(t_3322), .c(t_3319), .d(t_3316), .cin(t_8006), .o(t_8028), .co(t_8029), .cout(t_8030));
compressor_4_2 u2_2753(.a(t_3287), .b(t_3284), .c(t_3281), .d(s_132_62), .cin(t_8009), .o(t_8031), .co(t_8032), .cout(t_8033));
compressor_4_2 u2_2754(.a(t_3299), .b(t_3296), .c(t_3293), .d(t_3290), .cin(t_8012), .o(t_8034), .co(t_8035), .cout(t_8036));
compressor_4_2 u2_2755(.a(t_3311), .b(t_3308), .c(t_3305), .d(t_3302), .cin(t_8015), .o(t_8037), .co(t_8038), .cout(t_8039));
compressor_4_2 u2_2756(.a(t_3323), .b(t_3320), .c(t_3317), .d(t_3314), .cin(t_8018), .o(t_8040), .co(t_8041), .cout(t_8042));
compressor_4_2 u2_2757(.a(t_3334), .b(t_3331), .c(t_3328), .d(t_3326), .cin(t_8021), .o(t_8043), .co(t_8044), .cout(t_8045));
compressor_4_2 u2_2758(.a(t_3346), .b(t_3343), .c(t_3340), .d(t_3337), .cin(t_8024), .o(t_8046), .co(t_8047), .cout(t_8048));
compressor_4_2 u2_2759(.a(t_3358), .b(t_3355), .c(t_3352), .d(t_3349), .cin(t_8027), .o(t_8049), .co(t_8050), .cout(t_8051));
compressor_4_2 u2_2760(.a(t_3370), .b(t_3367), .c(t_3364), .d(t_3361), .cin(t_8030), .o(t_8052), .co(t_8053), .cout(t_8054));
compressor_4_2 u2_2761(.a(t_3338), .b(t_3335), .c(t_3332), .d(t_3329), .cin(t_8033), .o(t_8055), .co(t_8056), .cout(t_8057));
compressor_4_2 u2_2762(.a(t_3350), .b(t_3347), .c(t_3344), .d(t_3341), .cin(t_8036), .o(t_8058), .co(t_8059), .cout(t_8060));
compressor_4_2 u2_2763(.a(t_3362), .b(t_3359), .c(t_3356), .d(t_3353), .cin(t_8039), .o(t_8061), .co(t_8062), .cout(t_8063));
compressor_4_2 u2_2764(.a(t_3374), .b(t_3371), .c(t_3368), .d(t_3365), .cin(t_8042), .o(t_8064), .co(t_8065), .cout(t_8066));
compressor_4_2 u2_2765(.a(t_3384), .b(t_3381), .c(t_3378), .d(t_3375), .cin(t_8045), .o(t_8067), .co(t_8068), .cout(t_8069));
compressor_4_2 u2_2766(.a(t_3396), .b(t_3393), .c(t_3390), .d(t_3387), .cin(t_8048), .o(t_8070), .co(t_8071), .cout(t_8072));
compressor_4_2 u2_2767(.a(t_3408), .b(t_3405), .c(t_3402), .d(t_3399), .cin(t_8051), .o(t_8073), .co(t_8074), .cout(t_8075));
compressor_4_2 u2_2768(.a(t_3420), .b(t_3417), .c(t_3414), .d(t_3411), .cin(t_8054), .o(t_8076), .co(t_8077), .cout(t_8078));
compressor_4_2 u2_2769(.a(t_3385), .b(t_3382), .c(t_3379), .d(t_3376), .cin(t_8057), .o(t_8079), .co(t_8080), .cout(t_8081));
compressor_4_2 u2_2770(.a(t_3397), .b(t_3394), .c(t_3391), .d(t_3388), .cin(t_8060), .o(t_8082), .co(t_8083), .cout(t_8084));
compressor_4_2 u2_2771(.a(t_3409), .b(t_3406), .c(t_3403), .d(t_3400), .cin(t_8063), .o(t_8085), .co(t_8086), .cout(t_8087));
compressor_4_2 u2_2772(.a(t_3421), .b(t_3418), .c(t_3415), .d(t_3412), .cin(t_8066), .o(t_8088), .co(t_8089), .cout(t_8090));
compressor_4_2 u2_2773(.a(t_3431), .b(t_3428), .c(t_3425), .d(t_3422), .cin(t_8069), .o(t_8091), .co(t_8092), .cout(t_8093));
compressor_4_2 u2_2774(.a(t_3443), .b(t_3440), .c(t_3437), .d(t_3434), .cin(t_8072), .o(t_8094), .co(t_8095), .cout(t_8096));
compressor_4_2 u2_2775(.a(t_3455), .b(t_3452), .c(t_3449), .d(t_3446), .cin(t_8075), .o(t_8097), .co(t_8098), .cout(t_8099));
compressor_4_2 u2_2776(.a(t_3467), .b(t_3464), .c(t_3461), .d(t_3458), .cin(t_8078), .o(t_8100), .co(t_8101), .cout(t_8102));
compressor_4_2 u2_2777(.a(t_3432), .b(t_3429), .c(t_3426), .d(t_3423), .cin(t_8081), .o(t_8103), .co(t_8104), .cout(t_8105));
compressor_4_2 u2_2778(.a(t_3444), .b(t_3441), .c(t_3438), .d(t_3435), .cin(t_8084), .o(t_8106), .co(t_8107), .cout(t_8108));
compressor_4_2 u2_2779(.a(t_3456), .b(t_3453), .c(t_3450), .d(t_3447), .cin(t_8087), .o(t_8109), .co(t_8110), .cout(t_8111));
compressor_4_2 u2_2780(.a(t_3468), .b(t_3465), .c(t_3462), .d(t_3459), .cin(t_8090), .o(t_8112), .co(t_8113), .cout(t_8114));
compressor_4_2 u2_2781(.a(t_3478), .b(t_3475), .c(t_3472), .d(t_3469), .cin(t_8093), .o(t_8115), .co(t_8116), .cout(t_8117));
compressor_4_2 u2_2782(.a(t_3490), .b(t_3487), .c(t_3484), .d(t_3481), .cin(t_8096), .o(t_8118), .co(t_8119), .cout(t_8120));
compressor_4_2 u2_2783(.a(t_3502), .b(t_3499), .c(t_3496), .d(t_3493), .cin(t_8099), .o(t_8121), .co(t_8122), .cout(t_8123));
compressor_4_2 u2_2784(.a(t_3514), .b(t_3511), .c(t_3508), .d(t_3505), .cin(t_8102), .o(t_8124), .co(t_8125), .cout(t_8126));
compressor_4_2 u2_2785(.a(t_3476), .b(t_3473), .c(t_3470), .d(s_136_60), .cin(t_8105), .o(t_8127), .co(t_8128), .cout(t_8129));
compressor_4_2 u2_2786(.a(t_3488), .b(t_3485), .c(t_3482), .d(t_3479), .cin(t_8108), .o(t_8130), .co(t_8131), .cout(t_8132));
compressor_4_2 u2_2787(.a(t_3500), .b(t_3497), .c(t_3494), .d(t_3491), .cin(t_8111), .o(t_8133), .co(t_8134), .cout(t_8135));
compressor_4_2 u2_2788(.a(t_3512), .b(t_3509), .c(t_3506), .d(t_3503), .cin(t_8114), .o(t_8136), .co(t_8137), .cout(t_8138));
compressor_4_2 u2_2789(.a(t_3522), .b(t_3519), .c(t_3516), .d(t_3515), .cin(t_8117), .o(t_8139), .co(t_8140), .cout(t_8141));
compressor_4_2 u2_2790(.a(t_3534), .b(t_3531), .c(t_3528), .d(t_3525), .cin(t_8120), .o(t_8142), .co(t_8143), .cout(t_8144));
compressor_4_2 u2_2791(.a(t_3546), .b(t_3543), .c(t_3540), .d(t_3537), .cin(t_8123), .o(t_8145), .co(t_8146), .cout(t_8147));
compressor_4_2 u2_2792(.a(t_3558), .b(t_3555), .c(t_3552), .d(t_3549), .cin(t_8126), .o(t_8148), .co(t_8149), .cout(t_8150));
compressor_4_2 u2_2793(.a(t_3523), .b(t_3520), .c(t_3517), .d(s_137_60), .cin(t_8129), .o(t_8151), .co(t_8152), .cout(t_8153));
compressor_4_2 u2_2794(.a(t_3535), .b(t_3532), .c(t_3529), .d(t_3526), .cin(t_8132), .o(t_8154), .co(t_8155), .cout(t_8156));
compressor_4_2 u2_2795(.a(t_3547), .b(t_3544), .c(t_3541), .d(t_3538), .cin(t_8135), .o(t_8157), .co(t_8158), .cout(t_8159));
compressor_4_2 u2_2796(.a(t_3559), .b(t_3556), .c(t_3553), .d(t_3550), .cin(t_8138), .o(t_8160), .co(t_8161), .cout(t_8162));
compressor_4_2 u2_2797(.a(t_3570), .b(t_3567), .c(t_3564), .d(t_3561), .cin(t_8141), .o(t_8163), .co(t_8164), .cout(t_8165));
compressor_4_2 u2_2798(.a(t_3582), .b(t_3579), .c(t_3576), .d(t_3573), .cin(t_8144), .o(t_8166), .co(t_8167), .cout(t_8168));
compressor_4_2 u2_2799(.a(t_3594), .b(t_3591), .c(t_3588), .d(t_3585), .cin(t_8147), .o(t_8169), .co(t_8170), .cout(t_8171));
compressor_3_2 u1_2800(.a(t_3600), .b(t_3597), .cin(t_8150), .o(t_8172), .cout(t_8173));
compressor_4_2 u2_2801(.a(t_3571), .b(t_3568), .c(t_3565), .d(t_3562), .cin(t_8153), .o(t_8174), .co(t_8175), .cout(t_8176));
compressor_4_2 u2_2802(.a(t_3583), .b(t_3580), .c(t_3577), .d(t_3574), .cin(t_8156), .o(t_8177), .co(t_8178), .cout(t_8179));
compressor_4_2 u2_2803(.a(t_3595), .b(t_3592), .c(t_3589), .d(t_3586), .cin(t_8159), .o(t_8180), .co(t_8181), .cout(t_8182));
compressor_4_2 u2_2804(.a(t_3606), .b(t_3604), .c(t_3601), .d(t_3598), .cin(t_8162), .o(t_8183), .co(t_8184), .cout(t_8185));
compressor_4_2 u2_2805(.a(t_3618), .b(t_3615), .c(t_3612), .d(t_3609), .cin(t_8165), .o(t_8186), .co(t_8187), .cout(t_8188));
compressor_4_2 u2_2806(.a(t_3630), .b(t_3627), .c(t_3624), .d(t_3621), .cin(t_8168), .o(t_8189), .co(t_8190), .cout(t_8191));
compressor_4_2 u2_2807(.a(t_3642), .b(t_3639), .c(t_3636), .d(t_3633), .cin(t_8171), .o(t_8192), .co(t_8193), .cout(t_8194));
half_adder u0_2808(.a(t_3648), .b(t_3645), .o(t_8195), .cout(t_8196));
compressor_4_2 u2_2809(.a(t_3616), .b(t_3613), .c(t_3610), .d(t_3607), .cin(t_8176), .o(t_8197), .co(t_8198), .cout(t_8199));
compressor_4_2 u2_2810(.a(t_3628), .b(t_3625), .c(t_3622), .d(t_3619), .cin(t_8179), .o(t_8200), .co(t_8201), .cout(t_8202));
compressor_4_2 u2_2811(.a(t_3640), .b(t_3637), .c(t_3634), .d(t_3631), .cin(t_8182), .o(t_8203), .co(t_8204), .cout(t_8205));
compressor_4_2 u2_2812(.a(t_3651), .b(t_3649), .c(t_3646), .d(t_3643), .cin(t_8185), .o(t_8206), .co(t_8207), .cout(t_8208));
compressor_4_2 u2_2813(.a(t_3663), .b(t_3660), .c(t_3657), .d(t_3654), .cin(t_8188), .o(t_8209), .co(t_8210), .cout(t_8211));
compressor_4_2 u2_2814(.a(t_3675), .b(t_3672), .c(t_3669), .d(t_3666), .cin(t_8191), .o(t_8212), .co(t_8213), .cout(t_8214));
compressor_4_2 u2_2815(.a(t_3687), .b(t_3684), .c(t_3681), .d(t_3678), .cin(t_8194), .o(t_8215), .co(t_8216), .cout(t_8217));
half_adder u0_2816(.a(t_3693), .b(t_3690), .o(t_8218), .cout(t_8219));
compressor_4_2 u2_2817(.a(t_3658), .b(t_3655), .c(t_3652), .d(s_140_58), .cin(t_8199), .o(t_8220), .co(t_8221), .cout(t_8222));
compressor_4_2 u2_2818(.a(t_3670), .b(t_3667), .c(t_3664), .d(t_3661), .cin(t_8202), .o(t_8223), .co(t_8224), .cout(t_8225));
compressor_4_2 u2_2819(.a(t_3682), .b(t_3679), .c(t_3676), .d(t_3673), .cin(t_8205), .o(t_8226), .co(t_8227), .cout(t_8228));
compressor_4_2 u2_2820(.a(t_3694), .b(t_3691), .c(t_3688), .d(t_3685), .cin(t_8208), .o(t_8229), .co(t_8230), .cout(t_8231));
compressor_4_2 u2_2821(.a(t_3705), .b(t_3702), .c(t_3699), .d(t_3696), .cin(t_8211), .o(t_8232), .co(t_8233), .cout(t_8234));
compressor_4_2 u2_2822(.a(t_3717), .b(t_3714), .c(t_3711), .d(t_3708), .cin(t_8214), .o(t_8235), .co(t_8236), .cout(t_8237));
compressor_4_2 u2_2823(.a(t_3729), .b(t_3726), .c(t_3723), .d(t_3720), .cin(t_8217), .o(t_8238), .co(t_8239), .cout(t_8240));
compressor_3_2 u1_2824(.a(t_3738), .b(t_3735), .cin(t_3732), .o(t_8241), .cout(t_8242));
compressor_4_2 u2_2825(.a(t_3706), .b(t_3703), .c(t_3700), .d(t_3697), .cin(t_8222), .o(t_8243), .co(t_8244), .cout(t_8245));
compressor_4_2 u2_2826(.a(t_3718), .b(t_3715), .c(t_3712), .d(t_3709), .cin(t_8225), .o(t_8246), .co(t_8247), .cout(t_8248));
compressor_4_2 u2_2827(.a(t_3730), .b(t_3727), .c(t_3724), .d(t_3721), .cin(t_8228), .o(t_8249), .co(t_8250), .cout(t_8251));
compressor_4_2 u2_2828(.a(t_3740), .b(t_3739), .c(t_3736), .d(t_3733), .cin(t_8231), .o(t_8252), .co(t_8253), .cout(t_8254));
compressor_4_2 u2_2829(.a(t_3752), .b(t_3749), .c(t_3746), .d(t_3743), .cin(t_8234), .o(t_8255), .co(t_8256), .cout(t_8257));
compressor_4_2 u2_2830(.a(t_3764), .b(t_3761), .c(t_3758), .d(t_3755), .cin(t_8237), .o(t_8258), .co(t_8259), .cout(t_8260));
compressor_4_2 u2_2831(.a(t_3776), .b(t_3773), .c(t_3770), .d(t_3767), .cin(t_8240), .o(t_8261), .co(t_8262), .cout(t_8263));
half_adder u0_2832(.a(t_3782), .b(t_3779), .o(t_8264), .cout(t_8265));
compressor_4_2 u2_2833(.a(t_3750), .b(t_3747), .c(t_3744), .d(t_3741), .cin(t_8245), .o(t_8266), .co(t_8267), .cout(t_8268));
compressor_4_2 u2_2834(.a(t_3762), .b(t_3759), .c(t_3756), .d(t_3753), .cin(t_8248), .o(t_8269), .co(t_8270), .cout(t_8271));
compressor_4_2 u2_2835(.a(t_3774), .b(t_3771), .c(t_3768), .d(t_3765), .cin(t_8251), .o(t_8272), .co(t_8273), .cout(t_8274));
compressor_4_2 u2_2836(.a(t_3784), .b(t_3783), .c(t_3780), .d(t_3777), .cin(t_8254), .o(t_8275), .co(t_8276), .cout(t_8277));
compressor_4_2 u2_2837(.a(t_3796), .b(t_3793), .c(t_3790), .d(t_3787), .cin(t_8257), .o(t_8278), .co(t_8279), .cout(t_8280));
compressor_4_2 u2_2838(.a(t_3808), .b(t_3805), .c(t_3802), .d(t_3799), .cin(t_8260), .o(t_8281), .co(t_8282), .cout(t_8283));
compressor_4_2 u2_2839(.a(t_3820), .b(t_3817), .c(t_3814), .d(t_3811), .cin(t_8263), .o(t_8284), .co(t_8285), .cout(t_8286));
half_adder u0_2840(.a(t_3826), .b(t_3823), .o(t_8287), .cout(t_8288));
compressor_4_2 u2_2841(.a(t_3794), .b(t_3791), .c(t_3788), .d(t_3785), .cin(t_8268), .o(t_8289), .co(t_8290), .cout(t_8291));
compressor_4_2 u2_2842(.a(t_3806), .b(t_3803), .c(t_3800), .d(t_3797), .cin(t_8271), .o(t_8292), .co(t_8293), .cout(t_8294));
compressor_4_2 u2_2843(.a(t_3818), .b(t_3815), .c(t_3812), .d(t_3809), .cin(t_8274), .o(t_8295), .co(t_8296), .cout(t_8297));
compressor_4_2 u2_2844(.a(t_3828), .b(t_3827), .c(t_3824), .d(t_3821), .cin(t_8277), .o(t_8298), .co(t_8299), .cout(t_8300));
compressor_4_2 u2_2845(.a(t_3840), .b(t_3837), .c(t_3834), .d(t_3831), .cin(t_8280), .o(t_8301), .co(t_8302), .cout(t_8303));
compressor_4_2 u2_2846(.a(t_3852), .b(t_3849), .c(t_3846), .d(t_3843), .cin(t_8283), .o(t_8304), .co(t_8305), .cout(t_8306));
compressor_4_2 u2_2847(.a(t_3864), .b(t_3861), .c(t_3858), .d(t_3855), .cin(t_8286), .o(t_8307), .co(t_8308), .cout(t_8309));
half_adder u0_2848(.a(t_3870), .b(t_3867), .o(t_8310), .cout(t_8311));
compressor_4_2 u2_2849(.a(t_3835), .b(t_3832), .c(t_3829), .d(s_144_56), .cin(t_8291), .o(t_8312), .co(t_8313), .cout(t_8314));
compressor_4_2 u2_2850(.a(t_3847), .b(t_3844), .c(t_3841), .d(t_3838), .cin(t_8294), .o(t_8315), .co(t_8316), .cout(t_8317));
compressor_4_2 u2_2851(.a(t_3859), .b(t_3856), .c(t_3853), .d(t_3850), .cin(t_8297), .o(t_8318), .co(t_8319), .cout(t_8320));
compressor_4_2 u2_2852(.a(t_3871), .b(t_3868), .c(t_3865), .d(t_3862), .cin(t_8300), .o(t_8321), .co(t_8322), .cout(t_8323));
compressor_4_2 u2_2853(.a(t_3881), .b(t_3878), .c(t_3875), .d(t_3872), .cin(t_8303), .o(t_8324), .co(t_8325), .cout(t_8326));
compressor_4_2 u2_2854(.a(t_3893), .b(t_3890), .c(t_3887), .d(t_3884), .cin(t_8306), .o(t_8327), .co(t_8328), .cout(t_8329));
compressor_4_2 u2_2855(.a(t_3905), .b(t_3902), .c(t_3899), .d(t_3896), .cin(t_8309), .o(t_8330), .co(t_8331), .cout(t_8332));
half_adder u0_2856(.a(t_3911), .b(t_3908), .o(t_8333), .cout(t_8334));
compressor_4_2 u2_2857(.a(t_3879), .b(t_3876), .c(t_3873), .d(s_145_56), .cin(t_8314), .o(t_8335), .co(t_8336), .cout(t_8337));
compressor_4_2 u2_2858(.a(t_3891), .b(t_3888), .c(t_3885), .d(t_3882), .cin(t_8317), .o(t_8338), .co(t_8339), .cout(t_8340));
compressor_4_2 u2_2859(.a(t_3903), .b(t_3900), .c(t_3897), .d(t_3894), .cin(t_8320), .o(t_8341), .co(t_8342), .cout(t_8343));
compressor_4_2 u2_2860(.a(t_3914), .b(t_3912), .c(t_3909), .d(t_3906), .cin(t_8323), .o(t_8344), .co(t_8345), .cout(t_8346));
compressor_4_2 u2_2861(.a(t_3926), .b(t_3923), .c(t_3920), .d(t_3917), .cin(t_8326), .o(t_8347), .co(t_8348), .cout(t_8349));
compressor_4_2 u2_2862(.a(t_3938), .b(t_3935), .c(t_3932), .d(t_3929), .cin(t_8329), .o(t_8350), .co(t_8351), .cout(t_8352));
compressor_4_2 u2_2863(.a(t_3950), .b(t_3947), .c(t_3944), .d(t_3941), .cin(t_8332), .o(t_8353), .co(t_8354), .cout(t_8355));
compressor_4_2 u2_2864(.a(t_3924), .b(t_3921), .c(t_3918), .d(t_3915), .cin(t_8337), .o(t_8356), .co(t_8357), .cout(t_8358));
compressor_4_2 u2_2865(.a(t_3936), .b(t_3933), .c(t_3930), .d(t_3927), .cin(t_8340), .o(t_8359), .co(t_8360), .cout(t_8361));
compressor_4_2 u2_2866(.a(t_3948), .b(t_3945), .c(t_3942), .d(t_3939), .cin(t_8343), .o(t_8362), .co(t_8363), .cout(t_8364));
compressor_4_2 u2_2867(.a(t_3959), .b(t_3956), .c(t_3954), .d(t_3951), .cin(t_8346), .o(t_8365), .co(t_8366), .cout(t_8367));
compressor_4_2 u2_2868(.a(t_3971), .b(t_3968), .c(t_3965), .d(t_3962), .cin(t_8349), .o(t_8368), .co(t_8369), .cout(t_8370));
compressor_4_2 u2_2869(.a(t_3983), .b(t_3980), .c(t_3977), .d(t_3974), .cin(t_8352), .o(t_8371), .co(t_8372), .cout(t_8373));
compressor_4_2 u2_2870(.a(t_3995), .b(t_3992), .c(t_3989), .d(t_3986), .cin(t_8355), .o(t_8374), .co(t_8375), .cout(t_8376));
compressor_4_2 u2_2871(.a(t_3966), .b(t_3963), .c(t_3960), .d(t_3957), .cin(t_8358), .o(t_8377), .co(t_8378), .cout(t_8379));
compressor_4_2 u2_2872(.a(t_3978), .b(t_3975), .c(t_3972), .d(t_3969), .cin(t_8361), .o(t_8380), .co(t_8381), .cout(t_8382));
compressor_4_2 u2_2873(.a(t_3990), .b(t_3987), .c(t_3984), .d(t_3981), .cin(t_8364), .o(t_8383), .co(t_8384), .cout(t_8385));
compressor_4_2 u2_2874(.a(t_4001), .b(t_3998), .c(t_3996), .d(t_3993), .cin(t_8367), .o(t_8386), .co(t_8387), .cout(t_8388));
compressor_4_2 u2_2875(.a(t_4013), .b(t_4010), .c(t_4007), .d(t_4004), .cin(t_8370), .o(t_8389), .co(t_8390), .cout(t_8391));
compressor_4_2 u2_2876(.a(t_4025), .b(t_4022), .c(t_4019), .d(t_4016), .cin(t_8373), .o(t_8392), .co(t_8393), .cout(t_8394));
compressor_4_2 u2_2877(.a(t_4037), .b(t_4034), .c(t_4031), .d(t_4028), .cin(t_8376), .o(t_8395), .co(t_8396), .cout(t_8397));
compressor_4_2 u2_2878(.a(t_4005), .b(t_4002), .c(t_3999), .d(s_148_54), .cin(t_8379), .o(t_8398), .co(t_8399), .cout(t_8400));
compressor_4_2 u2_2879(.a(t_4017), .b(t_4014), .c(t_4011), .d(t_4008), .cin(t_8382), .o(t_8401), .co(t_8402), .cout(t_8403));
compressor_4_2 u2_2880(.a(t_4029), .b(t_4026), .c(t_4023), .d(t_4020), .cin(t_8385), .o(t_8404), .co(t_8405), .cout(t_8406));
compressor_4_2 u2_2881(.a(t_4040), .b(t_4038), .c(t_4035), .d(t_4032), .cin(t_8388), .o(t_8407), .co(t_8408), .cout(t_8409));
compressor_4_2 u2_2882(.a(t_4052), .b(t_4049), .c(t_4046), .d(t_4043), .cin(t_8391), .o(t_8410), .co(t_8411), .cout(t_8412));
compressor_4_2 u2_2883(.a(t_4064), .b(t_4061), .c(t_4058), .d(t_4055), .cin(t_8394), .o(t_8413), .co(t_8414), .cout(t_8415));
compressor_4_2 u2_2884(.a(t_4076), .b(t_4073), .c(t_4070), .d(t_4067), .cin(t_8397), .o(t_8416), .co(t_8417), .cout(t_8418));
compressor_4_2 u2_2885(.a(t_4050), .b(t_4047), .c(t_4044), .d(t_4041), .cin(t_8400), .o(t_8419), .co(t_8420), .cout(t_8421));
compressor_4_2 u2_2886(.a(t_4062), .b(t_4059), .c(t_4056), .d(t_4053), .cin(t_8403), .o(t_8422), .co(t_8423), .cout(t_8424));
compressor_4_2 u2_2887(.a(t_4074), .b(t_4071), .c(t_4068), .d(t_4065), .cin(t_8406), .o(t_8425), .co(t_8426), .cout(t_8427));
compressor_4_2 u2_2888(.a(t_4084), .b(t_4081), .c(t_4080), .d(t_4077), .cin(t_8409), .o(t_8428), .co(t_8429), .cout(t_8430));
compressor_4_2 u2_2889(.a(t_4096), .b(t_4093), .c(t_4090), .d(t_4087), .cin(t_8412), .o(t_8431), .co(t_8432), .cout(t_8433));
compressor_4_2 u2_2890(.a(t_4108), .b(t_4105), .c(t_4102), .d(t_4099), .cin(t_8415), .o(t_8434), .co(t_8435), .cout(t_8436));
compressor_4_2 u2_2891(.a(t_4120), .b(t_4117), .c(t_4114), .d(t_4111), .cin(t_8418), .o(t_8437), .co(t_8438), .cout(t_8439));
compressor_4_2 u2_2892(.a(t_4091), .b(t_4088), .c(t_4085), .d(t_4082), .cin(t_8421), .o(t_8440), .co(t_8441), .cout(t_8442));
compressor_4_2 u2_2893(.a(t_4103), .b(t_4100), .c(t_4097), .d(t_4094), .cin(t_8424), .o(t_8443), .co(t_8444), .cout(t_8445));
compressor_4_2 u2_2894(.a(t_4115), .b(t_4112), .c(t_4109), .d(t_4106), .cin(t_8427), .o(t_8446), .co(t_8447), .cout(t_8448));
compressor_4_2 u2_2895(.a(t_4125), .b(t_4122), .c(t_4121), .d(t_4118), .cin(t_8430), .o(t_8449), .co(t_8450), .cout(t_8451));
compressor_4_2 u2_2896(.a(t_4137), .b(t_4134), .c(t_4131), .d(t_4128), .cin(t_8433), .o(t_8452), .co(t_8453), .cout(t_8454));
compressor_4_2 u2_2897(.a(t_4149), .b(t_4146), .c(t_4143), .d(t_4140), .cin(t_8436), .o(t_8455), .co(t_8456), .cout(t_8457));
compressor_4_2 u2_2898(.a(t_4161), .b(t_4158), .c(t_4155), .d(t_4152), .cin(t_8439), .o(t_8458), .co(t_8459), .cout(t_8460));
compressor_4_2 u2_2899(.a(t_4132), .b(t_4129), .c(t_4126), .d(t_4123), .cin(t_8442), .o(t_8461), .co(t_8462), .cout(t_8463));
compressor_4_2 u2_2900(.a(t_4144), .b(t_4141), .c(t_4138), .d(t_4135), .cin(t_8445), .o(t_8464), .co(t_8465), .cout(t_8466));
compressor_4_2 u2_2901(.a(t_4156), .b(t_4153), .c(t_4150), .d(t_4147), .cin(t_8448), .o(t_8467), .co(t_8468), .cout(t_8469));
compressor_4_2 u2_2902(.a(t_4166), .b(t_4163), .c(t_4162), .d(t_4159), .cin(t_8451), .o(t_8470), .co(t_8471), .cout(t_8472));
compressor_4_2 u2_2903(.a(t_4178), .b(t_4175), .c(t_4172), .d(t_4169), .cin(t_8454), .o(t_8473), .co(t_8474), .cout(t_8475));
compressor_4_2 u2_2904(.a(t_4190), .b(t_4187), .c(t_4184), .d(t_4181), .cin(t_8457), .o(t_8476), .co(t_8477), .cout(t_8478));
compressor_4_2 u2_2905(.a(t_4202), .b(t_4199), .c(t_4196), .d(t_4193), .cin(t_8460), .o(t_8479), .co(t_8480), .cout(t_8481));
compressor_4_2 u2_2906(.a(t_4170), .b(t_4167), .c(t_4164), .d(s_152_52), .cin(t_8463), .o(t_8482), .co(t_8483), .cout(t_8484));
compressor_4_2 u2_2907(.a(t_4182), .b(t_4179), .c(t_4176), .d(t_4173), .cin(t_8466), .o(t_8485), .co(t_8486), .cout(t_8487));
compressor_4_2 u2_2908(.a(t_4194), .b(t_4191), .c(t_4188), .d(t_4185), .cin(t_8469), .o(t_8488), .co(t_8489), .cout(t_8490));
compressor_4_2 u2_2909(.a(t_4204), .b(t_4203), .c(t_4200), .d(t_4197), .cin(t_8472), .o(t_8491), .co(t_8492), .cout(t_8493));
compressor_4_2 u2_2910(.a(t_4216), .b(t_4213), .c(t_4210), .d(t_4207), .cin(t_8475), .o(t_8494), .co(t_8495), .cout(t_8496));
compressor_4_2 u2_2911(.a(t_4228), .b(t_4225), .c(t_4222), .d(t_4219), .cin(t_8478), .o(t_8497), .co(t_8498), .cout(t_8499));
compressor_4_2 u2_2912(.a(t_4240), .b(t_4237), .c(t_4234), .d(t_4231), .cin(t_8481), .o(t_8500), .co(t_8501), .cout(t_8502));
compressor_4_2 u2_2913(.a(t_4211), .b(t_4208), .c(t_4205), .d(s_153_52), .cin(t_8484), .o(t_8503), .co(t_8504), .cout(t_8505));
compressor_4_2 u2_2914(.a(t_4223), .b(t_4220), .c(t_4217), .d(t_4214), .cin(t_8487), .o(t_8506), .co(t_8507), .cout(t_8508));
compressor_4_2 u2_2915(.a(t_4235), .b(t_4232), .c(t_4229), .d(t_4226), .cin(t_8490), .o(t_8509), .co(t_8510), .cout(t_8511));
compressor_4_2 u2_2916(.a(t_4246), .b(t_4243), .c(t_4241), .d(t_4238), .cin(t_8493), .o(t_8512), .co(t_8513), .cout(t_8514));
compressor_4_2 u2_2917(.a(t_4258), .b(t_4255), .c(t_4252), .d(t_4249), .cin(t_8496), .o(t_8515), .co(t_8516), .cout(t_8517));
compressor_4_2 u2_2918(.a(t_4270), .b(t_4267), .c(t_4264), .d(t_4261), .cin(t_8499), .o(t_8518), .co(t_8519), .cout(t_8520));
compressor_3_2 u1_2919(.a(t_4276), .b(t_4273), .cin(t_8502), .o(t_8521), .cout(t_8522));
compressor_4_2 u2_2920(.a(t_4253), .b(t_4250), .c(t_4247), .d(t_4244), .cin(t_8505), .o(t_8523), .co(t_8524), .cout(t_8525));
compressor_4_2 u2_2921(.a(t_4265), .b(t_4262), .c(t_4259), .d(t_4256), .cin(t_8508), .o(t_8526), .co(t_8527), .cout(t_8528));
compressor_4_2 u2_2922(.a(t_4277), .b(t_4274), .c(t_4271), .d(t_4268), .cin(t_8511), .o(t_8529), .co(t_8530), .cout(t_8531));
compressor_4_2 u2_2923(.a(t_4288), .b(t_4285), .c(t_4282), .d(t_4280), .cin(t_8514), .o(t_8532), .co(t_8533), .cout(t_8534));
compressor_4_2 u2_2924(.a(t_4300), .b(t_4297), .c(t_4294), .d(t_4291), .cin(t_8517), .o(t_8535), .co(t_8536), .cout(t_8537));
compressor_4_2 u2_2925(.a(t_4312), .b(t_4309), .c(t_4306), .d(t_4303), .cin(t_8520), .o(t_8538), .co(t_8539), .cout(t_8540));
half_adder u0_2926(.a(t_4318), .b(t_4315), .o(t_8541), .cout(t_8542));
compressor_4_2 u2_2927(.a(t_4292), .b(t_4289), .c(t_4286), .d(t_4283), .cin(t_8525), .o(t_8543), .co(t_8544), .cout(t_8545));
compressor_4_2 u2_2928(.a(t_4304), .b(t_4301), .c(t_4298), .d(t_4295), .cin(t_8528), .o(t_8546), .co(t_8547), .cout(t_8548));
compressor_4_2 u2_2929(.a(t_4316), .b(t_4313), .c(t_4310), .d(t_4307), .cin(t_8531), .o(t_8549), .co(t_8550), .cout(t_8551));
compressor_4_2 u2_2930(.a(t_4327), .b(t_4324), .c(t_4321), .d(t_4319), .cin(t_8534), .o(t_8552), .co(t_8553), .cout(t_8554));
compressor_4_2 u2_2931(.a(t_4339), .b(t_4336), .c(t_4333), .d(t_4330), .cin(t_8537), .o(t_8555), .co(t_8556), .cout(t_8557));
compressor_4_2 u2_2932(.a(t_4351), .b(t_4348), .c(t_4345), .d(t_4342), .cin(t_8540), .o(t_8558), .co(t_8559), .cout(t_8560));
half_adder u0_2933(.a(t_4357), .b(t_4354), .o(t_8561), .cout(t_8562));
compressor_4_2 u2_2934(.a(t_4328), .b(t_4325), .c(t_4322), .d(s_156_50), .cin(t_8545), .o(t_8563), .co(t_8564), .cout(t_8565));
compressor_4_2 u2_2935(.a(t_4340), .b(t_4337), .c(t_4334), .d(t_4331), .cin(t_8548), .o(t_8566), .co(t_8567), .cout(t_8568));
compressor_4_2 u2_2936(.a(t_4352), .b(t_4349), .c(t_4346), .d(t_4343), .cin(t_8551), .o(t_8569), .co(t_8570), .cout(t_8571));
compressor_4_2 u2_2937(.a(t_4363), .b(t_4360), .c(t_4358), .d(t_4355), .cin(t_8554), .o(t_8572), .co(t_8573), .cout(t_8574));
compressor_4_2 u2_2938(.a(t_4375), .b(t_4372), .c(t_4369), .d(t_4366), .cin(t_8557), .o(t_8575), .co(t_8576), .cout(t_8577));
compressor_4_2 u2_2939(.a(t_4387), .b(t_4384), .c(t_4381), .d(t_4378), .cin(t_8560), .o(t_8578), .co(t_8579), .cout(t_8580));
compressor_3_2 u1_2940(.a(t_4396), .b(t_4393), .cin(t_4390), .o(t_8581), .cout(t_8582));
compressor_4_2 u2_2941(.a(t_4370), .b(t_4367), .c(t_4364), .d(t_4361), .cin(t_8565), .o(t_8583), .co(t_8584), .cout(t_8585));
compressor_4_2 u2_2942(.a(t_4382), .b(t_4379), .c(t_4376), .d(t_4373), .cin(t_8568), .o(t_8586), .co(t_8587), .cout(t_8588));
compressor_4_2 u2_2943(.a(t_4394), .b(t_4391), .c(t_4388), .d(t_4385), .cin(t_8571), .o(t_8589), .co(t_8590), .cout(t_8591));
compressor_4_2 u2_2944(.a(t_4404), .b(t_4401), .c(t_4398), .d(t_4397), .cin(t_8574), .o(t_8592), .co(t_8593), .cout(t_8594));
compressor_4_2 u2_2945(.a(t_4416), .b(t_4413), .c(t_4410), .d(t_4407), .cin(t_8577), .o(t_8595), .co(t_8596), .cout(t_8597));
compressor_4_2 u2_2946(.a(t_4428), .b(t_4425), .c(t_4422), .d(t_4419), .cin(t_8580), .o(t_8598), .co(t_8599), .cout(t_8600));
half_adder u0_2947(.a(t_4434), .b(t_4431), .o(t_8601), .cout(t_8602));
compressor_4_2 u2_2948(.a(t_4408), .b(t_4405), .c(t_4402), .d(t_4399), .cin(t_8585), .o(t_8603), .co(t_8604), .cout(t_8605));
compressor_4_2 u2_2949(.a(t_4420), .b(t_4417), .c(t_4414), .d(t_4411), .cin(t_8588), .o(t_8606), .co(t_8607), .cout(t_8608));
compressor_4_2 u2_2950(.a(t_4432), .b(t_4429), .c(t_4426), .d(t_4423), .cin(t_8591), .o(t_8609), .co(t_8610), .cout(t_8611));
compressor_4_2 u2_2951(.a(t_4442), .b(t_4439), .c(t_4436), .d(t_4435), .cin(t_8594), .o(t_8612), .co(t_8613), .cout(t_8614));
compressor_4_2 u2_2952(.a(t_4454), .b(t_4451), .c(t_4448), .d(t_4445), .cin(t_8597), .o(t_8615), .co(t_8616), .cout(t_8617));
compressor_4_2 u2_2953(.a(t_4466), .b(t_4463), .c(t_4460), .d(t_4457), .cin(t_8600), .o(t_8618), .co(t_8619), .cout(t_8620));
half_adder u0_2954(.a(t_4472), .b(t_4469), .o(t_8621), .cout(t_8622));
compressor_4_2 u2_2955(.a(t_4446), .b(t_4443), .c(t_4440), .d(t_4437), .cin(t_8605), .o(t_8623), .co(t_8624), .cout(t_8625));
compressor_4_2 u2_2956(.a(t_4458), .b(t_4455), .c(t_4452), .d(t_4449), .cin(t_8608), .o(t_8626), .co(t_8627), .cout(t_8628));
compressor_4_2 u2_2957(.a(t_4470), .b(t_4467), .c(t_4464), .d(t_4461), .cin(t_8611), .o(t_8629), .co(t_8630), .cout(t_8631));
compressor_4_2 u2_2958(.a(t_4480), .b(t_4477), .c(t_4474), .d(t_4473), .cin(t_8614), .o(t_8632), .co(t_8633), .cout(t_8634));
compressor_4_2 u2_2959(.a(t_4492), .b(t_4489), .c(t_4486), .d(t_4483), .cin(t_8617), .o(t_8635), .co(t_8636), .cout(t_8637));
compressor_4_2 u2_2960(.a(t_4504), .b(t_4501), .c(t_4498), .d(t_4495), .cin(t_8620), .o(t_8638), .co(t_8639), .cout(t_8640));
half_adder u0_2961(.a(t_4510), .b(t_4507), .o(t_8641), .cout(t_8642));
compressor_4_2 u2_2962(.a(t_4481), .b(t_4478), .c(t_4475), .d(s_160_48), .cin(t_8625), .o(t_8643), .co(t_8644), .cout(t_8645));
compressor_4_2 u2_2963(.a(t_4493), .b(t_4490), .c(t_4487), .d(t_4484), .cin(t_8628), .o(t_8646), .co(t_8647), .cout(t_8648));
compressor_4_2 u2_2964(.a(t_4505), .b(t_4502), .c(t_4499), .d(t_4496), .cin(t_8631), .o(t_8649), .co(t_8650), .cout(t_8651));
compressor_4_2 u2_2965(.a(t_4515), .b(t_4512), .c(t_4511), .d(t_4508), .cin(t_8634), .o(t_8652), .co(t_8653), .cout(t_8654));
compressor_4_2 u2_2966(.a(t_4527), .b(t_4524), .c(t_4521), .d(t_4518), .cin(t_8637), .o(t_8655), .co(t_8656), .cout(t_8657));
compressor_4_2 u2_2967(.a(t_4539), .b(t_4536), .c(t_4533), .d(t_4530), .cin(t_8640), .o(t_8658), .co(t_8659), .cout(t_8660));
half_adder u0_2968(.a(t_4545), .b(t_4542), .o(t_8661), .cout(t_8662));
compressor_4_2 u2_2969(.a(t_4519), .b(t_4516), .c(t_4513), .d(s_161_48), .cin(t_8645), .o(t_8663), .co(t_8664), .cout(t_8665));
compressor_4_2 u2_2970(.a(t_4531), .b(t_4528), .c(t_4525), .d(t_4522), .cin(t_8648), .o(t_8666), .co(t_8667), .cout(t_8668));
compressor_4_2 u2_2971(.a(t_4543), .b(t_4540), .c(t_4537), .d(t_4534), .cin(t_8651), .o(t_8669), .co(t_8670), .cout(t_8671));
compressor_4_2 u2_2972(.a(t_4554), .b(t_4551), .c(t_4548), .d(t_4546), .cin(t_8654), .o(t_8672), .co(t_8673), .cout(t_8674));
compressor_4_2 u2_2973(.a(t_4566), .b(t_4563), .c(t_4560), .d(t_4557), .cin(t_8657), .o(t_8675), .co(t_8676), .cout(t_8677));
compressor_4_2 u2_2974(.a(t_4578), .b(t_4575), .c(t_4572), .d(t_4569), .cin(t_8660), .o(t_8678), .co(t_8679), .cout(t_8680));
compressor_4_2 u2_2975(.a(t_4558), .b(t_4555), .c(t_4552), .d(t_4549), .cin(t_8665), .o(t_8681), .co(t_8682), .cout(t_8683));
compressor_4_2 u2_2976(.a(t_4570), .b(t_4567), .c(t_4564), .d(t_4561), .cin(t_8668), .o(t_8684), .co(t_8685), .cout(t_8686));
compressor_4_2 u2_2977(.a(t_4582), .b(t_4579), .c(t_4576), .d(t_4573), .cin(t_8671), .o(t_8687), .co(t_8688), .cout(t_8689));
compressor_4_2 u2_2978(.a(t_4593), .b(t_4590), .c(t_4587), .d(t_4584), .cin(t_8674), .o(t_8690), .co(t_8691), .cout(t_8692));
compressor_4_2 u2_2979(.a(t_4605), .b(t_4602), .c(t_4599), .d(t_4596), .cin(t_8677), .o(t_8693), .co(t_8694), .cout(t_8695));
compressor_4_2 u2_2980(.a(t_4617), .b(t_4614), .c(t_4611), .d(t_4608), .cin(t_8680), .o(t_8696), .co(t_8697), .cout(t_8698));
compressor_4_2 u2_2981(.a(t_4594), .b(t_4591), .c(t_4588), .d(t_4585), .cin(t_8683), .o(t_8699), .co(t_8700), .cout(t_8701));
compressor_4_2 u2_2982(.a(t_4606), .b(t_4603), .c(t_4600), .d(t_4597), .cin(t_8686), .o(t_8702), .co(t_8703), .cout(t_8704));
compressor_4_2 u2_2983(.a(t_4618), .b(t_4615), .c(t_4612), .d(t_4609), .cin(t_8689), .o(t_8705), .co(t_8706), .cout(t_8707));
compressor_4_2 u2_2984(.a(t_4629), .b(t_4626), .c(t_4623), .d(t_4620), .cin(t_8692), .o(t_8708), .co(t_8709), .cout(t_8710));
compressor_4_2 u2_2985(.a(t_4641), .b(t_4638), .c(t_4635), .d(t_4632), .cin(t_8695), .o(t_8711), .co(t_8712), .cout(t_8713));
compressor_4_2 u2_2986(.a(t_4653), .b(t_4650), .c(t_4647), .d(t_4644), .cin(t_8698), .o(t_8714), .co(t_8715), .cout(t_8716));
compressor_4_2 u2_2987(.a(t_4627), .b(t_4624), .c(t_4621), .d(s_164_46), .cin(t_8701), .o(t_8717), .co(t_8718), .cout(t_8719));
compressor_4_2 u2_2988(.a(t_4639), .b(t_4636), .c(t_4633), .d(t_4630), .cin(t_8704), .o(t_8720), .co(t_8721), .cout(t_8722));
compressor_4_2 u2_2989(.a(t_4651), .b(t_4648), .c(t_4645), .d(t_4642), .cin(t_8707), .o(t_8723), .co(t_8724), .cout(t_8725));
compressor_4_2 u2_2990(.a(t_4662), .b(t_4659), .c(t_4656), .d(t_4654), .cin(t_8710), .o(t_8726), .co(t_8727), .cout(t_8728));
compressor_4_2 u2_2991(.a(t_4674), .b(t_4671), .c(t_4668), .d(t_4665), .cin(t_8713), .o(t_8729), .co(t_8730), .cout(t_8731));
compressor_4_2 u2_2992(.a(t_4686), .b(t_4683), .c(t_4680), .d(t_4677), .cin(t_8716), .o(t_8732), .co(t_8733), .cout(t_8734));
compressor_4_2 u2_2993(.a(t_4666), .b(t_4663), .c(t_4660), .d(t_4657), .cin(t_8719), .o(t_8735), .co(t_8736), .cout(t_8737));
compressor_4_2 u2_2994(.a(t_4678), .b(t_4675), .c(t_4672), .d(t_4669), .cin(t_8722), .o(t_8738), .co(t_8739), .cout(t_8740));
compressor_4_2 u2_2995(.a(t_4690), .b(t_4687), .c(t_4684), .d(t_4681), .cin(t_8725), .o(t_8741), .co(t_8742), .cout(t_8743));
compressor_4_2 u2_2996(.a(t_4700), .b(t_4697), .c(t_4694), .d(t_4691), .cin(t_8728), .o(t_8744), .co(t_8745), .cout(t_8746));
compressor_4_2 u2_2997(.a(t_4712), .b(t_4709), .c(t_4706), .d(t_4703), .cin(t_8731), .o(t_8747), .co(t_8748), .cout(t_8749));
compressor_4_2 u2_2998(.a(t_4724), .b(t_4721), .c(t_4718), .d(t_4715), .cin(t_8734), .o(t_8750), .co(t_8751), .cout(t_8752));
compressor_4_2 u2_2999(.a(t_4701), .b(t_4698), .c(t_4695), .d(t_4692), .cin(t_8737), .o(t_8753), .co(t_8754), .cout(t_8755));
compressor_4_2 u2_3000(.a(t_4713), .b(t_4710), .c(t_4707), .d(t_4704), .cin(t_8740), .o(t_8756), .co(t_8757), .cout(t_8758));
compressor_4_2 u2_3001(.a(t_4725), .b(t_4722), .c(t_4719), .d(t_4716), .cin(t_8743), .o(t_8759), .co(t_8760), .cout(t_8761));
compressor_4_2 u2_3002(.a(t_4735), .b(t_4732), .c(t_4729), .d(t_4726), .cin(t_8746), .o(t_8762), .co(t_8763), .cout(t_8764));
compressor_4_2 u2_3003(.a(t_4747), .b(t_4744), .c(t_4741), .d(t_4738), .cin(t_8749), .o(t_8765), .co(t_8766), .cout(t_8767));
compressor_4_2 u2_3004(.a(t_4759), .b(t_4756), .c(t_4753), .d(t_4750), .cin(t_8752), .o(t_8768), .co(t_8769), .cout(t_8770));
compressor_4_2 u2_3005(.a(t_4736), .b(t_4733), .c(t_4730), .d(t_4727), .cin(t_8755), .o(t_8771), .co(t_8772), .cout(t_8773));
compressor_4_2 u2_3006(.a(t_4748), .b(t_4745), .c(t_4742), .d(t_4739), .cin(t_8758), .o(t_8774), .co(t_8775), .cout(t_8776));
compressor_4_2 u2_3007(.a(t_4760), .b(t_4757), .c(t_4754), .d(t_4751), .cin(t_8761), .o(t_8777), .co(t_8778), .cout(t_8779));
compressor_4_2 u2_3008(.a(t_4770), .b(t_4767), .c(t_4764), .d(t_4761), .cin(t_8764), .o(t_8780), .co(t_8781), .cout(t_8782));
compressor_4_2 u2_3009(.a(t_4782), .b(t_4779), .c(t_4776), .d(t_4773), .cin(t_8767), .o(t_8783), .co(t_8784), .cout(t_8785));
compressor_4_2 u2_3010(.a(t_4794), .b(t_4791), .c(t_4788), .d(t_4785), .cin(t_8770), .o(t_8786), .co(t_8787), .cout(t_8788));
compressor_4_2 u2_3011(.a(t_4768), .b(t_4765), .c(t_4762), .d(s_168_44), .cin(t_8773), .o(t_8789), .co(t_8790), .cout(t_8791));
compressor_4_2 u2_3012(.a(t_4780), .b(t_4777), .c(t_4774), .d(t_4771), .cin(t_8776), .o(t_8792), .co(t_8793), .cout(t_8794));
compressor_4_2 u2_3013(.a(t_4792), .b(t_4789), .c(t_4786), .d(t_4783), .cin(t_8779), .o(t_8795), .co(t_8796), .cout(t_8797));
compressor_4_2 u2_3014(.a(t_4802), .b(t_4799), .c(t_4796), .d(t_4795), .cin(t_8782), .o(t_8798), .co(t_8799), .cout(t_8800));
compressor_4_2 u2_3015(.a(t_4814), .b(t_4811), .c(t_4808), .d(t_4805), .cin(t_8785), .o(t_8801), .co(t_8802), .cout(t_8803));
compressor_4_2 u2_3016(.a(t_4826), .b(t_4823), .c(t_4820), .d(t_4817), .cin(t_8788), .o(t_8804), .co(t_8805), .cout(t_8806));
compressor_4_2 u2_3017(.a(t_4803), .b(t_4800), .c(t_4797), .d(s_169_44), .cin(t_8791), .o(t_8807), .co(t_8808), .cout(t_8809));
compressor_4_2 u2_3018(.a(t_4815), .b(t_4812), .c(t_4809), .d(t_4806), .cin(t_8794), .o(t_8810), .co(t_8811), .cout(t_8812));
compressor_4_2 u2_3019(.a(t_4827), .b(t_4824), .c(t_4821), .d(t_4818), .cin(t_8797), .o(t_8813), .co(t_8814), .cout(t_8815));
compressor_4_2 u2_3020(.a(t_4838), .b(t_4835), .c(t_4832), .d(t_4829), .cin(t_8800), .o(t_8816), .co(t_8817), .cout(t_8818));
compressor_4_2 u2_3021(.a(t_4850), .b(t_4847), .c(t_4844), .d(t_4841), .cin(t_8803), .o(t_8819), .co(t_8820), .cout(t_8821));
compressor_3_2 u1_3022(.a(t_4856), .b(t_4853), .cin(t_8806), .o(t_8822), .cout(t_8823));
compressor_4_2 u2_3023(.a(t_4839), .b(t_4836), .c(t_4833), .d(t_4830), .cin(t_8809), .o(t_8824), .co(t_8825), .cout(t_8826));
compressor_4_2 u2_3024(.a(t_4851), .b(t_4848), .c(t_4845), .d(t_4842), .cin(t_8812), .o(t_8827), .co(t_8828), .cout(t_8829));
compressor_4_2 u2_3025(.a(t_4862), .b(t_4860), .c(t_4857), .d(t_4854), .cin(t_8815), .o(t_8830), .co(t_8831), .cout(t_8832));
compressor_4_2 u2_3026(.a(t_4874), .b(t_4871), .c(t_4868), .d(t_4865), .cin(t_8818), .o(t_8833), .co(t_8834), .cout(t_8835));
compressor_4_2 u2_3027(.a(t_4886), .b(t_4883), .c(t_4880), .d(t_4877), .cin(t_8821), .o(t_8836), .co(t_8837), .cout(t_8838));
half_adder u0_3028(.a(t_4892), .b(t_4889), .o(t_8839), .cout(t_8840));
compressor_4_2 u2_3029(.a(t_4872), .b(t_4869), .c(t_4866), .d(t_4863), .cin(t_8826), .o(t_8841), .co(t_8842), .cout(t_8843));
compressor_4_2 u2_3030(.a(t_4884), .b(t_4881), .c(t_4878), .d(t_4875), .cin(t_8829), .o(t_8844), .co(t_8845), .cout(t_8846));
compressor_4_2 u2_3031(.a(t_4895), .b(t_4893), .c(t_4890), .d(t_4887), .cin(t_8832), .o(t_8847), .co(t_8848), .cout(t_8849));
compressor_4_2 u2_3032(.a(t_4907), .b(t_4904), .c(t_4901), .d(t_4898), .cin(t_8835), .o(t_8850), .co(t_8851), .cout(t_8852));
compressor_4_2 u2_3033(.a(t_4919), .b(t_4916), .c(t_4913), .d(t_4910), .cin(t_8838), .o(t_8853), .co(t_8854), .cout(t_8855));
half_adder u0_3034(.a(t_4925), .b(t_4922), .o(t_8856), .cout(t_8857));
compressor_4_2 u2_3035(.a(t_4902), .b(t_4899), .c(t_4896), .d(s_172_42), .cin(t_8843), .o(t_8858), .co(t_8859), .cout(t_8860));
compressor_4_2 u2_3036(.a(t_4914), .b(t_4911), .c(t_4908), .d(t_4905), .cin(t_8846), .o(t_8861), .co(t_8862), .cout(t_8863));
compressor_4_2 u2_3037(.a(t_4926), .b(t_4923), .c(t_4920), .d(t_4917), .cin(t_8849), .o(t_8864), .co(t_8865), .cout(t_8866));
compressor_4_2 u2_3038(.a(t_4937), .b(t_4934), .c(t_4931), .d(t_4928), .cin(t_8852), .o(t_8867), .co(t_8868), .cout(t_8869));
compressor_4_2 u2_3039(.a(t_4949), .b(t_4946), .c(t_4943), .d(t_4940), .cin(t_8855), .o(t_8870), .co(t_8871), .cout(t_8872));
compressor_3_2 u1_3040(.a(t_4958), .b(t_4955), .cin(t_4952), .o(t_8873), .cout(t_8874));
compressor_4_2 u2_3041(.a(t_4938), .b(t_4935), .c(t_4932), .d(t_4929), .cin(t_8860), .o(t_8875), .co(t_8876), .cout(t_8877));
compressor_4_2 u2_3042(.a(t_4950), .b(t_4947), .c(t_4944), .d(t_4941), .cin(t_8863), .o(t_8878), .co(t_8879), .cout(t_8880));
compressor_4_2 u2_3043(.a(t_4960), .b(t_4959), .c(t_4956), .d(t_4953), .cin(t_8866), .o(t_8881), .co(t_8882), .cout(t_8883));
compressor_4_2 u2_3044(.a(t_4972), .b(t_4969), .c(t_4966), .d(t_4963), .cin(t_8869), .o(t_8884), .co(t_8885), .cout(t_8886));
compressor_4_2 u2_3045(.a(t_4984), .b(t_4981), .c(t_4978), .d(t_4975), .cin(t_8872), .o(t_8887), .co(t_8888), .cout(t_8889));
half_adder u0_3046(.a(t_4990), .b(t_4987), .o(t_8890), .cout(t_8891));
compressor_4_2 u2_3047(.a(t_4970), .b(t_4967), .c(t_4964), .d(t_4961), .cin(t_8877), .o(t_8892), .co(t_8893), .cout(t_8894));
compressor_4_2 u2_3048(.a(t_4982), .b(t_4979), .c(t_4976), .d(t_4973), .cin(t_8880), .o(t_8895), .co(t_8896), .cout(t_8897));
compressor_4_2 u2_3049(.a(t_4992), .b(t_4991), .c(t_4988), .d(t_4985), .cin(t_8883), .o(t_8898), .co(t_8899), .cout(t_8900));
compressor_4_2 u2_3050(.a(t_5004), .b(t_5001), .c(t_4998), .d(t_4995), .cin(t_8886), .o(t_8901), .co(t_8902), .cout(t_8903));
compressor_4_2 u2_3051(.a(t_5016), .b(t_5013), .c(t_5010), .d(t_5007), .cin(t_8889), .o(t_8904), .co(t_8905), .cout(t_8906));
half_adder u0_3052(.a(t_5022), .b(t_5019), .o(t_8907), .cout(t_8908));
compressor_4_2 u2_3053(.a(t_5002), .b(t_4999), .c(t_4996), .d(t_4993), .cin(t_8894), .o(t_8909), .co(t_8910), .cout(t_8911));
compressor_4_2 u2_3054(.a(t_5014), .b(t_5011), .c(t_5008), .d(t_5005), .cin(t_8897), .o(t_8912), .co(t_8913), .cout(t_8914));
compressor_4_2 u2_3055(.a(t_5024), .b(t_5023), .c(t_5020), .d(t_5017), .cin(t_8900), .o(t_8915), .co(t_8916), .cout(t_8917));
compressor_4_2 u2_3056(.a(t_5036), .b(t_5033), .c(t_5030), .d(t_5027), .cin(t_8903), .o(t_8918), .co(t_8919), .cout(t_8920));
compressor_4_2 u2_3057(.a(t_5048), .b(t_5045), .c(t_5042), .d(t_5039), .cin(t_8906), .o(t_8921), .co(t_8922), .cout(t_8923));
half_adder u0_3058(.a(t_5054), .b(t_5051), .o(t_8924), .cout(t_8925));
compressor_4_2 u2_3059(.a(t_5031), .b(t_5028), .c(t_5025), .d(s_176_40), .cin(t_8911), .o(t_8926), .co(t_8927), .cout(t_8928));
compressor_4_2 u2_3060(.a(t_5043), .b(t_5040), .c(t_5037), .d(t_5034), .cin(t_8914), .o(t_8929), .co(t_8930), .cout(t_8931));
compressor_4_2 u2_3061(.a(t_5055), .b(t_5052), .c(t_5049), .d(t_5046), .cin(t_8917), .o(t_8932), .co(t_8933), .cout(t_8934));
compressor_4_2 u2_3062(.a(t_5065), .b(t_5062), .c(t_5059), .d(t_5056), .cin(t_8920), .o(t_8935), .co(t_8936), .cout(t_8937));
compressor_4_2 u2_3063(.a(t_5077), .b(t_5074), .c(t_5071), .d(t_5068), .cin(t_8923), .o(t_8938), .co(t_8939), .cout(t_8940));
half_adder u0_3064(.a(t_5083), .b(t_5080), .o(t_8941), .cout(t_8942));
compressor_4_2 u2_3065(.a(t_5063), .b(t_5060), .c(t_5057), .d(s_177_40), .cin(t_8928), .o(t_8943), .co(t_8944), .cout(t_8945));
compressor_4_2 u2_3066(.a(t_5075), .b(t_5072), .c(t_5069), .d(t_5066), .cin(t_8931), .o(t_8946), .co(t_8947), .cout(t_8948));
compressor_4_2 u2_3067(.a(t_5086), .b(t_5084), .c(t_5081), .d(t_5078), .cin(t_8934), .o(t_8949), .co(t_8950), .cout(t_8951));
compressor_4_2 u2_3068(.a(t_5098), .b(t_5095), .c(t_5092), .d(t_5089), .cin(t_8937), .o(t_8952), .co(t_8953), .cout(t_8954));
compressor_4_2 u2_3069(.a(t_5110), .b(t_5107), .c(t_5104), .d(t_5101), .cin(t_8940), .o(t_8955), .co(t_8956), .cout(t_8957));
compressor_4_2 u2_3070(.a(t_5096), .b(t_5093), .c(t_5090), .d(t_5087), .cin(t_8945), .o(t_8958), .co(t_8959), .cout(t_8960));
compressor_4_2 u2_3071(.a(t_5108), .b(t_5105), .c(t_5102), .d(t_5099), .cin(t_8948), .o(t_8961), .co(t_8962), .cout(t_8963));
compressor_4_2 u2_3072(.a(t_5119), .b(t_5116), .c(t_5114), .d(t_5111), .cin(t_8951), .o(t_8964), .co(t_8965), .cout(t_8966));
compressor_4_2 u2_3073(.a(t_5131), .b(t_5128), .c(t_5125), .d(t_5122), .cin(t_8954), .o(t_8967), .co(t_8968), .cout(t_8969));
compressor_4_2 u2_3074(.a(t_5143), .b(t_5140), .c(t_5137), .d(t_5134), .cin(t_8957), .o(t_8970), .co(t_8971), .cout(t_8972));
compressor_4_2 u2_3075(.a(t_5126), .b(t_5123), .c(t_5120), .d(t_5117), .cin(t_8960), .o(t_8973), .co(t_8974), .cout(t_8975));
compressor_4_2 u2_3076(.a(t_5138), .b(t_5135), .c(t_5132), .d(t_5129), .cin(t_8963), .o(t_8976), .co(t_8977), .cout(t_8978));
compressor_4_2 u2_3077(.a(t_5149), .b(t_5146), .c(t_5144), .d(t_5141), .cin(t_8966), .o(t_8979), .co(t_8980), .cout(t_8981));
compressor_4_2 u2_3078(.a(t_5161), .b(t_5158), .c(t_5155), .d(t_5152), .cin(t_8969), .o(t_8982), .co(t_8983), .cout(t_8984));
compressor_4_2 u2_3079(.a(t_5173), .b(t_5170), .c(t_5167), .d(t_5164), .cin(t_8972), .o(t_8985), .co(t_8986), .cout(t_8987));
compressor_4_2 u2_3080(.a(t_5153), .b(t_5150), .c(t_5147), .d(s_180_38), .cin(t_8975), .o(t_8988), .co(t_8989), .cout(t_8990));
compressor_4_2 u2_3081(.a(t_5165), .b(t_5162), .c(t_5159), .d(t_5156), .cin(t_8978), .o(t_8991), .co(t_8992), .cout(t_8993));
compressor_4_2 u2_3082(.a(t_5176), .b(t_5174), .c(t_5171), .d(t_5168), .cin(t_8981), .o(t_8994), .co(t_8995), .cout(t_8996));
compressor_4_2 u2_3083(.a(t_5188), .b(t_5185), .c(t_5182), .d(t_5179), .cin(t_8984), .o(t_8997), .co(t_8998), .cout(t_8999));
compressor_4_2 u2_3084(.a(t_5200), .b(t_5197), .c(t_5194), .d(t_5191), .cin(t_8987), .o(t_9000), .co(t_9001), .cout(t_9002));
compressor_4_2 u2_3085(.a(t_5186), .b(t_5183), .c(t_5180), .d(t_5177), .cin(t_8990), .o(t_9003), .co(t_9004), .cout(t_9005));
compressor_4_2 u2_3086(.a(t_5198), .b(t_5195), .c(t_5192), .d(t_5189), .cin(t_8993), .o(t_9006), .co(t_9007), .cout(t_9008));
compressor_4_2 u2_3087(.a(t_5208), .b(t_5205), .c(t_5204), .d(t_5201), .cin(t_8996), .o(t_9009), .co(t_9010), .cout(t_9011));
compressor_4_2 u2_3088(.a(t_5220), .b(t_5217), .c(t_5214), .d(t_5211), .cin(t_8999), .o(t_9012), .co(t_9013), .cout(t_9014));
compressor_4_2 u2_3089(.a(t_5232), .b(t_5229), .c(t_5226), .d(t_5223), .cin(t_9002), .o(t_9015), .co(t_9016), .cout(t_9017));
compressor_4_2 u2_3090(.a(t_5215), .b(t_5212), .c(t_5209), .d(t_5206), .cin(t_9005), .o(t_9018), .co(t_9019), .cout(t_9020));
compressor_4_2 u2_3091(.a(t_5227), .b(t_5224), .c(t_5221), .d(t_5218), .cin(t_9008), .o(t_9021), .co(t_9022), .cout(t_9023));
compressor_4_2 u2_3092(.a(t_5237), .b(t_5234), .c(t_5233), .d(t_5230), .cin(t_9011), .o(t_9024), .co(t_9025), .cout(t_9026));
compressor_4_2 u2_3093(.a(t_5249), .b(t_5246), .c(t_5243), .d(t_5240), .cin(t_9014), .o(t_9027), .co(t_9028), .cout(t_9029));
compressor_4_2 u2_3094(.a(t_5261), .b(t_5258), .c(t_5255), .d(t_5252), .cin(t_9017), .o(t_9030), .co(t_9031), .cout(t_9032));
compressor_4_2 u2_3095(.a(t_5244), .b(t_5241), .c(t_5238), .d(t_5235), .cin(t_9020), .o(t_9033), .co(t_9034), .cout(t_9035));
compressor_4_2 u2_3096(.a(t_5256), .b(t_5253), .c(t_5250), .d(t_5247), .cin(t_9023), .o(t_9036), .co(t_9037), .cout(t_9038));
compressor_4_2 u2_3097(.a(t_5266), .b(t_5263), .c(t_5262), .d(t_5259), .cin(t_9026), .o(t_9039), .co(t_9040), .cout(t_9041));
compressor_4_2 u2_3098(.a(t_5278), .b(t_5275), .c(t_5272), .d(t_5269), .cin(t_9029), .o(t_9042), .co(t_9043), .cout(t_9044));
compressor_4_2 u2_3099(.a(t_5290), .b(t_5287), .c(t_5284), .d(t_5281), .cin(t_9032), .o(t_9045), .co(t_9046), .cout(t_9047));
compressor_4_2 u2_3100(.a(t_5270), .b(t_5267), .c(t_5264), .d(s_184_36), .cin(t_9035), .o(t_9048), .co(t_9049), .cout(t_9050));
compressor_4_2 u2_3101(.a(t_5282), .b(t_5279), .c(t_5276), .d(t_5273), .cin(t_9038), .o(t_9051), .co(t_9052), .cout(t_9053));
compressor_4_2 u2_3102(.a(t_5292), .b(t_5291), .c(t_5288), .d(t_5285), .cin(t_9041), .o(t_9054), .co(t_9055), .cout(t_9056));
compressor_4_2 u2_3103(.a(t_5304), .b(t_5301), .c(t_5298), .d(t_5295), .cin(t_9044), .o(t_9057), .co(t_9058), .cout(t_9059));
compressor_4_2 u2_3104(.a(t_5316), .b(t_5313), .c(t_5310), .d(t_5307), .cin(t_9047), .o(t_9060), .co(t_9061), .cout(t_9062));
compressor_4_2 u2_3105(.a(t_5299), .b(t_5296), .c(t_5293), .d(s_185_36), .cin(t_9050), .o(t_9063), .co(t_9064), .cout(t_9065));
compressor_4_2 u2_3106(.a(t_5311), .b(t_5308), .c(t_5305), .d(t_5302), .cin(t_9053), .o(t_9066), .co(t_9067), .cout(t_9068));
compressor_4_2 u2_3107(.a(t_5322), .b(t_5319), .c(t_5317), .d(t_5314), .cin(t_9056), .o(t_9069), .co(t_9070), .cout(t_9071));
compressor_4_2 u2_3108(.a(t_5334), .b(t_5331), .c(t_5328), .d(t_5325), .cin(t_9059), .o(t_9072), .co(t_9073), .cout(t_9074));
compressor_3_2 u1_3109(.a(t_5340), .b(t_5337), .cin(t_9062), .o(t_9075), .cout(t_9076));
compressor_4_2 u2_3110(.a(t_5329), .b(t_5326), .c(t_5323), .d(t_5320), .cin(t_9065), .o(t_9077), .co(t_9078), .cout(t_9079));
compressor_4_2 u2_3111(.a(t_5341), .b(t_5338), .c(t_5335), .d(t_5332), .cin(t_9068), .o(t_9080), .co(t_9081), .cout(t_9082));
compressor_4_2 u2_3112(.a(t_5352), .b(t_5349), .c(t_5346), .d(t_5344), .cin(t_9071), .o(t_9083), .co(t_9084), .cout(t_9085));
compressor_4_2 u2_3113(.a(t_5364), .b(t_5361), .c(t_5358), .d(t_5355), .cin(t_9074), .o(t_9086), .co(t_9087), .cout(t_9088));
half_adder u0_3114(.a(t_5370), .b(t_5367), .o(t_9089), .cout(t_9090));
compressor_4_2 u2_3115(.a(t_5356), .b(t_5353), .c(t_5350), .d(t_5347), .cin(t_9079), .o(t_9091), .co(t_9092), .cout(t_9093));
compressor_4_2 u2_3116(.a(t_5368), .b(t_5365), .c(t_5362), .d(t_5359), .cin(t_9082), .o(t_9094), .co(t_9095), .cout(t_9096));
compressor_4_2 u2_3117(.a(t_5379), .b(t_5376), .c(t_5373), .d(t_5371), .cin(t_9085), .o(t_9097), .co(t_9098), .cout(t_9099));
compressor_4_2 u2_3118(.a(t_5391), .b(t_5388), .c(t_5385), .d(t_5382), .cin(t_9088), .o(t_9100), .co(t_9101), .cout(t_9102));
half_adder u0_3119(.a(t_5397), .b(t_5394), .o(t_9103), .cout(t_9104));
compressor_4_2 u2_3120(.a(t_5380), .b(t_5377), .c(t_5374), .d(s_188_34), .cin(t_9093), .o(t_9105), .co(t_9106), .cout(t_9107));
compressor_4_2 u2_3121(.a(t_5392), .b(t_5389), .c(t_5386), .d(t_5383), .cin(t_9096), .o(t_9108), .co(t_9109), .cout(t_9110));
compressor_4_2 u2_3122(.a(t_5403), .b(t_5400), .c(t_5398), .d(t_5395), .cin(t_9099), .o(t_9111), .co(t_9112), .cout(t_9113));
compressor_4_2 u2_3123(.a(t_5415), .b(t_5412), .c(t_5409), .d(t_5406), .cin(t_9102), .o(t_9114), .co(t_9115), .cout(t_9116));
compressor_3_2 u1_3124(.a(t_5424), .b(t_5421), .cin(t_5418), .o(t_9117), .cout(t_9118));
compressor_4_2 u2_3125(.a(t_5410), .b(t_5407), .c(t_5404), .d(t_5401), .cin(t_9107), .o(t_9119), .co(t_9120), .cout(t_9121));
compressor_4_2 u2_3126(.a(t_5422), .b(t_5419), .c(t_5416), .d(t_5413), .cin(t_9110), .o(t_9122), .co(t_9123), .cout(t_9124));
compressor_4_2 u2_3127(.a(t_5432), .b(t_5429), .c(t_5426), .d(t_5425), .cin(t_9113), .o(t_9125), .co(t_9126), .cout(t_9127));
compressor_4_2 u2_3128(.a(t_5444), .b(t_5441), .c(t_5438), .d(t_5435), .cin(t_9116), .o(t_9128), .co(t_9129), .cout(t_9130));
half_adder u0_3129(.a(t_5450), .b(t_5447), .o(t_9131), .cout(t_9132));
compressor_4_2 u2_3130(.a(t_5436), .b(t_5433), .c(t_5430), .d(t_5427), .cin(t_9121), .o(t_9133), .co(t_9134), .cout(t_9135));
compressor_4_2 u2_3131(.a(t_5448), .b(t_5445), .c(t_5442), .d(t_5439), .cin(t_9124), .o(t_9136), .co(t_9137), .cout(t_9138));
compressor_4_2 u2_3132(.a(t_5458), .b(t_5455), .c(t_5452), .d(t_5451), .cin(t_9127), .o(t_9139), .co(t_9140), .cout(t_9141));
compressor_4_2 u2_3133(.a(t_5470), .b(t_5467), .c(t_5464), .d(t_5461), .cin(t_9130), .o(t_9142), .co(t_9143), .cout(t_9144));
half_adder u0_3134(.a(t_5476), .b(t_5473), .o(t_9145), .cout(t_9146));
compressor_4_2 u2_3135(.a(t_5462), .b(t_5459), .c(t_5456), .d(t_5453), .cin(t_9135), .o(t_9147), .co(t_9148), .cout(t_9149));
compressor_4_2 u2_3136(.a(t_5474), .b(t_5471), .c(t_5468), .d(t_5465), .cin(t_9138), .o(t_9150), .co(t_9151), .cout(t_9152));
compressor_4_2 u2_3137(.a(t_5484), .b(t_5481), .c(t_5478), .d(t_5477), .cin(t_9141), .o(t_9153), .co(t_9154), .cout(t_9155));
compressor_4_2 u2_3138(.a(t_5496), .b(t_5493), .c(t_5490), .d(t_5487), .cin(t_9144), .o(t_9156), .co(t_9157), .cout(t_9158));
half_adder u0_3139(.a(t_5502), .b(t_5499), .o(t_9159), .cout(t_9160));
compressor_4_2 u2_3140(.a(t_5485), .b(t_5482), .c(t_5479), .d(s_192_32), .cin(t_9149), .o(t_9161), .co(t_9162), .cout(t_9163));
compressor_4_2 u2_3141(.a(t_5497), .b(t_5494), .c(t_5491), .d(t_5488), .cin(t_9152), .o(t_9164), .co(t_9165), .cout(t_9166));
compressor_4_2 u2_3142(.a(t_5507), .b(t_5504), .c(t_5503), .d(t_5500), .cin(t_9155), .o(t_9167), .co(t_9168), .cout(t_9169));
compressor_4_2 u2_3143(.a(t_5519), .b(t_5516), .c(t_5513), .d(t_5510), .cin(t_9158), .o(t_9170), .co(t_9171), .cout(t_9172));
half_adder u0_3144(.a(t_5525), .b(t_5522), .o(t_9173), .cout(t_9174));
compressor_4_2 u2_3145(.a(t_5511), .b(t_5508), .c(t_5505), .d(s_193_32), .cin(t_9163), .o(t_9175), .co(t_9176), .cout(t_9177));
compressor_4_2 u2_3146(.a(t_5523), .b(t_5520), .c(t_5517), .d(t_5514), .cin(t_9166), .o(t_9178), .co(t_9179), .cout(t_9180));
compressor_4_2 u2_3147(.a(t_5534), .b(t_5531), .c(t_5528), .d(t_5526), .cin(t_9169), .o(t_9181), .co(t_9182), .cout(t_9183));
compressor_4_2 u2_3148(.a(t_5546), .b(t_5543), .c(t_5540), .d(t_5537), .cin(t_9172), .o(t_9184), .co(t_9185), .cout(t_9186));
compressor_4_2 u2_3149(.a(t_5538), .b(t_5535), .c(t_5532), .d(t_5529), .cin(t_9177), .o(t_9187), .co(t_9188), .cout(t_9189));
compressor_4_2 u2_3150(.a(t_5550), .b(t_5547), .c(t_5544), .d(t_5541), .cin(t_9180), .o(t_9190), .co(t_9191), .cout(t_9192));
compressor_4_2 u2_3151(.a(t_5561), .b(t_5558), .c(t_5555), .d(t_5552), .cin(t_9183), .o(t_9193), .co(t_9194), .cout(t_9195));
compressor_4_2 u2_3152(.a(t_5573), .b(t_5570), .c(t_5567), .d(t_5564), .cin(t_9186), .o(t_9196), .co(t_9197), .cout(t_9198));
compressor_4_2 u2_3153(.a(t_5562), .b(t_5559), .c(t_5556), .d(t_5553), .cin(t_9189), .o(t_9199), .co(t_9200), .cout(t_9201));
compressor_4_2 u2_3154(.a(t_5574), .b(t_5571), .c(t_5568), .d(t_5565), .cin(t_9192), .o(t_9202), .co(t_9203), .cout(t_9204));
compressor_4_2 u2_3155(.a(t_5585), .b(t_5582), .c(t_5579), .d(t_5576), .cin(t_9195), .o(t_9205), .co(t_9206), .cout(t_9207));
compressor_4_2 u2_3156(.a(t_5597), .b(t_5594), .c(t_5591), .d(t_5588), .cin(t_9198), .o(t_9208), .co(t_9209), .cout(t_9210));
compressor_4_2 u2_3157(.a(t_5583), .b(t_5580), .c(t_5577), .d(s_196_30), .cin(t_9201), .o(t_9211), .co(t_9212), .cout(t_9213));
compressor_4_2 u2_3158(.a(t_5595), .b(t_5592), .c(t_5589), .d(t_5586), .cin(t_9204), .o(t_9214), .co(t_9215), .cout(t_9216));
compressor_4_2 u2_3159(.a(t_5606), .b(t_5603), .c(t_5600), .d(t_5598), .cin(t_9207), .o(t_9217), .co(t_9218), .cout(t_9219));
compressor_4_2 u2_3160(.a(t_5618), .b(t_5615), .c(t_5612), .d(t_5609), .cin(t_9210), .o(t_9220), .co(t_9221), .cout(t_9222));
compressor_4_2 u2_3161(.a(t_5610), .b(t_5607), .c(t_5604), .d(t_5601), .cin(t_9213), .o(t_9223), .co(t_9224), .cout(t_9225));
compressor_4_2 u2_3162(.a(t_5622), .b(t_5619), .c(t_5616), .d(t_5613), .cin(t_9216), .o(t_9226), .co(t_9227), .cout(t_9228));
compressor_4_2 u2_3163(.a(t_5632), .b(t_5629), .c(t_5626), .d(t_5623), .cin(t_9219), .o(t_9229), .co(t_9230), .cout(t_9231));
compressor_4_2 u2_3164(.a(t_5644), .b(t_5641), .c(t_5638), .d(t_5635), .cin(t_9222), .o(t_9232), .co(t_9233), .cout(t_9234));
compressor_4_2 u2_3165(.a(t_5633), .b(t_5630), .c(t_5627), .d(t_5624), .cin(t_9225), .o(t_9235), .co(t_9236), .cout(t_9237));
compressor_4_2 u2_3166(.a(t_5645), .b(t_5642), .c(t_5639), .d(t_5636), .cin(t_9228), .o(t_9238), .co(t_9239), .cout(t_9240));
compressor_4_2 u2_3167(.a(t_5655), .b(t_5652), .c(t_5649), .d(t_5646), .cin(t_9231), .o(t_9241), .co(t_9242), .cout(t_9243));
compressor_4_2 u2_3168(.a(t_5667), .b(t_5664), .c(t_5661), .d(t_5658), .cin(t_9234), .o(t_9244), .co(t_9245), .cout(t_9246));
compressor_4_2 u2_3169(.a(t_5656), .b(t_5653), .c(t_5650), .d(t_5647), .cin(t_9237), .o(t_9247), .co(t_9248), .cout(t_9249));
compressor_4_2 u2_3170(.a(t_5668), .b(t_5665), .c(t_5662), .d(t_5659), .cin(t_9240), .o(t_9250), .co(t_9251), .cout(t_9252));
compressor_4_2 u2_3171(.a(t_5678), .b(t_5675), .c(t_5672), .d(t_5669), .cin(t_9243), .o(t_9253), .co(t_9254), .cout(t_9255));
compressor_4_2 u2_3172(.a(t_5690), .b(t_5687), .c(t_5684), .d(t_5681), .cin(t_9246), .o(t_9256), .co(t_9257), .cout(t_9258));
compressor_4_2 u2_3173(.a(t_5676), .b(t_5673), .c(t_5670), .d(s_200_28), .cin(t_9249), .o(t_9259), .co(t_9260), .cout(t_9261));
compressor_4_2 u2_3174(.a(t_5688), .b(t_5685), .c(t_5682), .d(t_5679), .cin(t_9252), .o(t_9262), .co(t_9263), .cout(t_9264));
compressor_4_2 u2_3175(.a(t_5698), .b(t_5695), .c(t_5692), .d(t_5691), .cin(t_9255), .o(t_9265), .co(t_9266), .cout(t_9267));
compressor_4_2 u2_3176(.a(t_5710), .b(t_5707), .c(t_5704), .d(t_5701), .cin(t_9258), .o(t_9268), .co(t_9269), .cout(t_9270));
compressor_4_2 u2_3177(.a(t_5699), .b(t_5696), .c(t_5693), .d(s_201_28), .cin(t_9261), .o(t_9271), .co(t_9272), .cout(t_9273));
compressor_4_2 u2_3178(.a(t_5711), .b(t_5708), .c(t_5705), .d(t_5702), .cin(t_9264), .o(t_9274), .co(t_9275), .cout(t_9276));
compressor_4_2 u2_3179(.a(t_5722), .b(t_5719), .c(t_5716), .d(t_5713), .cin(t_9267), .o(t_9277), .co(t_9278), .cout(t_9279));
compressor_3_2 u1_3180(.a(t_5728), .b(t_5725), .cin(t_9270), .o(t_9280), .cout(t_9281));
compressor_4_2 u2_3181(.a(t_5723), .b(t_5720), .c(t_5717), .d(t_5714), .cin(t_9273), .o(t_9282), .co(t_9283), .cout(t_9284));
compressor_4_2 u2_3182(.a(t_5734), .b(t_5732), .c(t_5729), .d(t_5726), .cin(t_9276), .o(t_9285), .co(t_9286), .cout(t_9287));
compressor_4_2 u2_3183(.a(t_5746), .b(t_5743), .c(t_5740), .d(t_5737), .cin(t_9279), .o(t_9288), .co(t_9289), .cout(t_9290));
half_adder u0_3184(.a(t_5752), .b(t_5749), .o(t_9291), .cout(t_9292));
compressor_4_2 u2_3185(.a(t_5744), .b(t_5741), .c(t_5738), .d(t_5735), .cin(t_9284), .o(t_9293), .co(t_9294), .cout(t_9295));
compressor_4_2 u2_3186(.a(t_5755), .b(t_5753), .c(t_5750), .d(t_5747), .cin(t_9287), .o(t_9296), .co(t_9297), .cout(t_9298));
compressor_4_2 u2_3187(.a(t_5767), .b(t_5764), .c(t_5761), .d(t_5758), .cin(t_9290), .o(t_9299), .co(t_9300), .cout(t_9301));
half_adder u0_3188(.a(t_5773), .b(t_5770), .o(t_9302), .cout(t_9303));
compressor_4_2 u2_3189(.a(t_5762), .b(t_5759), .c(t_5756), .d(s_204_26), .cin(t_9295), .o(t_9304), .co(t_9305), .cout(t_9306));
compressor_4_2 u2_3190(.a(t_5774), .b(t_5771), .c(t_5768), .d(t_5765), .cin(t_9298), .o(t_9307), .co(t_9308), .cout(t_9309));
compressor_4_2 u2_3191(.a(t_5785), .b(t_5782), .c(t_5779), .d(t_5776), .cin(t_9301), .o(t_9310), .co(t_9311), .cout(t_9312));
compressor_3_2 u1_3192(.a(t_5794), .b(t_5791), .cin(t_5788), .o(t_9313), .cout(t_9314));
compressor_4_2 u2_3193(.a(t_5786), .b(t_5783), .c(t_5780), .d(t_5777), .cin(t_9306), .o(t_9315), .co(t_9316), .cout(t_9317));
compressor_4_2 u2_3194(.a(t_5796), .b(t_5795), .c(t_5792), .d(t_5789), .cin(t_9309), .o(t_9318), .co(t_9319), .cout(t_9320));
compressor_4_2 u2_3195(.a(t_5808), .b(t_5805), .c(t_5802), .d(t_5799), .cin(t_9312), .o(t_9321), .co(t_9322), .cout(t_9323));
half_adder u0_3196(.a(t_5814), .b(t_5811), .o(t_9324), .cout(t_9325));
compressor_4_2 u2_3197(.a(t_5806), .b(t_5803), .c(t_5800), .d(t_5797), .cin(t_9317), .o(t_9326), .co(t_9327), .cout(t_9328));
compressor_4_2 u2_3198(.a(t_5816), .b(t_5815), .c(t_5812), .d(t_5809), .cin(t_9320), .o(t_9329), .co(t_9330), .cout(t_9331));
compressor_4_2 u2_3199(.a(t_5828), .b(t_5825), .c(t_5822), .d(t_5819), .cin(t_9323), .o(t_9332), .co(t_9333), .cout(t_9334));
half_adder u0_3200(.a(t_5834), .b(t_5831), .o(t_9335), .cout(t_9336));
compressor_4_2 u2_3201(.a(t_5826), .b(t_5823), .c(t_5820), .d(t_5817), .cin(t_9328), .o(t_9337), .co(t_9338), .cout(t_9339));
compressor_4_2 u2_3202(.a(t_5836), .b(t_5835), .c(t_5832), .d(t_5829), .cin(t_9331), .o(t_9340), .co(t_9341), .cout(t_9342));
compressor_4_2 u2_3203(.a(t_5848), .b(t_5845), .c(t_5842), .d(t_5839), .cin(t_9334), .o(t_9343), .co(t_9344), .cout(t_9345));
half_adder u0_3204(.a(t_5854), .b(t_5851), .o(t_9346), .cout(t_9347));
compressor_4_2 u2_3205(.a(t_5843), .b(t_5840), .c(t_5837), .d(s_208_24), .cin(t_9339), .o(t_9348), .co(t_9349), .cout(t_9350));
compressor_4_2 u2_3206(.a(t_5855), .b(t_5852), .c(t_5849), .d(t_5846), .cin(t_9342), .o(t_9351), .co(t_9352), .cout(t_9353));
compressor_4_2 u2_3207(.a(t_5865), .b(t_5862), .c(t_5859), .d(t_5856), .cin(t_9345), .o(t_9354), .co(t_9355), .cout(t_9356));
half_adder u0_3208(.a(t_5871), .b(t_5868), .o(t_9357), .cout(t_9358));
compressor_4_2 u2_3209(.a(t_5863), .b(t_5860), .c(t_5857), .d(s_209_24), .cin(t_9350), .o(t_9359), .co(t_9360), .cout(t_9361));
compressor_4_2 u2_3210(.a(t_5874), .b(t_5872), .c(t_5869), .d(t_5866), .cin(t_9353), .o(t_9362), .co(t_9363), .cout(t_9364));
compressor_4_2 u2_3211(.a(t_5886), .b(t_5883), .c(t_5880), .d(t_5877), .cin(t_9356), .o(t_9365), .co(t_9366), .cout(t_9367));
compressor_4_2 u2_3212(.a(t_5884), .b(t_5881), .c(t_5878), .d(t_5875), .cin(t_9361), .o(t_9368), .co(t_9369), .cout(t_9370));
compressor_4_2 u2_3213(.a(t_5895), .b(t_5892), .c(t_5890), .d(t_5887), .cin(t_9364), .o(t_9371), .co(t_9372), .cout(t_9373));
compressor_4_2 u2_3214(.a(t_5907), .b(t_5904), .c(t_5901), .d(t_5898), .cin(t_9367), .o(t_9374), .co(t_9375), .cout(t_9376));
compressor_4_2 u2_3215(.a(t_5902), .b(t_5899), .c(t_5896), .d(t_5893), .cin(t_9370), .o(t_9377), .co(t_9378), .cout(t_9379));
compressor_4_2 u2_3216(.a(t_5913), .b(t_5910), .c(t_5908), .d(t_5905), .cin(t_9373), .o(t_9380), .co(t_9381), .cout(t_9382));
compressor_4_2 u2_3217(.a(t_5925), .b(t_5922), .c(t_5919), .d(t_5916), .cin(t_9376), .o(t_9383), .co(t_9384), .cout(t_9385));
compressor_4_2 u2_3218(.a(t_5917), .b(t_5914), .c(t_5911), .d(s_212_22), .cin(t_9379), .o(t_9386), .co(t_9387), .cout(t_9388));
compressor_4_2 u2_3219(.a(t_5928), .b(t_5926), .c(t_5923), .d(t_5920), .cin(t_9382), .o(t_9389), .co(t_9390), .cout(t_9391));
compressor_4_2 u2_3220(.a(t_5940), .b(t_5937), .c(t_5934), .d(t_5931), .cin(t_9385), .o(t_9392), .co(t_9393), .cout(t_9394));
compressor_4_2 u2_3221(.a(t_5938), .b(t_5935), .c(t_5932), .d(t_5929), .cin(t_9388), .o(t_9395), .co(t_9396), .cout(t_9397));
compressor_4_2 u2_3222(.a(t_5948), .b(t_5945), .c(t_5944), .d(t_5941), .cin(t_9391), .o(t_9398), .co(t_9399), .cout(t_9400));
compressor_4_2 u2_3223(.a(t_5960), .b(t_5957), .c(t_5954), .d(t_5951), .cin(t_9394), .o(t_9401), .co(t_9402), .cout(t_9403));
compressor_4_2 u2_3224(.a(t_5955), .b(t_5952), .c(t_5949), .d(t_5946), .cin(t_9397), .o(t_9404), .co(t_9405), .cout(t_9406));
compressor_4_2 u2_3225(.a(t_5965), .b(t_5962), .c(t_5961), .d(t_5958), .cin(t_9400), .o(t_9407), .co(t_9408), .cout(t_9409));
compressor_4_2 u2_3226(.a(t_5977), .b(t_5974), .c(t_5971), .d(t_5968), .cin(t_9403), .o(t_9410), .co(t_9411), .cout(t_9412));
compressor_4_2 u2_3227(.a(t_5972), .b(t_5969), .c(t_5966), .d(t_5963), .cin(t_9406), .o(t_9413), .co(t_9414), .cout(t_9415));
compressor_4_2 u2_3228(.a(t_5982), .b(t_5979), .c(t_5978), .d(t_5975), .cin(t_9409), .o(t_9416), .co(t_9417), .cout(t_9418));
compressor_4_2 u2_3229(.a(t_5994), .b(t_5991), .c(t_5988), .d(t_5985), .cin(t_9412), .o(t_9419), .co(t_9420), .cout(t_9421));
compressor_4_2 u2_3230(.a(t_5986), .b(t_5983), .c(t_5980), .d(s_216_20), .cin(t_9415), .o(t_9422), .co(t_9423), .cout(t_9424));
compressor_4_2 u2_3231(.a(t_5996), .b(t_5995), .c(t_5992), .d(t_5989), .cin(t_9418), .o(t_9425), .co(t_9426), .cout(t_9427));
compressor_4_2 u2_3232(.a(t_6008), .b(t_6005), .c(t_6002), .d(t_5999), .cin(t_9421), .o(t_9428), .co(t_9429), .cout(t_9430));
compressor_4_2 u2_3233(.a(t_6003), .b(t_6000), .c(t_5997), .d(s_217_20), .cin(t_9424), .o(t_9431), .co(t_9432), .cout(t_9433));
compressor_4_2 u2_3234(.a(t_6014), .b(t_6011), .c(t_6009), .d(t_6006), .cin(t_9427), .o(t_9434), .co(t_9435), .cout(t_9436));
compressor_3_2 u1_3235(.a(t_6020), .b(t_6017), .cin(t_9430), .o(t_9437), .cout(t_9438));
compressor_4_2 u2_3236(.a(t_6021), .b(t_6018), .c(t_6015), .d(t_6012), .cin(t_9433), .o(t_9439), .co(t_9440), .cout(t_9441));
compressor_4_2 u2_3237(.a(t_6032), .b(t_6029), .c(t_6026), .d(t_6024), .cin(t_9436), .o(t_9442), .co(t_9443), .cout(t_9444));
half_adder u0_3238(.a(t_6038), .b(t_6035), .o(t_9445), .cout(t_9446));
compressor_4_2 u2_3239(.a(t_6036), .b(t_6033), .c(t_6030), .d(t_6027), .cin(t_9441), .o(t_9447), .co(t_9448), .cout(t_9449));
compressor_4_2 u2_3240(.a(t_6047), .b(t_6044), .c(t_6041), .d(t_6039), .cin(t_9444), .o(t_9450), .co(t_9451), .cout(t_9452));
half_adder u0_3241(.a(t_6053), .b(t_6050), .o(t_9453), .cout(t_9454));
compressor_4_2 u2_3242(.a(t_6048), .b(t_6045), .c(t_6042), .d(s_220_18), .cin(t_9449), .o(t_9455), .co(t_9456), .cout(t_9457));
compressor_4_2 u2_3243(.a(t_6059), .b(t_6056), .c(t_6054), .d(t_6051), .cin(t_9452), .o(t_9458), .co(t_9459), .cout(t_9460));
compressor_3_2 u1_3244(.a(t_6068), .b(t_6065), .cin(t_6062), .o(t_9461), .cout(t_9462));
compressor_4_2 u2_3245(.a(t_6066), .b(t_6063), .c(t_6060), .d(t_6057), .cin(t_9457), .o(t_9463), .co(t_9464), .cout(t_9465));
compressor_4_2 u2_3246(.a(t_6076), .b(t_6073), .c(t_6070), .d(t_6069), .cin(t_9460), .o(t_9466), .co(t_9467), .cout(t_9468));
half_adder u0_3247(.a(t_6082), .b(t_6079), .o(t_9469), .cout(t_9470));
compressor_4_2 u2_3248(.a(t_6080), .b(t_6077), .c(t_6074), .d(t_6071), .cin(t_9465), .o(t_9471), .co(t_9472), .cout(t_9473));
compressor_4_2 u2_3249(.a(t_6090), .b(t_6087), .c(t_6084), .d(t_6083), .cin(t_9468), .o(t_9474), .co(t_9475), .cout(t_9476));
half_adder u0_3250(.a(t_6096), .b(t_6093), .o(t_9477), .cout(t_9478));
compressor_4_2 u2_3251(.a(t_6094), .b(t_6091), .c(t_6088), .d(t_6085), .cin(t_9473), .o(t_9479), .co(t_9480), .cout(t_9481));
compressor_4_2 u2_3252(.a(t_6104), .b(t_6101), .c(t_6098), .d(t_6097), .cin(t_9476), .o(t_9482), .co(t_9483), .cout(t_9484));
half_adder u0_3253(.a(t_6110), .b(t_6107), .o(t_9485), .cout(t_9486));
compressor_4_2 u2_3254(.a(t_6105), .b(t_6102), .c(t_6099), .d(s_224_16), .cin(t_9481), .o(t_9487), .co(t_9488), .cout(t_9489));
compressor_4_2 u2_3255(.a(t_6115), .b(t_6112), .c(t_6111), .d(t_6108), .cin(t_9484), .o(t_9490), .co(t_9491), .cout(t_9492));
half_adder u0_3256(.a(t_6121), .b(t_6118), .o(t_9493), .cout(t_9494));
compressor_4_2 u2_3257(.a(t_6119), .b(t_6116), .c(t_6113), .d(s_225_16), .cin(t_9489), .o(t_9495), .co(t_9496), .cout(t_9497));
compressor_4_2 u2_3258(.a(t_6130), .b(t_6127), .c(t_6124), .d(t_6122), .cin(t_9492), .o(t_9498), .co(t_9499), .cout(t_9500));
compressor_4_2 u2_3259(.a(t_6134), .b(t_6131), .c(t_6128), .d(t_6125), .cin(t_9497), .o(t_9501), .co(t_9502), .cout(t_9503));
compressor_4_2 u2_3260(.a(t_6145), .b(t_6142), .c(t_6139), .d(t_6136), .cin(t_9500), .o(t_9504), .co(t_9505), .cout(t_9506));
compressor_4_2 u2_3261(.a(t_6146), .b(t_6143), .c(t_6140), .d(t_6137), .cin(t_9503), .o(t_9507), .co(t_9508), .cout(t_9509));
compressor_4_2 u2_3262(.a(t_6157), .b(t_6154), .c(t_6151), .d(t_6148), .cin(t_9506), .o(t_9510), .co(t_9511), .cout(t_9512));
compressor_4_2 u2_3263(.a(t_6155), .b(t_6152), .c(t_6149), .d(s_228_14), .cin(t_9509), .o(t_9513), .co(t_9514), .cout(t_9515));
compressor_4_2 u2_3264(.a(t_6166), .b(t_6163), .c(t_6160), .d(t_6158), .cin(t_9512), .o(t_9516), .co(t_9517), .cout(t_9518));
compressor_4_2 u2_3265(.a(t_6170), .b(t_6167), .c(t_6164), .d(t_6161), .cin(t_9515), .o(t_9519), .co(t_9520), .cout(t_9521));
compressor_4_2 u2_3266(.a(t_6180), .b(t_6177), .c(t_6174), .d(t_6171), .cin(t_9518), .o(t_9522), .co(t_9523), .cout(t_9524));
compressor_4_2 u2_3267(.a(t_6181), .b(t_6178), .c(t_6175), .d(t_6172), .cin(t_9521), .o(t_9525), .co(t_9526), .cout(t_9527));
compressor_4_2 u2_3268(.a(t_6191), .b(t_6188), .c(t_6185), .d(t_6182), .cin(t_9524), .o(t_9528), .co(t_9529), .cout(t_9530));
compressor_4_2 u2_3269(.a(t_6192), .b(t_6189), .c(t_6186), .d(t_6183), .cin(t_9527), .o(t_9531), .co(t_9532), .cout(t_9533));
compressor_4_2 u2_3270(.a(t_6202), .b(t_6199), .c(t_6196), .d(t_6193), .cin(t_9530), .o(t_9534), .co(t_9535), .cout(t_9536));
compressor_4_2 u2_3271(.a(t_6200), .b(t_6197), .c(t_6194), .d(s_232_12), .cin(t_9533), .o(t_9537), .co(t_9538), .cout(t_9539));
compressor_4_2 u2_3272(.a(t_6210), .b(t_6207), .c(t_6204), .d(t_6203), .cin(t_9536), .o(t_9540), .co(t_9541), .cout(t_9542));
compressor_4_2 u2_3273(.a(t_6211), .b(t_6208), .c(t_6205), .d(s_233_12), .cin(t_9539), .o(t_9543), .co(t_9544), .cout(t_9545));
compressor_3_2 u1_3274(.a(t_6216), .b(t_6213), .cin(t_9542), .o(t_9546), .cout(t_9547));
compressor_4_2 u2_3275(.a(t_6222), .b(t_6220), .c(t_6217), .d(t_6214), .cin(t_9545), .o(t_9548), .co(t_9549), .cout(t_9550));
half_adder u0_3276(.a(t_6228), .b(t_6225), .o(t_9551), .cout(t_9552));
compressor_4_2 u2_3277(.a(t_6231), .b(t_6229), .c(t_6226), .d(t_6223), .cin(t_9550), .o(t_9553), .co(t_9554), .cout(t_9555));
half_adder u0_3278(.a(t_6237), .b(t_6234), .o(t_9556), .cout(t_9557));
compressor_4_2 u2_3279(.a(t_6238), .b(t_6235), .c(t_6232), .d(s_236_10), .cin(t_9555), .o(t_9558), .co(t_9559), .cout(t_9560));
compressor_3_2 u1_3280(.a(t_6246), .b(t_6243), .cin(t_6240), .o(t_9561), .cout(t_9562));
compressor_4_2 u2_3281(.a(t_6248), .b(t_6247), .c(t_6244), .d(t_6241), .cin(t_9560), .o(t_9563), .co(t_9564), .cout(t_9565));
half_adder u0_3282(.a(t_6254), .b(t_6251), .o(t_9566), .cout(t_9567));
compressor_4_2 u2_3283(.a(t_6256), .b(t_6255), .c(t_6252), .d(t_6249), .cin(t_9565), .o(t_9568), .co(t_9569), .cout(t_9570));
half_adder u0_3284(.a(t_6262), .b(t_6259), .o(t_9571), .cout(t_9572));
compressor_4_2 u2_3285(.a(t_6264), .b(t_6263), .c(t_6260), .d(t_6257), .cin(t_9570), .o(t_9573), .co(t_9574), .cout(t_9575));
half_adder u0_3286(.a(t_6270), .b(t_6267), .o(t_9576), .cout(t_9577));
compressor_4_2 u2_3287(.a(t_6271), .b(t_6268), .c(t_6265), .d(s_240_8), .cin(t_9575), .o(t_9578), .co(t_9579), .cout(t_9580));
half_adder u0_3288(.a(t_6275), .b(t_6272), .o(t_9581), .cout(t_9582));
compressor_4_2 u2_3289(.a(t_6278), .b(t_6276), .c(t_6273), .d(s_241_8), .cin(t_9580), .o(t_9583), .co(t_9584), .cout(t_9585));
compressor_4_2 u2_3290(.a(t_6287), .b(t_6284), .c(t_6282), .d(t_6279), .cin(t_9585), .o(t_9586), .co(t_9587), .cout(t_9588));
compressor_4_2 u2_3291(.a(t_6293), .b(t_6290), .c(t_6288), .d(t_6285), .cin(t_9588), .o(t_9589), .co(t_9590), .cout(t_9591));
compressor_4_2 u2_3292(.a(t_6296), .b(t_6294), .c(t_6291), .d(s_244_6), .cin(t_9591), .o(t_9592), .co(t_9593), .cout(t_9594));
compressor_4_2 u2_3293(.a(t_6304), .b(t_6301), .c(t_6300), .d(t_6297), .cin(t_9594), .o(t_9595), .co(t_9596), .cout(t_9597));
compressor_4_2 u2_3294(.a(t_6309), .b(t_6306), .c(t_6305), .d(t_6302), .cin(t_9597), .o(t_9598), .co(t_9599), .cout(t_9600));
compressor_4_2 u2_3295(.a(t_6314), .b(t_6311), .c(t_6310), .d(t_6307), .cin(t_9600), .o(t_9601), .co(t_9602), .cout(t_9603));
compressor_4_2 u2_3296(.a(t_6316), .b(t_6315), .c(t_6312), .d(s_248_4), .cin(t_9603), .o(t_9604), .co(t_9605), .cout(t_9606));
compressor_3_2 u1_3297(.a(t_6317), .b(s_249_4), .cin(t_9606), .o(t_9607), .cout(t_9608));
half_adder u0_3298(.a(t_6322), .b(t_6320), .o(t_9609), .cout(t_9610));
half_adder u0_3299(.a(t_6325), .b(t_6323), .o(t_9611), .cout(t_9612));
compressor_3_2 u1_3300(.a(t_6328), .b(t_6326), .cin(s_252_2), .o(t_9613), .cout(t_9614));
half_adder u0_3301(.a(t_6330), .b(t_6329), .o(t_9615), .cout(t_9616));
half_adder u0_3302(.a(t_6332), .b(t_6331), .o(t_9617), .cout(t_9618));
half_adder u0_3303(.a(t_6334), .b(t_6333), .o(t_9619), .cout());

/* u0_3304 Output nets */
wire t_9620,   t_9621;
/* u0_3305 Output nets */
wire t_9622,   t_9623;
/* u0_3306 Output nets */
wire t_9624,   t_9625;
/* u0_3307 Output nets */
wire t_9626,   t_9627;
/* u0_3308 Output nets */
wire t_9628,   t_9629;
/* u0_3309 Output nets */
wire t_9630,   t_9631;
/* u1_3310 Output nets */
wire t_9632,   t_9633;
/* u0_3311 Output nets */
wire t_9634,   t_9635;
/* u1_3312 Output nets */
wire t_9636,   t_9637;
/* u0_3313 Output nets */
wire t_9638,   t_9639;
/* u0_3314 Output nets */
wire t_9640,   t_9641;
/* u0_3315 Output nets */
wire t_9642,   t_9643;
/* u0_3316 Output nets */
wire t_9644,   t_9645;
/* u1_3317 Output nets */
wire t_9646,   t_9647;
/* u1_3318 Output nets */
wire t_9648,   t_9649;
/* u1_3319 Output nets */
wire t_9650,   t_9651;
/* u1_3320 Output nets */
wire t_9652,   t_9653;
/* u1_3321 Output nets */
wire t_9654,   t_9655;
/* u1_3322 Output nets */
wire t_9656,   t_9657;
/* u1_3323 Output nets */
wire t_9658,   t_9659;
/* u1_3324 Output nets */
wire t_9660,   t_9661;
/* u1_3325 Output nets */
wire t_9662,   t_9663;
/* u2_3326 Output nets */
wire t_9664,   t_9665,   t_9666;
/* u2_3327 Output nets */
wire t_9667,   t_9668,   t_9669;
/* u2_3328 Output nets */
wire t_9670,   t_9671,   t_9672;
/* u2_3329 Output nets */
wire t_9673,   t_9674,   t_9675;
/* u2_3330 Output nets */
wire t_9676,   t_9677,   t_9678;
/* u2_3331 Output nets */
wire t_9679,   t_9680,   t_9681;
/* u2_3332 Output nets */
wire t_9682,   t_9683,   t_9684;
/* u2_3333 Output nets */
wire t_9685,   t_9686,   t_9687;
/* u2_3334 Output nets */
wire t_9688,   t_9689,   t_9690;
/* u2_3335 Output nets */
wire t_9691,   t_9692,   t_9693;
/* u0_3336 Output nets */
wire t_9694,   t_9695;
/* u2_3337 Output nets */
wire t_9696,   t_9697,   t_9698;
/* u2_3338 Output nets */
wire t_9699,   t_9700,   t_9701;
/* u0_3339 Output nets */
wire t_9702,   t_9703;
/* u2_3340 Output nets */
wire t_9704,   t_9705,   t_9706;
/* u0_3341 Output nets */
wire t_9707,   t_9708;
/* u2_3342 Output nets */
wire t_9709,   t_9710,   t_9711;
/* u0_3343 Output nets */
wire t_9712,   t_9713;
/* u2_3344 Output nets */
wire t_9714,   t_9715,   t_9716;
/* u0_3345 Output nets */
wire t_9717,   t_9718;
/* u2_3346 Output nets */
wire t_9719,   t_9720,   t_9721;
/* u0_3347 Output nets */
wire t_9722,   t_9723;
/* u2_3348 Output nets */
wire t_9724,   t_9725,   t_9726;
/* u1_3349 Output nets */
wire t_9727,   t_9728;
/* u2_3350 Output nets */
wire t_9729,   t_9730,   t_9731;
/* u0_3351 Output nets */
wire t_9732,   t_9733;
/* u2_3352 Output nets */
wire t_9734,   t_9735,   t_9736;
/* u1_3353 Output nets */
wire t_9737,   t_9738;
/* u2_3354 Output nets */
wire t_9739,   t_9740,   t_9741;
/* u0_3355 Output nets */
wire t_9742,   t_9743;
/* u2_3356 Output nets */
wire t_9744,   t_9745,   t_9746;
/* u0_3357 Output nets */
wire t_9747,   t_9748;
/* u2_3358 Output nets */
wire t_9749,   t_9750,   t_9751;
/* u0_3359 Output nets */
wire t_9752,   t_9753;
/* u2_3360 Output nets */
wire t_9754,   t_9755,   t_9756;
/* u0_3361 Output nets */
wire t_9757,   t_9758;
/* u2_3362 Output nets */
wire t_9759,   t_9760,   t_9761;
/* u1_3363 Output nets */
wire t_9762,   t_9763;
/* u2_3364 Output nets */
wire t_9764,   t_9765,   t_9766;
/* u1_3365 Output nets */
wire t_9767,   t_9768;
/* u2_3366 Output nets */
wire t_9769,   t_9770,   t_9771;
/* u1_3367 Output nets */
wire t_9772,   t_9773;
/* u2_3368 Output nets */
wire t_9774,   t_9775,   t_9776;
/* u1_3369 Output nets */
wire t_9777,   t_9778;
/* u2_3370 Output nets */
wire t_9779,   t_9780,   t_9781;
/* u1_3371 Output nets */
wire t_9782,   t_9783;
/* u2_3372 Output nets */
wire t_9784,   t_9785,   t_9786;
/* u1_3373 Output nets */
wire t_9787,   t_9788;
/* u2_3374 Output nets */
wire t_9789,   t_9790,   t_9791;
/* u1_3375 Output nets */
wire t_9792,   t_9793;
/* u2_3376 Output nets */
wire t_9794,   t_9795,   t_9796;
/* u1_3377 Output nets */
wire t_9797,   t_9798;
/* u2_3378 Output nets */
wire t_9799,   t_9800,   t_9801;
/* u1_3379 Output nets */
wire t_9802,   t_9803;
/* u2_3380 Output nets */
wire t_9804,   t_9805,   t_9806;
/* u2_3381 Output nets */
wire t_9807,   t_9808,   t_9809;
/* u2_3382 Output nets */
wire t_9810,   t_9811,   t_9812;
/* u2_3383 Output nets */
wire t_9813,   t_9814,   t_9815;
/* u2_3384 Output nets */
wire t_9816,   t_9817,   t_9818;
/* u2_3385 Output nets */
wire t_9819,   t_9820,   t_9821;
/* u2_3386 Output nets */
wire t_9822,   t_9823,   t_9824;
/* u2_3387 Output nets */
wire t_9825,   t_9826,   t_9827;
/* u2_3388 Output nets */
wire t_9828,   t_9829,   t_9830;
/* u2_3389 Output nets */
wire t_9831,   t_9832,   t_9833;
/* u2_3390 Output nets */
wire t_9834,   t_9835,   t_9836;
/* u2_3391 Output nets */
wire t_9837,   t_9838,   t_9839;
/* u2_3392 Output nets */
wire t_9840,   t_9841,   t_9842;
/* u2_3393 Output nets */
wire t_9843,   t_9844,   t_9845;
/* u2_3394 Output nets */
wire t_9846,   t_9847,   t_9848;
/* u2_3395 Output nets */
wire t_9849,   t_9850,   t_9851;
/* u2_3396 Output nets */
wire t_9852,   t_9853,   t_9854;
/* u2_3397 Output nets */
wire t_9855,   t_9856,   t_9857;
/* u2_3398 Output nets */
wire t_9858,   t_9859,   t_9860;
/* u2_3399 Output nets */
wire t_9861,   t_9862,   t_9863;
/* u0_3400 Output nets */
wire t_9864,   t_9865;
/* u2_3401 Output nets */
wire t_9866,   t_9867,   t_9868;
/* u2_3402 Output nets */
wire t_9869,   t_9870,   t_9871;
/* u2_3403 Output nets */
wire t_9872,   t_9873,   t_9874;
/* u2_3404 Output nets */
wire t_9875,   t_9876,   t_9877;
/* u0_3405 Output nets */
wire t_9878,   t_9879;
/* u2_3406 Output nets */
wire t_9880,   t_9881,   t_9882;
/* u2_3407 Output nets */
wire t_9883,   t_9884,   t_9885;
/* u0_3408 Output nets */
wire t_9886,   t_9887;
/* u2_3409 Output nets */
wire t_9888,   t_9889,   t_9890;
/* u2_3410 Output nets */
wire t_9891,   t_9892,   t_9893;
/* u0_3411 Output nets */
wire t_9894,   t_9895;
/* u2_3412 Output nets */
wire t_9896,   t_9897,   t_9898;
/* u2_3413 Output nets */
wire t_9899,   t_9900,   t_9901;
/* u0_3414 Output nets */
wire t_9902,   t_9903;
/* u2_3415 Output nets */
wire t_9904,   t_9905,   t_9906;
/* u2_3416 Output nets */
wire t_9907,   t_9908,   t_9909;
/* u0_3417 Output nets */
wire t_9910,   t_9911;
/* u2_3418 Output nets */
wire t_9912,   t_9913,   t_9914;
/* u2_3419 Output nets */
wire t_9915,   t_9916,   t_9917;
/* u1_3420 Output nets */
wire t_9918,   t_9919;
/* u2_3421 Output nets */
wire t_9920,   t_9921,   t_9922;
/* u2_3422 Output nets */
wire t_9923,   t_9924,   t_9925;
/* u0_3423 Output nets */
wire t_9926,   t_9927;
/* u2_3424 Output nets */
wire t_9928,   t_9929,   t_9930;
/* u2_3425 Output nets */
wire t_9931,   t_9932,   t_9933;
/* u1_3426 Output nets */
wire t_9934,   t_9935;
/* u2_3427 Output nets */
wire t_9936,   t_9937,   t_9938;
/* u2_3428 Output nets */
wire t_9939,   t_9940,   t_9941;
/* u0_3429 Output nets */
wire t_9942,   t_9943;
/* u2_3430 Output nets */
wire t_9944,   t_9945,   t_9946;
/* u2_3431 Output nets */
wire t_9947,   t_9948,   t_9949;
/* u0_3432 Output nets */
wire t_9950,   t_9951;
/* u2_3433 Output nets */
wire t_9952,   t_9953,   t_9954;
/* u2_3434 Output nets */
wire t_9955,   t_9956,   t_9957;
/* u0_3435 Output nets */
wire t_9958,   t_9959;
/* u2_3436 Output nets */
wire t_9960,   t_9961,   t_9962;
/* u2_3437 Output nets */
wire t_9963,   t_9964,   t_9965;
/* u0_3438 Output nets */
wire t_9966,   t_9967;
/* u2_3439 Output nets */
wire t_9968,   t_9969,   t_9970;
/* u2_3440 Output nets */
wire t_9971,   t_9972,   t_9973;
/* u1_3441 Output nets */
wire t_9974,   t_9975;
/* u2_3442 Output nets */
wire t_9976,   t_9977,   t_9978;
/* u2_3443 Output nets */
wire t_9979,   t_9980,   t_9981;
/* u1_3444 Output nets */
wire t_9982,   t_9983;
/* u2_3445 Output nets */
wire t_9984,   t_9985,   t_9986;
/* u2_3446 Output nets */
wire t_9987,   t_9988,   t_9989;
/* u1_3447 Output nets */
wire t_9990,   t_9991;
/* u2_3448 Output nets */
wire t_9992,   t_9993,   t_9994;
/* u2_3449 Output nets */
wire t_9995,   t_9996,   t_9997;
/* u1_3450 Output nets */
wire t_9998,   t_9999;
/* u2_3451 Output nets */
wire t_10000,  t_10001,  t_10002;
/* u2_3452 Output nets */
wire t_10003,  t_10004,  t_10005;
/* u1_3453 Output nets */
wire t_10006,  t_10007;
/* u2_3454 Output nets */
wire t_10008,  t_10009,  t_10010;
/* u2_3455 Output nets */
wire t_10011,  t_10012,  t_10013;
/* u1_3456 Output nets */
wire t_10014,  t_10015;
/* u2_3457 Output nets */
wire t_10016,  t_10017,  t_10018;
/* u2_3458 Output nets */
wire t_10019,  t_10020,  t_10021;
/* u1_3459 Output nets */
wire t_10022,  t_10023;
/* u2_3460 Output nets */
wire t_10024,  t_10025,  t_10026;
/* u2_3461 Output nets */
wire t_10027,  t_10028,  t_10029;
/* u1_3462 Output nets */
wire t_10030,  t_10031;
/* u2_3463 Output nets */
wire t_10032,  t_10033,  t_10034;
/* u2_3464 Output nets */
wire t_10035,  t_10036,  t_10037;
/* u1_3465 Output nets */
wire t_10038,  t_10039;
/* u2_3466 Output nets */
wire t_10040,  t_10041,  t_10042;
/* u2_3467 Output nets */
wire t_10043,  t_10044,  t_10045;
/* u2_3468 Output nets */
wire t_10046,  t_10047,  t_10048;
/* u2_3469 Output nets */
wire t_10049,  t_10050,  t_10051;
/* u2_3470 Output nets */
wire t_10052,  t_10053,  t_10054;
/* u2_3471 Output nets */
wire t_10055,  t_10056,  t_10057;
/* u2_3472 Output nets */
wire t_10058,  t_10059,  t_10060;
/* u2_3473 Output nets */
wire t_10061,  t_10062,  t_10063;
/* u2_3474 Output nets */
wire t_10064,  t_10065,  t_10066;
/* u2_3475 Output nets */
wire t_10067,  t_10068,  t_10069;
/* u2_3476 Output nets */
wire t_10070,  t_10071,  t_10072;
/* u2_3477 Output nets */
wire t_10073,  t_10074,  t_10075;
/* u2_3478 Output nets */
wire t_10076,  t_10077,  t_10078;
/* u2_3479 Output nets */
wire t_10079,  t_10080,  t_10081;
/* u2_3480 Output nets */
wire t_10082,  t_10083,  t_10084;
/* u2_3481 Output nets */
wire t_10085,  t_10086,  t_10087;
/* u2_3482 Output nets */
wire t_10088,  t_10089,  t_10090;
/* u2_3483 Output nets */
wire t_10091,  t_10092,  t_10093;
/* u2_3484 Output nets */
wire t_10094,  t_10095,  t_10096;
/* u2_3485 Output nets */
wire t_10097,  t_10098,  t_10099;
/* u2_3486 Output nets */
wire t_10100,  t_10101,  t_10102;
/* u2_3487 Output nets */
wire t_10103,  t_10104,  t_10105;
/* u2_3488 Output nets */
wire t_10106,  t_10107,  t_10108;
/* u2_3489 Output nets */
wire t_10109,  t_10110,  t_10111;
/* u2_3490 Output nets */
wire t_10112,  t_10113,  t_10114;
/* u2_3491 Output nets */
wire t_10115,  t_10116,  t_10117;
/* u2_3492 Output nets */
wire t_10118,  t_10119,  t_10120;
/* u2_3493 Output nets */
wire t_10121,  t_10122,  t_10123;
/* u2_3494 Output nets */
wire t_10124,  t_10125,  t_10126;
/* u2_3495 Output nets */
wire t_10127,  t_10128,  t_10129;
/* u0_3496 Output nets */
wire t_10130,  t_10131;
/* u2_3497 Output nets */
wire t_10132,  t_10133,  t_10134;
/* u2_3498 Output nets */
wire t_10135,  t_10136,  t_10137;
/* u2_3499 Output nets */
wire t_10138,  t_10139,  t_10140;
/* u2_3500 Output nets */
wire t_10141,  t_10142,  t_10143;
/* u2_3501 Output nets */
wire t_10144,  t_10145,  t_10146;
/* u2_3502 Output nets */
wire t_10147,  t_10148,  t_10149;
/* u0_3503 Output nets */
wire t_10150,  t_10151;
/* u2_3504 Output nets */
wire t_10152,  t_10153,  t_10154;
/* u2_3505 Output nets */
wire t_10155,  t_10156,  t_10157;
/* u2_3506 Output nets */
wire t_10158,  t_10159,  t_10160;
/* u0_3507 Output nets */
wire t_10161,  t_10162;
/* u2_3508 Output nets */
wire t_10163,  t_10164,  t_10165;
/* u2_3509 Output nets */
wire t_10166,  t_10167,  t_10168;
/* u2_3510 Output nets */
wire t_10169,  t_10170,  t_10171;
/* u0_3511 Output nets */
wire t_10172,  t_10173;
/* u2_3512 Output nets */
wire t_10174,  t_10175,  t_10176;
/* u2_3513 Output nets */
wire t_10177,  t_10178,  t_10179;
/* u2_3514 Output nets */
wire t_10180,  t_10181,  t_10182;
/* u0_3515 Output nets */
wire t_10183,  t_10184;
/* u2_3516 Output nets */
wire t_10185,  t_10186,  t_10187;
/* u2_3517 Output nets */
wire t_10188,  t_10189,  t_10190;
/* u2_3518 Output nets */
wire t_10191,  t_10192,  t_10193;
/* u0_3519 Output nets */
wire t_10194,  t_10195;
/* u2_3520 Output nets */
wire t_10196,  t_10197,  t_10198;
/* u2_3521 Output nets */
wire t_10199,  t_10200,  t_10201;
/* u2_3522 Output nets */
wire t_10202,  t_10203,  t_10204;
/* u1_3523 Output nets */
wire t_10205,  t_10206;
/* u2_3524 Output nets */
wire t_10207,  t_10208,  t_10209;
/* u2_3525 Output nets */
wire t_10210,  t_10211,  t_10212;
/* u2_3526 Output nets */
wire t_10213,  t_10214,  t_10215;
/* u0_3527 Output nets */
wire t_10216,  t_10217;
/* u2_3528 Output nets */
wire t_10218,  t_10219,  t_10220;
/* u2_3529 Output nets */
wire t_10221,  t_10222,  t_10223;
/* u2_3530 Output nets */
wire t_10224,  t_10225,  t_10226;
/* u1_3531 Output nets */
wire t_10227,  t_10228;
/* u2_3532 Output nets */
wire t_10229,  t_10230,  t_10231;
/* u2_3533 Output nets */
wire t_10232,  t_10233,  t_10234;
/* u2_3534 Output nets */
wire t_10235,  t_10236,  t_10237;
/* u0_3535 Output nets */
wire t_10238,  t_10239;
/* u2_3536 Output nets */
wire t_10240,  t_10241,  t_10242;
/* u2_3537 Output nets */
wire t_10243,  t_10244,  t_10245;
/* u2_3538 Output nets */
wire t_10246,  t_10247,  t_10248;
/* u0_3539 Output nets */
wire t_10249,  t_10250;
/* u2_3540 Output nets */
wire t_10251,  t_10252,  t_10253;
/* u2_3541 Output nets */
wire t_10254,  t_10255,  t_10256;
/* u2_3542 Output nets */
wire t_10257,  t_10258,  t_10259;
/* u0_3543 Output nets */
wire t_10260,  t_10261;
/* u2_3544 Output nets */
wire t_10262,  t_10263,  t_10264;
/* u2_3545 Output nets */
wire t_10265,  t_10266,  t_10267;
/* u2_3546 Output nets */
wire t_10268,  t_10269,  t_10270;
/* u0_3547 Output nets */
wire t_10271,  t_10272;
/* u2_3548 Output nets */
wire t_10273,  t_10274,  t_10275;
/* u2_3549 Output nets */
wire t_10276,  t_10277,  t_10278;
/* u2_3550 Output nets */
wire t_10279,  t_10280,  t_10281;
/* u1_3551 Output nets */
wire t_10282,  t_10283;
/* u2_3552 Output nets */
wire t_10284,  t_10285,  t_10286;
/* u2_3553 Output nets */
wire t_10287,  t_10288,  t_10289;
/* u2_3554 Output nets */
wire t_10290,  t_10291,  t_10292;
/* u1_3555 Output nets */
wire t_10293,  t_10294;
/* u2_3556 Output nets */
wire t_10295,  t_10296,  t_10297;
/* u2_3557 Output nets */
wire t_10298,  t_10299,  t_10300;
/* u2_3558 Output nets */
wire t_10301,  t_10302,  t_10303;
/* u1_3559 Output nets */
wire t_10304,  t_10305;
/* u2_3560 Output nets */
wire t_10306,  t_10307,  t_10308;
/* u2_3561 Output nets */
wire t_10309,  t_10310,  t_10311;
/* u2_3562 Output nets */
wire t_10312,  t_10313,  t_10314;
/* u1_3563 Output nets */
wire t_10315,  t_10316;
/* u2_3564 Output nets */
wire t_10317,  t_10318,  t_10319;
/* u2_3565 Output nets */
wire t_10320,  t_10321,  t_10322;
/* u2_3566 Output nets */
wire t_10323,  t_10324,  t_10325;
/* u1_3567 Output nets */
wire t_10326,  t_10327;
/* u2_3568 Output nets */
wire t_10328,  t_10329,  t_10330;
/* u2_3569 Output nets */
wire t_10331,  t_10332,  t_10333;
/* u2_3570 Output nets */
wire t_10334,  t_10335,  t_10336;
/* u1_3571 Output nets */
wire t_10337,  t_10338;
/* u2_3572 Output nets */
wire t_10339,  t_10340,  t_10341;
/* u2_3573 Output nets */
wire t_10342,  t_10343,  t_10344;
/* u2_3574 Output nets */
wire t_10345,  t_10346,  t_10347;
/* u1_3575 Output nets */
wire t_10348,  t_10349;
/* u2_3576 Output nets */
wire t_10350,  t_10351,  t_10352;
/* u2_3577 Output nets */
wire t_10353,  t_10354,  t_10355;
/* u2_3578 Output nets */
wire t_10356,  t_10357,  t_10358;
/* u1_3579 Output nets */
wire t_10359,  t_10360;
/* u2_3580 Output nets */
wire t_10361,  t_10362,  t_10363;
/* u2_3581 Output nets */
wire t_10364,  t_10365,  t_10366;
/* u2_3582 Output nets */
wire t_10367,  t_10368,  t_10369;
/* u1_3583 Output nets */
wire t_10370,  t_10371;
/* u2_3584 Output nets */
wire t_10372,  t_10373,  t_10374;
/* u2_3585 Output nets */
wire t_10375,  t_10376,  t_10377;
/* u2_3586 Output nets */
wire t_10378,  t_10379,  t_10380;
/* u2_3587 Output nets */
wire t_10381,  t_10382,  t_10383;
/* u2_3588 Output nets */
wire t_10384,  t_10385,  t_10386;
/* u2_3589 Output nets */
wire t_10387,  t_10388,  t_10389;
/* u2_3590 Output nets */
wire t_10390,  t_10391,  t_10392;
/* u2_3591 Output nets */
wire t_10393,  t_10394,  t_10395;
/* u2_3592 Output nets */
wire t_10396,  t_10397,  t_10398;
/* u2_3593 Output nets */
wire t_10399,  t_10400,  t_10401;
/* u2_3594 Output nets */
wire t_10402,  t_10403,  t_10404;
/* u2_3595 Output nets */
wire t_10405,  t_10406,  t_10407;
/* u2_3596 Output nets */
wire t_10408,  t_10409,  t_10410;
/* u2_3597 Output nets */
wire t_10411,  t_10412,  t_10413;
/* u2_3598 Output nets */
wire t_10414,  t_10415,  t_10416;
/* u2_3599 Output nets */
wire t_10417,  t_10418,  t_10419;
/* u2_3600 Output nets */
wire t_10420,  t_10421,  t_10422;
/* u2_3601 Output nets */
wire t_10423,  t_10424,  t_10425;
/* u2_3602 Output nets */
wire t_10426,  t_10427,  t_10428;
/* u2_3603 Output nets */
wire t_10429,  t_10430,  t_10431;
/* u2_3604 Output nets */
wire t_10432,  t_10433,  t_10434;
/* u2_3605 Output nets */
wire t_10435,  t_10436,  t_10437;
/* u2_3606 Output nets */
wire t_10438,  t_10439,  t_10440;
/* u2_3607 Output nets */
wire t_10441,  t_10442,  t_10443;
/* u2_3608 Output nets */
wire t_10444,  t_10445,  t_10446;
/* u2_3609 Output nets */
wire t_10447,  t_10448,  t_10449;
/* u2_3610 Output nets */
wire t_10450,  t_10451,  t_10452;
/* u2_3611 Output nets */
wire t_10453,  t_10454,  t_10455;
/* u2_3612 Output nets */
wire t_10456,  t_10457,  t_10458;
/* u2_3613 Output nets */
wire t_10459,  t_10460,  t_10461;
/* u2_3614 Output nets */
wire t_10462,  t_10463,  t_10464;
/* u2_3615 Output nets */
wire t_10465,  t_10466,  t_10467;
/* u2_3616 Output nets */
wire t_10468,  t_10469,  t_10470;
/* u2_3617 Output nets */
wire t_10471,  t_10472,  t_10473;
/* u2_3618 Output nets */
wire t_10474,  t_10475,  t_10476;
/* u2_3619 Output nets */
wire t_10477,  t_10478,  t_10479;
/* u2_3620 Output nets */
wire t_10480,  t_10481,  t_10482;
/* u2_3621 Output nets */
wire t_10483,  t_10484,  t_10485;
/* u2_3622 Output nets */
wire t_10486,  t_10487,  t_10488;
/* u2_3623 Output nets */
wire t_10489,  t_10490,  t_10491;
/* u2_3624 Output nets */
wire t_10492,  t_10493,  t_10494;
/* u2_3625 Output nets */
wire t_10495,  t_10496,  t_10497;
/* u2_3626 Output nets */
wire t_10498,  t_10499,  t_10500;
/* u2_3627 Output nets */
wire t_10501,  t_10502,  t_10503;
/* u2_3628 Output nets */
wire t_10504,  t_10505,  t_10506;
/* u2_3629 Output nets */
wire t_10507,  t_10508,  t_10509;
/* u2_3630 Output nets */
wire t_10510,  t_10511,  t_10512;
/* u2_3631 Output nets */
wire t_10513,  t_10514,  t_10515;
/* u2_3632 Output nets */
wire t_10516,  t_10517,  t_10518;
/* u2_3633 Output nets */
wire t_10519,  t_10520,  t_10521;
/* u2_3634 Output nets */
wire t_10522,  t_10523,  t_10524;
/* u2_3635 Output nets */
wire t_10525,  t_10526,  t_10527;
/* u2_3636 Output nets */
wire t_10528,  t_10529,  t_10530;
/* u2_3637 Output nets */
wire t_10531,  t_10532,  t_10533;
/* u2_3638 Output nets */
wire t_10534,  t_10535,  t_10536;
/* u2_3639 Output nets */
wire t_10537,  t_10538,  t_10539;
/* u2_3640 Output nets */
wire t_10540,  t_10541,  t_10542;
/* u2_3641 Output nets */
wire t_10543,  t_10544,  t_10545;
/* u2_3642 Output nets */
wire t_10546,  t_10547,  t_10548;
/* u2_3643 Output nets */
wire t_10549,  t_10550,  t_10551;
/* u2_3644 Output nets */
wire t_10552,  t_10553,  t_10554;
/* u2_3645 Output nets */
wire t_10555,  t_10556,  t_10557;
/* u2_3646 Output nets */
wire t_10558,  t_10559,  t_10560;
/* u2_3647 Output nets */
wire t_10561,  t_10562,  t_10563;
/* u2_3648 Output nets */
wire t_10564,  t_10565,  t_10566;
/* u2_3649 Output nets */
wire t_10567,  t_10568,  t_10569;
/* u2_3650 Output nets */
wire t_10570,  t_10571,  t_10572;
/* u2_3651 Output nets */
wire t_10573,  t_10574,  t_10575;
/* u2_3652 Output nets */
wire t_10576,  t_10577,  t_10578;
/* u2_3653 Output nets */
wire t_10579,  t_10580,  t_10581;
/* u2_3654 Output nets */
wire t_10582,  t_10583,  t_10584;
/* u2_3655 Output nets */
wire t_10585,  t_10586,  t_10587;
/* u2_3656 Output nets */
wire t_10588,  t_10589,  t_10590;
/* u2_3657 Output nets */
wire t_10591,  t_10592,  t_10593;
/* u2_3658 Output nets */
wire t_10594,  t_10595,  t_10596;
/* u2_3659 Output nets */
wire t_10597,  t_10598,  t_10599;
/* u2_3660 Output nets */
wire t_10600,  t_10601,  t_10602;
/* u2_3661 Output nets */
wire t_10603,  t_10604,  t_10605;
/* u2_3662 Output nets */
wire t_10606,  t_10607,  t_10608;
/* u2_3663 Output nets */
wire t_10609,  t_10610,  t_10611;
/* u2_3664 Output nets */
wire t_10612,  t_10613,  t_10614;
/* u2_3665 Output nets */
wire t_10615,  t_10616,  t_10617;
/* u2_3666 Output nets */
wire t_10618,  t_10619,  t_10620;
/* u2_3667 Output nets */
wire t_10621,  t_10622,  t_10623;
/* u2_3668 Output nets */
wire t_10624,  t_10625,  t_10626;
/* u2_3669 Output nets */
wire t_10627,  t_10628,  t_10629;
/* u2_3670 Output nets */
wire t_10630,  t_10631,  t_10632;
/* u2_3671 Output nets */
wire t_10633,  t_10634,  t_10635;
/* u2_3672 Output nets */
wire t_10636,  t_10637,  t_10638;
/* u2_3673 Output nets */
wire t_10639,  t_10640,  t_10641;
/* u2_3674 Output nets */
wire t_10642,  t_10643,  t_10644;
/* u2_3675 Output nets */
wire t_10645,  t_10646,  t_10647;
/* u2_3676 Output nets */
wire t_10648,  t_10649,  t_10650;
/* u2_3677 Output nets */
wire t_10651,  t_10652,  t_10653;
/* u2_3678 Output nets */
wire t_10654,  t_10655,  t_10656;
/* u2_3679 Output nets */
wire t_10657,  t_10658,  t_10659;
/* u2_3680 Output nets */
wire t_10660,  t_10661,  t_10662;
/* u2_3681 Output nets */
wire t_10663,  t_10664,  t_10665;
/* u2_3682 Output nets */
wire t_10666,  t_10667,  t_10668;
/* u2_3683 Output nets */
wire t_10669,  t_10670,  t_10671;
/* u2_3684 Output nets */
wire t_10672,  t_10673,  t_10674;
/* u2_3685 Output nets */
wire t_10675,  t_10676,  t_10677;
/* u2_3686 Output nets */
wire t_10678,  t_10679,  t_10680;
/* u1_3687 Output nets */
wire t_10681,  t_10682;
/* u2_3688 Output nets */
wire t_10683,  t_10684,  t_10685;
/* u2_3689 Output nets */
wire t_10686,  t_10687,  t_10688;
/* u2_3690 Output nets */
wire t_10689,  t_10690,  t_10691;
/* u0_3691 Output nets */
wire t_10692,  t_10693;
/* u2_3692 Output nets */
wire t_10694,  t_10695,  t_10696;
/* u2_3693 Output nets */
wire t_10697,  t_10698,  t_10699;
/* u2_3694 Output nets */
wire t_10700,  t_10701,  t_10702;
/* u1_3695 Output nets */
wire t_10703,  t_10704;
/* u2_3696 Output nets */
wire t_10705,  t_10706,  t_10707;
/* u2_3697 Output nets */
wire t_10708,  t_10709,  t_10710;
/* u2_3698 Output nets */
wire t_10711,  t_10712,  t_10713;
/* u0_3699 Output nets */
wire t_10714,  t_10715;
/* u2_3700 Output nets */
wire t_10716,  t_10717,  t_10718;
/* u2_3701 Output nets */
wire t_10719,  t_10720,  t_10721;
/* u2_3702 Output nets */
wire t_10722,  t_10723,  t_10724;
/* u0_3703 Output nets */
wire t_10725,  t_10726;
/* u2_3704 Output nets */
wire t_10727,  t_10728,  t_10729;
/* u2_3705 Output nets */
wire t_10730,  t_10731,  t_10732;
/* u2_3706 Output nets */
wire t_10733,  t_10734,  t_10735;
/* u0_3707 Output nets */
wire t_10736,  t_10737;
/* u2_3708 Output nets */
wire t_10738,  t_10739,  t_10740;
/* u2_3709 Output nets */
wire t_10741,  t_10742,  t_10743;
/* u2_3710 Output nets */
wire t_10744,  t_10745,  t_10746;
/* u0_3711 Output nets */
wire t_10747,  t_10748;
/* u2_3712 Output nets */
wire t_10749,  t_10750,  t_10751;
/* u2_3713 Output nets */
wire t_10752,  t_10753,  t_10754;
/* u2_3714 Output nets */
wire t_10755,  t_10756,  t_10757;
/* u1_3715 Output nets */
wire t_10758,  t_10759;
/* u2_3716 Output nets */
wire t_10760,  t_10761,  t_10762;
/* u2_3717 Output nets */
wire t_10763,  t_10764,  t_10765;
/* u2_3718 Output nets */
wire t_10766,  t_10767,  t_10768;
/* u0_3719 Output nets */
wire t_10769,  t_10770;
/* u2_3720 Output nets */
wire t_10771,  t_10772,  t_10773;
/* u2_3721 Output nets */
wire t_10774,  t_10775,  t_10776;
/* u2_3722 Output nets */
wire t_10777,  t_10778,  t_10779;
/* u0_3723 Output nets */
wire t_10780,  t_10781;
/* u2_3724 Output nets */
wire t_10782,  t_10783,  t_10784;
/* u2_3725 Output nets */
wire t_10785,  t_10786,  t_10787;
/* u2_3726 Output nets */
wire t_10788,  t_10789,  t_10790;
/* u0_3727 Output nets */
wire t_10791,  t_10792;
/* u2_3728 Output nets */
wire t_10793,  t_10794,  t_10795;
/* u2_3729 Output nets */
wire t_10796,  t_10797,  t_10798;
/* u2_3730 Output nets */
wire t_10799,  t_10800,  t_10801;
/* u0_3731 Output nets */
wire t_10802,  t_10803;
/* u2_3732 Output nets */
wire t_10804,  t_10805,  t_10806;
/* u2_3733 Output nets */
wire t_10807,  t_10808,  t_10809;
/* u2_3734 Output nets */
wire t_10810,  t_10811,  t_10812;
/* u0_3735 Output nets */
wire t_10813,  t_10814;
/* u2_3736 Output nets */
wire t_10815,  t_10816,  t_10817;
/* u2_3737 Output nets */
wire t_10818,  t_10819,  t_10820;
/* u2_3738 Output nets */
wire t_10821,  t_10822,  t_10823;
/* u0_3739 Output nets */
wire t_10824,  t_10825;
/* u2_3740 Output nets */
wire t_10826,  t_10827,  t_10828;
/* u2_3741 Output nets */
wire t_10829,  t_10830,  t_10831;
/* u2_3742 Output nets */
wire t_10832,  t_10833,  t_10834;
/* u0_3743 Output nets */
wire t_10835,  t_10836;
/* u2_3744 Output nets */
wire t_10837,  t_10838,  t_10839;
/* u2_3745 Output nets */
wire t_10840,  t_10841,  t_10842;
/* u2_3746 Output nets */
wire t_10843,  t_10844,  t_10845;
/* u0_3747 Output nets */
wire t_10846,  t_10847;
/* u2_3748 Output nets */
wire t_10848,  t_10849,  t_10850;
/* u2_3749 Output nets */
wire t_10851,  t_10852,  t_10853;
/* u2_3750 Output nets */
wire t_10854,  t_10855,  t_10856;
/* u2_3751 Output nets */
wire t_10857,  t_10858,  t_10859;
/* u2_3752 Output nets */
wire t_10860,  t_10861,  t_10862;
/* u2_3753 Output nets */
wire t_10863,  t_10864,  t_10865;
/* u2_3754 Output nets */
wire t_10866,  t_10867,  t_10868;
/* u2_3755 Output nets */
wire t_10869,  t_10870,  t_10871;
/* u2_3756 Output nets */
wire t_10872,  t_10873,  t_10874;
/* u2_3757 Output nets */
wire t_10875,  t_10876,  t_10877;
/* u2_3758 Output nets */
wire t_10878,  t_10879,  t_10880;
/* u2_3759 Output nets */
wire t_10881,  t_10882,  t_10883;
/* u2_3760 Output nets */
wire t_10884,  t_10885,  t_10886;
/* u2_3761 Output nets */
wire t_10887,  t_10888,  t_10889;
/* u2_3762 Output nets */
wire t_10890,  t_10891,  t_10892;
/* u2_3763 Output nets */
wire t_10893,  t_10894,  t_10895;
/* u2_3764 Output nets */
wire t_10896,  t_10897,  t_10898;
/* u2_3765 Output nets */
wire t_10899,  t_10900,  t_10901;
/* u2_3766 Output nets */
wire t_10902,  t_10903,  t_10904;
/* u2_3767 Output nets */
wire t_10905,  t_10906,  t_10907;
/* u2_3768 Output nets */
wire t_10908,  t_10909,  t_10910;
/* u2_3769 Output nets */
wire t_10911,  t_10912,  t_10913;
/* u2_3770 Output nets */
wire t_10914,  t_10915,  t_10916;
/* u2_3771 Output nets */
wire t_10917,  t_10918,  t_10919;
/* u2_3772 Output nets */
wire t_10920,  t_10921,  t_10922;
/* u2_3773 Output nets */
wire t_10923,  t_10924,  t_10925;
/* u2_3774 Output nets */
wire t_10926,  t_10927,  t_10928;
/* u2_3775 Output nets */
wire t_10929,  t_10930,  t_10931;
/* u2_3776 Output nets */
wire t_10932,  t_10933,  t_10934;
/* u2_3777 Output nets */
wire t_10935,  t_10936,  t_10937;
/* u2_3778 Output nets */
wire t_10938,  t_10939,  t_10940;
/* u2_3779 Output nets */
wire t_10941,  t_10942,  t_10943;
/* u2_3780 Output nets */
wire t_10944,  t_10945,  t_10946;
/* u2_3781 Output nets */
wire t_10947,  t_10948,  t_10949;
/* u2_3782 Output nets */
wire t_10950,  t_10951,  t_10952;
/* u2_3783 Output nets */
wire t_10953,  t_10954,  t_10955;
/* u2_3784 Output nets */
wire t_10956,  t_10957,  t_10958;
/* u2_3785 Output nets */
wire t_10959,  t_10960,  t_10961;
/* u2_3786 Output nets */
wire t_10962,  t_10963,  t_10964;
/* u2_3787 Output nets */
wire t_10965,  t_10966,  t_10967;
/* u2_3788 Output nets */
wire t_10968,  t_10969,  t_10970;
/* u2_3789 Output nets */
wire t_10971,  t_10972,  t_10973;
/* u2_3790 Output nets */
wire t_10974,  t_10975,  t_10976;
/* u2_3791 Output nets */
wire t_10977,  t_10978,  t_10979;
/* u2_3792 Output nets */
wire t_10980,  t_10981,  t_10982;
/* u2_3793 Output nets */
wire t_10983,  t_10984,  t_10985;
/* u2_3794 Output nets */
wire t_10986,  t_10987,  t_10988;
/* u2_3795 Output nets */
wire t_10989,  t_10990,  t_10991;
/* u2_3796 Output nets */
wire t_10992,  t_10993,  t_10994;
/* u2_3797 Output nets */
wire t_10995,  t_10996,  t_10997;
/* u1_3798 Output nets */
wire t_10998,  t_10999;
/* u2_3799 Output nets */
wire t_11000,  t_11001,  t_11002;
/* u2_3800 Output nets */
wire t_11003,  t_11004,  t_11005;
/* u0_3801 Output nets */
wire t_11006,  t_11007;
/* u2_3802 Output nets */
wire t_11008,  t_11009,  t_11010;
/* u2_3803 Output nets */
wire t_11011,  t_11012,  t_11013;
/* u1_3804 Output nets */
wire t_11014,  t_11015;
/* u2_3805 Output nets */
wire t_11016,  t_11017,  t_11018;
/* u2_3806 Output nets */
wire t_11019,  t_11020,  t_11021;
/* u0_3807 Output nets */
wire t_11022,  t_11023;
/* u2_3808 Output nets */
wire t_11024,  t_11025,  t_11026;
/* u2_3809 Output nets */
wire t_11027,  t_11028,  t_11029;
/* u0_3810 Output nets */
wire t_11030,  t_11031;
/* u2_3811 Output nets */
wire t_11032,  t_11033,  t_11034;
/* u2_3812 Output nets */
wire t_11035,  t_11036,  t_11037;
/* u0_3813 Output nets */
wire t_11038,  t_11039;
/* u2_3814 Output nets */
wire t_11040,  t_11041,  t_11042;
/* u2_3815 Output nets */
wire t_11043,  t_11044,  t_11045;
/* u0_3816 Output nets */
wire t_11046,  t_11047;
/* u2_3817 Output nets */
wire t_11048,  t_11049,  t_11050;
/* u2_3818 Output nets */
wire t_11051,  t_11052,  t_11053;
/* u1_3819 Output nets */
wire t_11054,  t_11055;
/* u2_3820 Output nets */
wire t_11056,  t_11057,  t_11058;
/* u2_3821 Output nets */
wire t_11059,  t_11060,  t_11061;
/* u0_3822 Output nets */
wire t_11062,  t_11063;
/* u2_3823 Output nets */
wire t_11064,  t_11065,  t_11066;
/* u2_3824 Output nets */
wire t_11067,  t_11068,  t_11069;
/* u0_3825 Output nets */
wire t_11070,  t_11071;
/* u2_3826 Output nets */
wire t_11072,  t_11073,  t_11074;
/* u2_3827 Output nets */
wire t_11075,  t_11076,  t_11077;
/* u0_3828 Output nets */
wire t_11078,  t_11079;
/* u2_3829 Output nets */
wire t_11080,  t_11081,  t_11082;
/* u2_3830 Output nets */
wire t_11083,  t_11084,  t_11085;
/* u0_3831 Output nets */
wire t_11086,  t_11087;
/* u2_3832 Output nets */
wire t_11088,  t_11089,  t_11090;
/* u2_3833 Output nets */
wire t_11091,  t_11092,  t_11093;
/* u0_3834 Output nets */
wire t_11094,  t_11095;
/* u2_3835 Output nets */
wire t_11096,  t_11097,  t_11098;
/* u2_3836 Output nets */
wire t_11099,  t_11100,  t_11101;
/* u0_3837 Output nets */
wire t_11102,  t_11103;
/* u2_3838 Output nets */
wire t_11104,  t_11105,  t_11106;
/* u2_3839 Output nets */
wire t_11107,  t_11108,  t_11109;
/* u0_3840 Output nets */
wire t_11110,  t_11111;
/* u2_3841 Output nets */
wire t_11112,  t_11113,  t_11114;
/* u2_3842 Output nets */
wire t_11115,  t_11116,  t_11117;
/* u0_3843 Output nets */
wire t_11118,  t_11119;
/* u2_3844 Output nets */
wire t_11120,  t_11121,  t_11122;
/* u2_3845 Output nets */
wire t_11123,  t_11124,  t_11125;
/* u2_3846 Output nets */
wire t_11126,  t_11127,  t_11128;
/* u2_3847 Output nets */
wire t_11129,  t_11130,  t_11131;
/* u2_3848 Output nets */
wire t_11132,  t_11133,  t_11134;
/* u2_3849 Output nets */
wire t_11135,  t_11136,  t_11137;
/* u2_3850 Output nets */
wire t_11138,  t_11139,  t_11140;
/* u2_3851 Output nets */
wire t_11141,  t_11142,  t_11143;
/* u2_3852 Output nets */
wire t_11144,  t_11145,  t_11146;
/* u2_3853 Output nets */
wire t_11147,  t_11148,  t_11149;
/* u2_3854 Output nets */
wire t_11150,  t_11151,  t_11152;
/* u2_3855 Output nets */
wire t_11153,  t_11154,  t_11155;
/* u2_3856 Output nets */
wire t_11156,  t_11157,  t_11158;
/* u2_3857 Output nets */
wire t_11159,  t_11160,  t_11161;
/* u2_3858 Output nets */
wire t_11162,  t_11163,  t_11164;
/* u2_3859 Output nets */
wire t_11165,  t_11166,  t_11167;
/* u2_3860 Output nets */
wire t_11168,  t_11169,  t_11170;
/* u2_3861 Output nets */
wire t_11171,  t_11172,  t_11173;
/* u2_3862 Output nets */
wire t_11174,  t_11175,  t_11176;
/* u2_3863 Output nets */
wire t_11177,  t_11178,  t_11179;
/* u2_3864 Output nets */
wire t_11180,  t_11181,  t_11182;
/* u2_3865 Output nets */
wire t_11183,  t_11184,  t_11185;
/* u2_3866 Output nets */
wire t_11186,  t_11187,  t_11188;
/* u2_3867 Output nets */
wire t_11189,  t_11190,  t_11191;
/* u2_3868 Output nets */
wire t_11192,  t_11193,  t_11194;
/* u2_3869 Output nets */
wire t_11195,  t_11196,  t_11197;
/* u2_3870 Output nets */
wire t_11198,  t_11199,  t_11200;
/* u2_3871 Output nets */
wire t_11201,  t_11202,  t_11203;
/* u2_3872 Output nets */
wire t_11204,  t_11205,  t_11206;
/* u2_3873 Output nets */
wire t_11207,  t_11208,  t_11209;
/* u2_3874 Output nets */
wire t_11210,  t_11211,  t_11212;
/* u2_3875 Output nets */
wire t_11213,  t_11214,  t_11215;
/* u2_3876 Output nets */
wire t_11216,  t_11217,  t_11218;
/* u1_3877 Output nets */
wire t_11219,  t_11220;
/* u2_3878 Output nets */
wire t_11221,  t_11222,  t_11223;
/* u0_3879 Output nets */
wire t_11224,  t_11225;
/* u2_3880 Output nets */
wire t_11226,  t_11227,  t_11228;
/* u1_3881 Output nets */
wire t_11229,  t_11230;
/* u2_3882 Output nets */
wire t_11231,  t_11232,  t_11233;
/* u0_3883 Output nets */
wire t_11234,  t_11235;
/* u2_3884 Output nets */
wire t_11236,  t_11237,  t_11238;
/* u0_3885 Output nets */
wire t_11239,  t_11240;
/* u2_3886 Output nets */
wire t_11241,  t_11242,  t_11243;
/* u0_3887 Output nets */
wire t_11244,  t_11245;
/* u2_3888 Output nets */
wire t_11246,  t_11247,  t_11248;
/* u0_3889 Output nets */
wire t_11249,  t_11250;
/* u2_3890 Output nets */
wire t_11251,  t_11252,  t_11253;
/* u1_3891 Output nets */
wire t_11254,  t_11255;
/* u2_3892 Output nets */
wire t_11256,  t_11257,  t_11258;
/* u0_3893 Output nets */
wire t_11259,  t_11260;
/* u2_3894 Output nets */
wire t_11261,  t_11262,  t_11263;
/* u0_3895 Output nets */
wire t_11264,  t_11265;
/* u2_3896 Output nets */
wire t_11266,  t_11267,  t_11268;
/* u0_3897 Output nets */
wire t_11269,  t_11270;
/* u2_3898 Output nets */
wire t_11271,  t_11272,  t_11273;
/* u0_3899 Output nets */
wire t_11274,  t_11275;
/* u2_3900 Output nets */
wire t_11276,  t_11277,  t_11278;
/* u0_3901 Output nets */
wire t_11279,  t_11280;
/* u2_3902 Output nets */
wire t_11281,  t_11282,  t_11283;
/* u0_3903 Output nets */
wire t_11284,  t_11285;
/* u2_3904 Output nets */
wire t_11286,  t_11287,  t_11288;
/* u0_3905 Output nets */
wire t_11289,  t_11290;
/* u2_3906 Output nets */
wire t_11291,  t_11292,  t_11293;
/* u0_3907 Output nets */
wire t_11294,  t_11295;
/* u2_3908 Output nets */
wire t_11296,  t_11297,  t_11298;
/* u2_3909 Output nets */
wire t_11299,  t_11300,  t_11301;
/* u2_3910 Output nets */
wire t_11302,  t_11303,  t_11304;
/* u2_3911 Output nets */
wire t_11305,  t_11306,  t_11307;
/* u2_3912 Output nets */
wire t_11308,  t_11309,  t_11310;
/* u2_3913 Output nets */
wire t_11311,  t_11312,  t_11313;
/* u2_3914 Output nets */
wire t_11314,  t_11315,  t_11316;
/* u2_3915 Output nets */
wire t_11317,  t_11318,  t_11319;
/* u2_3916 Output nets */
wire t_11320,  t_11321,  t_11322;
/* u2_3917 Output nets */
wire t_11323,  t_11324,  t_11325;
/* u2_3918 Output nets */
wire t_11326,  t_11327,  t_11328;
/* u2_3919 Output nets */
wire t_11329,  t_11330,  t_11331;
/* u2_3920 Output nets */
wire t_11332,  t_11333,  t_11334;
/* u2_3921 Output nets */
wire t_11335,  t_11336,  t_11337;
/* u2_3922 Output nets */
wire t_11338,  t_11339,  t_11340;
/* u2_3923 Output nets */
wire t_11341,  t_11342,  t_11343;
/* u1_3924 Output nets */
wire t_11344,  t_11345;
/* u0_3925 Output nets */
wire t_11346,  t_11347;
/* u1_3926 Output nets */
wire t_11348,  t_11349;
/* u0_3927 Output nets */
wire t_11350,  t_11351;
/* u0_3928 Output nets */
wire t_11352,  t_11353;
/* u0_3929 Output nets */
wire t_11354,  t_11355;
/* u0_3930 Output nets */
wire t_11356,  t_11357;
/* u1_3931 Output nets */
wire t_11358,  t_11359;
/* u0_3932 Output nets */
wire t_11360,  t_11361;
/* u0_3933 Output nets */
wire t_11362,  t_11363;
/* u0_3934 Output nets */
wire t_11364,  t_11365;
/* u0_3935 Output nets */
wire t_11366,  t_11367;
/* u0_3936 Output nets */
wire t_11368,  t_11369;
/* u0_3937 Output nets */
wire t_11370;

/* compress stage 3 */
half_adder u0_3304(.a(t_6336), .b(t_2), .o(t_9620), .cout(t_9621));
half_adder u0_3305(.a(t_6339), .b(t_6338), .o(t_9622), .cout(t_9623));
half_adder u0_3306(.a(t_6341), .b(t_6340), .o(t_9624), .cout(t_9625));
half_adder u0_3307(.a(t_6343), .b(t_6342), .o(t_9626), .cout(t_9627));
half_adder u0_3308(.a(t_6345), .b(t_6344), .o(t_9628), .cout(t_9629));
half_adder u0_3309(.a(t_6347), .b(t_6346), .o(t_9630), .cout(t_9631));
compressor_3_2 u1_3310(.a(t_6349), .b(t_6348), .cin(t_21), .o(t_9632), .cout(t_9633));
half_adder u0_3311(.a(t_6351), .b(t_6350), .o(t_9634), .cout(t_9635));
compressor_3_2 u1_3312(.a(t_6353), .b(t_6352), .cin(t_32), .o(t_9636), .cout(t_9637));
half_adder u0_3313(.a(t_6355), .b(t_6354), .o(t_9638), .cout(t_9639));
half_adder u0_3314(.a(t_6358), .b(t_6356), .o(t_9640), .cout(t_9641));
half_adder u0_3315(.a(t_6361), .b(t_6359), .o(t_9642), .cout(t_9643));
half_adder u0_3316(.a(t_6364), .b(t_6362), .o(t_9644), .cout(t_9645));
compressor_3_2 u1_3317(.a(t_6367), .b(t_6365), .cin(t_62), .o(t_9646), .cout(t_9647));
compressor_3_2 u1_3318(.a(t_6373), .b(t_6370), .cin(t_6368), .o(t_9648), .cout(t_9649));
compressor_3_2 u1_3319(.a(t_6374), .b(t_6371), .cin(t_76), .o(t_9650), .cout(t_9651));
compressor_3_2 u1_3320(.a(t_6381), .b(t_6378), .cin(t_6376), .o(t_9652), .cout(t_9653));
compressor_3_2 u1_3321(.a(t_6383), .b(t_6382), .cin(t_6379), .o(t_9654), .cout(t_9655));
compressor_3_2 u1_3322(.a(t_6388), .b(t_6387), .cin(t_6384), .o(t_9656), .cout(t_9657));
compressor_3_2 u1_3323(.a(t_6393), .b(t_6392), .cin(t_6389), .o(t_9658), .cout(t_9659));
compressor_3_2 u1_3324(.a(t_6398), .b(t_6397), .cin(t_6394), .o(t_9660), .cout(t_9661));
compressor_3_2 u1_3325(.a(t_6403), .b(t_6402), .cin(t_6399), .o(t_9662), .cout(t_9663));
compressor_4_2 u2_3326(.a(t_6411), .b(t_6408), .c(t_6407), .d(t_6404), .cin(t_137), .o(t_9664), .co(t_9665), .cout(t_9666));
compressor_4_2 u2_3327(.a(t_6416), .b(t_6413), .c(t_6412), .d(t_6409), .cin(t_9666), .o(t_9667), .co(t_9668), .cout(t_9669));
compressor_4_2 u2_3328(.a(t_6418), .b(t_6417), .c(t_6414), .d(t_160), .cin(t_9669), .o(t_9670), .co(t_9671), .cout(t_9672));
compressor_4_2 u2_3329(.a(t_6426), .b(t_6423), .c(t_6422), .d(t_6419), .cin(t_9672), .o(t_9673), .co(t_9674), .cout(t_9675));
compressor_4_2 u2_3330(.a(t_6432), .b(t_6429), .c(t_6427), .d(t_6424), .cin(t_9675), .o(t_9676), .co(t_9677), .cout(t_9678));
compressor_4_2 u2_3331(.a(t_6438), .b(t_6435), .c(t_6433), .d(t_6430), .cin(t_9678), .o(t_9679), .co(t_9680), .cout(t_9681));
compressor_4_2 u2_3332(.a(t_6444), .b(t_6441), .c(t_6439), .d(t_6436), .cin(t_9681), .o(t_9682), .co(t_9683), .cout(t_9684));
compressor_4_2 u2_3333(.a(t_6447), .b(t_6445), .c(t_6442), .d(t_220), .cin(t_9684), .o(t_9685), .co(t_9686), .cout(t_9687));
compressor_4_2 u2_3334(.a(t_6456), .b(t_6453), .c(t_6451), .d(t_6448), .cin(t_9687), .o(t_9688), .co(t_9689), .cout(t_9690));
compressor_4_2 u2_3335(.a(t_6460), .b(t_6457), .c(t_6454), .d(t_246), .cin(t_9690), .o(t_9691), .co(t_9692), .cout(t_9693));
half_adder u0_3336(.a(t_6464), .b(t_6461), .o(t_9694), .cout(t_9695));
compressor_4_2 u2_3337(.a(t_6470), .b(t_6467), .c(t_6465), .d(t_6462), .cin(t_9693), .o(t_9696), .co(t_9697), .cout(t_9698));
compressor_4_2 u2_3338(.a(t_6475), .b(t_6474), .c(t_6471), .d(t_6468), .cin(t_9698), .o(t_9699), .co(t_9700), .cout(t_9701));
half_adder u0_3339(.a(t_6481), .b(t_6478), .o(t_9702), .cout(t_9703));
compressor_4_2 u2_3340(.a(t_6483), .b(t_6482), .c(t_6479), .d(t_6476), .cin(t_9701), .o(t_9704), .co(t_9705), .cout(t_9706));
half_adder u0_3341(.a(t_6489), .b(t_6486), .o(t_9707), .cout(t_9708));
compressor_4_2 u2_3342(.a(t_6491), .b(t_6490), .c(t_6487), .d(t_6484), .cin(t_9706), .o(t_9709), .co(t_9710), .cout(t_9711));
half_adder u0_3343(.a(t_6497), .b(t_6494), .o(t_9712), .cout(t_9713));
compressor_4_2 u2_3344(.a(t_6499), .b(t_6498), .c(t_6495), .d(t_6492), .cin(t_9711), .o(t_9714), .co(t_9715), .cout(t_9716));
half_adder u0_3345(.a(t_6505), .b(t_6502), .o(t_9717), .cout(t_9718));
compressor_4_2 u2_3346(.a(t_6507), .b(t_6506), .c(t_6503), .d(t_6500), .cin(t_9716), .o(t_9719), .co(t_9720), .cout(t_9721));
half_adder u0_3347(.a(t_6513), .b(t_6510), .o(t_9722), .cout(t_9723));
compressor_4_2 u2_3348(.a(t_6514), .b(t_6511), .c(t_6508), .d(t_349), .cin(t_9721), .o(t_9724), .co(t_9725), .cout(t_9726));
compressor_3_2 u1_3349(.a(t_6521), .b(t_6518), .cin(t_6515), .o(t_9727), .cout(t_9728));
compressor_4_2 u2_3350(.a(t_6523), .b(t_6522), .c(t_6519), .d(t_6516), .cin(t_9726), .o(t_9729), .co(t_9730), .cout(t_9731));
half_adder u0_3351(.a(t_6529), .b(t_6526), .o(t_9732), .cout(t_9733));
compressor_4_2 u2_3352(.a(t_6530), .b(t_6527), .c(t_6524), .d(t_384), .cin(t_9731), .o(t_9734), .co(t_9735), .cout(t_9736));
compressor_3_2 u1_3353(.a(t_6537), .b(t_6534), .cin(t_6531), .o(t_9737), .cout(t_9738));
compressor_4_2 u2_3354(.a(t_6539), .b(t_6538), .c(t_6535), .d(t_6532), .cin(t_9736), .o(t_9739), .co(t_9740), .cout(t_9741));
half_adder u0_3355(.a(t_6545), .b(t_6542), .o(t_9742), .cout(t_9743));
compressor_4_2 u2_3356(.a(t_6548), .b(t_6546), .c(t_6543), .d(t_6540), .cin(t_9741), .o(t_9744), .co(t_9745), .cout(t_9746));
half_adder u0_3357(.a(t_6554), .b(t_6551), .o(t_9747), .cout(t_9748));
compressor_4_2 u2_3358(.a(t_6557), .b(t_6555), .c(t_6552), .d(t_6549), .cin(t_9746), .o(t_9749), .co(t_9750), .cout(t_9751));
half_adder u0_3359(.a(t_6563), .b(t_6560), .o(t_9752), .cout(t_9753));
compressor_4_2 u2_3360(.a(t_6566), .b(t_6564), .c(t_6561), .d(t_6558), .cin(t_9751), .o(t_9754), .co(t_9755), .cout(t_9756));
half_adder u0_3361(.a(t_6572), .b(t_6569), .o(t_9757), .cout(t_9758));
compressor_4_2 u2_3362(.a(t_6573), .b(t_6570), .c(t_6567), .d(t_474), .cin(t_9756), .o(t_9759), .co(t_9760), .cout(t_9761));
compressor_3_2 u1_3363(.a(t_6581), .b(t_6578), .cin(t_6575), .o(t_9762), .cout(t_9763));
compressor_4_2 u2_3364(.a(t_6584), .b(t_6582), .c(t_6579), .d(t_6576), .cin(t_9761), .o(t_9764), .co(t_9765), .cout(t_9766));
compressor_3_2 u1_3365(.a(t_6593), .b(t_6590), .cin(t_6587), .o(t_9767), .cout(t_9768));
compressor_4_2 u2_3366(.a(t_6591), .b(t_6588), .c(t_6585), .d(t_512), .cin(t_9766), .o(t_9769), .co(t_9770), .cout(t_9771));
compressor_3_2 u1_3367(.a(t_6598), .b(t_6595), .cin(t_6594), .o(t_9772), .cout(t_9773));
compressor_4_2 u2_3368(.a(t_6604), .b(t_6602), .c(t_6599), .d(t_6596), .cin(t_9771), .o(t_9774), .co(t_9775), .cout(t_9776));
compressor_3_2 u1_3369(.a(t_6613), .b(t_6610), .cin(t_6607), .o(t_9777), .cout(t_9778));
compressor_4_2 u2_3370(.a(t_6614), .b(t_6611), .c(t_6608), .d(t_6605), .cin(t_9776), .o(t_9779), .co(t_9780), .cout(t_9781));
compressor_3_2 u1_3371(.a(t_6621), .b(t_6618), .cin(t_6615), .o(t_9782), .cout(t_9783));
compressor_4_2 u2_3372(.a(t_6625), .b(t_6622), .c(t_6619), .d(t_6616), .cin(t_9781), .o(t_9784), .co(t_9785), .cout(t_9786));
compressor_3_2 u1_3373(.a(t_6632), .b(t_6629), .cin(t_6626), .o(t_9787), .cout(t_9788));
compressor_4_2 u2_3374(.a(t_6636), .b(t_6633), .c(t_6630), .d(t_6627), .cin(t_9786), .o(t_9789), .co(t_9790), .cout(t_9791));
compressor_3_2 u1_3375(.a(t_6643), .b(t_6640), .cin(t_6637), .o(t_9792), .cout(t_9793));
compressor_4_2 u2_3376(.a(t_6647), .b(t_6644), .c(t_6641), .d(t_6638), .cin(t_9791), .o(t_9794), .co(t_9795), .cout(t_9796));
compressor_3_2 u1_3377(.a(t_6654), .b(t_6651), .cin(t_6648), .o(t_9797), .cout(t_9798));
compressor_4_2 u2_3378(.a(t_6658), .b(t_6655), .c(t_6652), .d(t_6649), .cin(t_9796), .o(t_9799), .co(t_9800), .cout(t_9801));
compressor_3_2 u1_3379(.a(t_6665), .b(t_6662), .cin(t_6659), .o(t_9802), .cout(t_9803));
compressor_4_2 u2_3380(.a(t_6666), .b(t_6663), .c(t_6660), .d(t_657), .cin(t_9801), .o(t_9804), .co(t_9805), .cout(t_9806));
compressor_4_2 u2_3381(.a(t_6679), .b(t_6676), .c(t_6673), .d(t_6670), .cin(t_6669), .o(t_9807), .co(t_9808), .cout(t_9809));
compressor_4_2 u2_3382(.a(t_6680), .b(t_6677), .c(t_6674), .d(t_6671), .cin(t_9806), .o(t_9810), .co(t_9811), .cout(t_9812));
compressor_4_2 u2_3383(.a(t_6690), .b(t_6687), .c(t_6684), .d(t_6681), .cin(t_9809), .o(t_9813), .co(t_9814), .cout(t_9815));
compressor_4_2 u2_3384(.a(t_6688), .b(t_6685), .c(t_6682), .d(t_704), .cin(t_9812), .o(t_9816), .co(t_9817), .cout(t_9818));
compressor_4_2 u2_3385(.a(t_6698), .b(t_6695), .c(t_6692), .d(t_6691), .cin(t_9815), .o(t_9819), .co(t_9820), .cout(t_9821));
compressor_4_2 u2_3386(.a(t_6702), .b(t_6699), .c(t_6696), .d(t_6693), .cin(t_9818), .o(t_9822), .co(t_9823), .cout(t_9824));
compressor_4_2 u2_3387(.a(t_6712), .b(t_6709), .c(t_6706), .d(t_6703), .cin(t_9821), .o(t_9825), .co(t_9826), .cout(t_9827));
compressor_4_2 u2_3388(.a(t_6713), .b(t_6710), .c(t_6707), .d(t_6704), .cin(t_9824), .o(t_9828), .co(t_9829), .cout(t_9830));
compressor_4_2 u2_3389(.a(t_6724), .b(t_6721), .c(t_6718), .d(t_6715), .cin(t_9827), .o(t_9831), .co(t_9832), .cout(t_9833));
compressor_4_2 u2_3390(.a(t_6725), .b(t_6722), .c(t_6719), .d(t_6716), .cin(t_9830), .o(t_9834), .co(t_9835), .cout(t_9836));
compressor_4_2 u2_3391(.a(t_6736), .b(t_6733), .c(t_6730), .d(t_6727), .cin(t_9833), .o(t_9837), .co(t_9838), .cout(t_9839));
compressor_4_2 u2_3392(.a(t_6737), .b(t_6734), .c(t_6731), .d(t_6728), .cin(t_9836), .o(t_9840), .co(t_9841), .cout(t_9842));
compressor_4_2 u2_3393(.a(t_6748), .b(t_6745), .c(t_6742), .d(t_6739), .cin(t_9839), .o(t_9843), .co(t_9844), .cout(t_9845));
compressor_4_2 u2_3394(.a(t_6746), .b(t_6743), .c(t_6740), .d(t_824), .cin(t_9842), .o(t_9846), .co(t_9847), .cout(t_9848));
compressor_4_2 u2_3395(.a(t_6757), .b(t_6754), .c(t_6751), .d(t_6749), .cin(t_9845), .o(t_9849), .co(t_9850), .cout(t_9851));
compressor_4_2 u2_3396(.a(t_6761), .b(t_6758), .c(t_6755), .d(t_6752), .cin(t_9848), .o(t_9852), .co(t_9853), .cout(t_9854));
compressor_4_2 u2_3397(.a(t_6772), .b(t_6769), .c(t_6766), .d(t_6763), .cin(t_9851), .o(t_9855), .co(t_9856), .cout(t_9857));
compressor_4_2 u2_3398(.a(t_6770), .b(t_6767), .c(t_6764), .d(t_874), .cin(t_9854), .o(t_9858), .co(t_9859), .cout(t_9860));
compressor_4_2 u2_3399(.a(t_6780), .b(t_6777), .c(t_6776), .d(t_6773), .cin(t_9857), .o(t_9861), .co(t_9862), .cout(t_9863));
half_adder u0_3400(.a(t_6786), .b(t_6783), .o(t_9864), .cout(t_9865));
compressor_4_2 u2_3401(.a(t_6787), .b(t_6784), .c(t_6781), .d(t_6778), .cin(t_9860), .o(t_9866), .co(t_9867), .cout(t_9868));
compressor_4_2 u2_3402(.a(t_6798), .b(t_6795), .c(t_6792), .d(t_6789), .cin(t_9863), .o(t_9869), .co(t_9870), .cout(t_9871));
compressor_4_2 u2_3403(.a(t_6799), .b(t_6796), .c(t_6793), .d(t_6790), .cin(t_9868), .o(t_9872), .co(t_9873), .cout(t_9874));
compressor_4_2 u2_3404(.a(t_6809), .b(t_6806), .c(t_6803), .d(t_6802), .cin(t_9871), .o(t_9875), .co(t_9876), .cout(t_9877));
half_adder u0_3405(.a(t_6815), .b(t_6812), .o(t_9878), .cout(t_9879));
compressor_4_2 u2_3406(.a(t_6813), .b(t_6810), .c(t_6807), .d(t_6804), .cin(t_9874), .o(t_9880), .co(t_9881), .cout(t_9882));
compressor_4_2 u2_3407(.a(t_6823), .b(t_6820), .c(t_6817), .d(t_6816), .cin(t_9877), .o(t_9883), .co(t_9884), .cout(t_9885));
half_adder u0_3408(.a(t_6829), .b(t_6826), .o(t_9886), .cout(t_9887));
compressor_4_2 u2_3409(.a(t_6827), .b(t_6824), .c(t_6821), .d(t_6818), .cin(t_9882), .o(t_9888), .co(t_9889), .cout(t_9890));
compressor_4_2 u2_3410(.a(t_6837), .b(t_6834), .c(t_6831), .d(t_6830), .cin(t_9885), .o(t_9891), .co(t_9892), .cout(t_9893));
half_adder u0_3411(.a(t_6843), .b(t_6840), .o(t_9894), .cout(t_9895));
compressor_4_2 u2_3412(.a(t_6841), .b(t_6838), .c(t_6835), .d(t_6832), .cin(t_9890), .o(t_9896), .co(t_9897), .cout(t_9898));
compressor_4_2 u2_3413(.a(t_6851), .b(t_6848), .c(t_6845), .d(t_6844), .cin(t_9893), .o(t_9899), .co(t_9900), .cout(t_9901));
half_adder u0_3414(.a(t_6857), .b(t_6854), .o(t_9902), .cout(t_9903));
compressor_4_2 u2_3415(.a(t_6855), .b(t_6852), .c(t_6849), .d(t_6846), .cin(t_9898), .o(t_9904), .co(t_9905), .cout(t_9906));
compressor_4_2 u2_3416(.a(t_6865), .b(t_6862), .c(t_6859), .d(t_6858), .cin(t_9901), .o(t_9907), .co(t_9908), .cout(t_9909));
half_adder u0_3417(.a(t_6871), .b(t_6868), .o(t_9910), .cout(t_9911));
compressor_4_2 u2_3418(.a(t_6866), .b(t_6863), .c(t_6860), .d(t_1061), .cin(t_9906), .o(t_9912), .co(t_9913), .cout(t_9914));
compressor_4_2 u2_3419(.a(t_6876), .b(t_6873), .c(t_6872), .d(t_6869), .cin(t_9909), .o(t_9915), .co(t_9916), .cout(t_9917));
compressor_3_2 u1_3420(.a(t_6885), .b(t_6882), .cin(t_6879), .o(t_9918), .cout(t_9919));
compressor_4_2 u2_3421(.a(t_6883), .b(t_6880), .c(t_6877), .d(t_6874), .cin(t_9914), .o(t_9920), .co(t_9921), .cout(t_9922));
compressor_4_2 u2_3422(.a(t_6893), .b(t_6890), .c(t_6887), .d(t_6886), .cin(t_9917), .o(t_9923), .co(t_9924), .cout(t_9925));
half_adder u0_3423(.a(t_6899), .b(t_6896), .o(t_9926), .cout(t_9927));
compressor_4_2 u2_3424(.a(t_6894), .b(t_6891), .c(t_6888), .d(t_1120), .cin(t_9922), .o(t_9928), .co(t_9929), .cout(t_9930));
compressor_4_2 u2_3425(.a(t_6904), .b(t_6901), .c(t_6900), .d(t_6897), .cin(t_9925), .o(t_9931), .co(t_9932), .cout(t_9933));
compressor_3_2 u1_3426(.a(t_6913), .b(t_6910), .cin(t_6907), .o(t_9934), .cout(t_9935));
compressor_4_2 u2_3427(.a(t_6911), .b(t_6908), .c(t_6905), .d(t_6902), .cin(t_9930), .o(t_9936), .co(t_9937), .cout(t_9938));
compressor_4_2 u2_3428(.a(t_6921), .b(t_6918), .c(t_6915), .d(t_6914), .cin(t_9933), .o(t_9939), .co(t_9940), .cout(t_9941));
half_adder u0_3429(.a(t_6927), .b(t_6924), .o(t_9942), .cout(t_9943));
compressor_4_2 u2_3430(.a(t_6925), .b(t_6922), .c(t_6919), .d(t_6916), .cin(t_9938), .o(t_9944), .co(t_9945), .cout(t_9946));
compressor_4_2 u2_3431(.a(t_6936), .b(t_6933), .c(t_6930), .d(t_6928), .cin(t_9941), .o(t_9947), .co(t_9948), .cout(t_9949));
half_adder u0_3432(.a(t_6942), .b(t_6939), .o(t_9950), .cout(t_9951));
compressor_4_2 u2_3433(.a(t_6940), .b(t_6937), .c(t_6934), .d(t_6931), .cin(t_9946), .o(t_9952), .co(t_9953), .cout(t_9954));
compressor_4_2 u2_3434(.a(t_6951), .b(t_6948), .c(t_6945), .d(t_6943), .cin(t_9949), .o(t_9955), .co(t_9956), .cout(t_9957));
half_adder u0_3435(.a(t_6957), .b(t_6954), .o(t_9958), .cout(t_9959));
compressor_4_2 u2_3436(.a(t_6955), .b(t_6952), .c(t_6949), .d(t_6946), .cin(t_9954), .o(t_9960), .co(t_9961), .cout(t_9962));
compressor_4_2 u2_3437(.a(t_6966), .b(t_6963), .c(t_6960), .d(t_6958), .cin(t_9957), .o(t_9963), .co(t_9964), .cout(t_9965));
half_adder u0_3438(.a(t_6972), .b(t_6969), .o(t_9966), .cout(t_9967));
compressor_4_2 u2_3439(.a(t_6967), .b(t_6964), .c(t_6961), .d(t_1270), .cin(t_9962), .o(t_9968), .co(t_9969), .cout(t_9970));
compressor_4_2 u2_3440(.a(t_6978), .b(t_6975), .c(t_6973), .d(t_6970), .cin(t_9965), .o(t_9971), .co(t_9972), .cout(t_9973));
compressor_3_2 u1_3441(.a(t_6987), .b(t_6984), .cin(t_6981), .o(t_9974), .cout(t_9975));
compressor_4_2 u2_3442(.a(t_6985), .b(t_6982), .c(t_6979), .d(t_6976), .cin(t_9970), .o(t_9976), .co(t_9977), .cout(t_9978));
compressor_4_2 u2_3443(.a(t_6996), .b(t_6993), .c(t_6990), .d(t_6988), .cin(t_9973), .o(t_9979), .co(t_9980), .cout(t_9981));
compressor_3_2 u1_3444(.a(t_7005), .b(t_7002), .cin(t_6999), .o(t_9982), .cout(t_9983));
compressor_4_2 u2_3445(.a(t_6997), .b(t_6994), .c(t_6991), .d(t_1332), .cin(t_9978), .o(t_9984), .co(t_9985), .cout(t_9986));
compressor_4_2 u2_3446(.a(t_7007), .b(t_7006), .c(t_7003), .d(t_7000), .cin(t_9981), .o(t_9987), .co(t_9988), .cout(t_9989));
compressor_3_2 u1_3447(.a(t_7016), .b(t_7013), .cin(t_7010), .o(t_9990), .cout(t_9991));
compressor_4_2 u2_3448(.a(t_7017), .b(t_7014), .c(t_7011), .d(t_7008), .cin(t_9986), .o(t_9992), .co(t_9993), .cout(t_9994));
compressor_4_2 u2_3449(.a(t_7028), .b(t_7025), .c(t_7022), .d(t_7020), .cin(t_9989), .o(t_9995), .co(t_9996), .cout(t_9997));
compressor_3_2 u1_3450(.a(t_7037), .b(t_7034), .cin(t_7031), .o(t_9998), .cout(t_9999));
compressor_4_2 u2_3451(.a(t_7032), .b(t_7029), .c(t_7026), .d(t_7023), .cin(t_9994), .o(t_10000), .co(t_10001), .cout(t_10002));
compressor_4_2 u2_3452(.a(t_7042), .b(t_7039), .c(t_7038), .d(t_7035), .cin(t_9997), .o(t_10003), .co(t_10004), .cout(t_10005));
compressor_3_2 u1_3453(.a(t_7051), .b(t_7048), .cin(t_7045), .o(t_10006), .cout(t_10007));
compressor_4_2 u2_3454(.a(t_7049), .b(t_7046), .c(t_7043), .d(t_7040), .cin(t_10002), .o(t_10008), .co(t_10009), .cout(t_10010));
compressor_4_2 u2_3455(.a(t_7059), .b(t_7056), .c(t_7055), .d(t_7052), .cin(t_10005), .o(t_10011), .co(t_10012), .cout(t_10013));
compressor_3_2 u1_3456(.a(t_7068), .b(t_7065), .cin(t_7062), .o(t_10014), .cout(t_10015));
compressor_4_2 u2_3457(.a(t_7066), .b(t_7063), .c(t_7060), .d(t_7057), .cin(t_10010), .o(t_10016), .co(t_10017), .cout(t_10018));
compressor_4_2 u2_3458(.a(t_7076), .b(t_7073), .c(t_7072), .d(t_7069), .cin(t_10013), .o(t_10019), .co(t_10020), .cout(t_10021));
compressor_3_2 u1_3459(.a(t_7085), .b(t_7082), .cin(t_7079), .o(t_10022), .cout(t_10023));
compressor_4_2 u2_3460(.a(t_7083), .b(t_7080), .c(t_7077), .d(t_7074), .cin(t_10018), .o(t_10024), .co(t_10025), .cout(t_10026));
compressor_4_2 u2_3461(.a(t_7093), .b(t_7090), .c(t_7089), .d(t_7086), .cin(t_10021), .o(t_10027), .co(t_10028), .cout(t_10029));
compressor_3_2 u1_3462(.a(t_7102), .b(t_7099), .cin(t_7096), .o(t_10030), .cout(t_10031));
compressor_4_2 u2_3463(.a(t_7100), .b(t_7097), .c(t_7094), .d(t_7091), .cin(t_10026), .o(t_10032), .co(t_10033), .cout(t_10034));
compressor_4_2 u2_3464(.a(t_7110), .b(t_7107), .c(t_7106), .d(t_7103), .cin(t_10029), .o(t_10035), .co(t_10036), .cout(t_10037));
compressor_3_2 u1_3465(.a(t_7119), .b(t_7116), .cin(t_7113), .o(t_10038), .cout(t_10039));
compressor_4_2 u2_3466(.a(t_7114), .b(t_7111), .c(t_7108), .d(t_1561), .cin(t_10034), .o(t_10040), .co(t_10041), .cout(t_10042));
compressor_4_2 u2_3467(.a(t_7124), .b(t_7123), .c(t_7120), .d(t_7117), .cin(t_10037), .o(t_10043), .co(t_10044), .cout(t_10045));
compressor_4_2 u2_3468(.a(t_7139), .b(t_7136), .c(t_7133), .d(t_7130), .cin(t_7127), .o(t_10046), .co(t_10047), .cout(t_10048));
compressor_4_2 u2_3469(.a(t_7134), .b(t_7131), .c(t_7128), .d(t_7125), .cin(t_10042), .o(t_10049), .co(t_10050), .cout(t_10051));
compressor_4_2 u2_3470(.a(t_7144), .b(t_7141), .c(t_7140), .d(t_7137), .cin(t_10045), .o(t_10052), .co(t_10053), .cout(t_10054));
compressor_4_2 u2_3471(.a(t_7156), .b(t_7153), .c(t_7150), .d(t_7147), .cin(t_10048), .o(t_10055), .co(t_10056), .cout(t_10057));
compressor_4_2 u2_3472(.a(t_7148), .b(t_7145), .c(t_7142), .d(t_1632), .cin(t_10051), .o(t_10058), .co(t_10059), .cout(t_10060));
compressor_4_2 u2_3473(.a(t_7158), .b(t_7157), .c(t_7154), .d(t_7151), .cin(t_10054), .o(t_10061), .co(t_10062), .cout(t_10063));
compressor_4_2 u2_3474(.a(t_7170), .b(t_7167), .c(t_7164), .d(t_7161), .cin(t_10057), .o(t_10064), .co(t_10065), .cout(t_10066));
compressor_4_2 u2_3475(.a(t_7168), .b(t_7165), .c(t_7162), .d(t_7159), .cin(t_10060), .o(t_10067), .co(t_10068), .cout(t_10069));
compressor_4_2 u2_3476(.a(t_7178), .b(t_7175), .c(t_7174), .d(t_7171), .cin(t_10063), .o(t_10070), .co(t_10071), .cout(t_10072));
compressor_4_2 u2_3477(.a(t_7190), .b(t_7187), .c(t_7184), .d(t_7181), .cin(t_10066), .o(t_10073), .co(t_10074), .cout(t_10075));
compressor_4_2 u2_3478(.a(t_7185), .b(t_7182), .c(t_7179), .d(t_7176), .cin(t_10069), .o(t_10076), .co(t_10077), .cout(t_10078));
compressor_4_2 u2_3479(.a(t_7196), .b(t_7193), .c(t_7191), .d(t_7188), .cin(t_10072), .o(t_10079), .co(t_10080), .cout(t_10081));
compressor_4_2 u2_3480(.a(t_7208), .b(t_7205), .c(t_7202), .d(t_7199), .cin(t_10075), .o(t_10082), .co(t_10083), .cout(t_10084));
compressor_4_2 u2_3481(.a(t_7203), .b(t_7200), .c(t_7197), .d(t_7194), .cin(t_10078), .o(t_10085), .co(t_10086), .cout(t_10087));
compressor_4_2 u2_3482(.a(t_7214), .b(t_7211), .c(t_7209), .d(t_7206), .cin(t_10081), .o(t_10088), .co(t_10089), .cout(t_10090));
compressor_4_2 u2_3483(.a(t_7226), .b(t_7223), .c(t_7220), .d(t_7217), .cin(t_10084), .o(t_10091), .co(t_10092), .cout(t_10093));
compressor_4_2 u2_3484(.a(t_7221), .b(t_7218), .c(t_7215), .d(t_7212), .cin(t_10087), .o(t_10094), .co(t_10095), .cout(t_10096));
compressor_4_2 u2_3485(.a(t_7232), .b(t_7229), .c(t_7227), .d(t_7224), .cin(t_10090), .o(t_10097), .co(t_10098), .cout(t_10099));
compressor_4_2 u2_3486(.a(t_7244), .b(t_7241), .c(t_7238), .d(t_7235), .cin(t_10093), .o(t_10100), .co(t_10101), .cout(t_10102));
compressor_4_2 u2_3487(.a(t_7236), .b(t_7233), .c(t_7230), .d(t_1812), .cin(t_10096), .o(t_10103), .co(t_10104), .cout(t_10105));
compressor_4_2 u2_3488(.a(t_7247), .b(t_7245), .c(t_7242), .d(t_7239), .cin(t_10099), .o(t_10106), .co(t_10107), .cout(t_10108));
compressor_4_2 u2_3489(.a(t_7259), .b(t_7256), .c(t_7253), .d(t_7250), .cin(t_10102), .o(t_10109), .co(t_10110), .cout(t_10111));
compressor_4_2 u2_3490(.a(t_7257), .b(t_7254), .c(t_7251), .d(t_7248), .cin(t_10105), .o(t_10112), .co(t_10113), .cout(t_10114));
compressor_4_2 u2_3491(.a(t_7268), .b(t_7265), .c(t_7263), .d(t_7260), .cin(t_10108), .o(t_10115), .co(t_10116), .cout(t_10117));
compressor_4_2 u2_3492(.a(t_7280), .b(t_7277), .c(t_7274), .d(t_7271), .cin(t_10111), .o(t_10118), .co(t_10119), .cout(t_10120));
compressor_4_2 u2_3493(.a(t_7272), .b(t_7269), .c(t_7266), .d(t_1886), .cin(t_10114), .o(t_10121), .co(t_10122), .cout(t_10123));
compressor_4_2 u2_3494(.a(t_7284), .b(t_7281), .c(t_7278), .d(t_7275), .cin(t_10117), .o(t_10124), .co(t_10125), .cout(t_10126));
compressor_4_2 u2_3495(.a(t_7294), .b(t_7291), .c(t_7288), .d(t_7285), .cin(t_10120), .o(t_10127), .co(t_10128), .cout(t_10129));
half_adder u0_3496(.a(t_7300), .b(t_7297), .o(t_10130), .cout(t_10131));
compressor_4_2 u2_3497(.a(t_7295), .b(t_7292), .c(t_7289), .d(t_7286), .cin(t_10123), .o(t_10132), .co(t_10133), .cout(t_10134));
compressor_4_2 u2_3498(.a(t_7306), .b(t_7303), .c(t_7301), .d(t_7298), .cin(t_10126), .o(t_10135), .co(t_10136), .cout(t_10137));
compressor_4_2 u2_3499(.a(t_7318), .b(t_7315), .c(t_7312), .d(t_7309), .cin(t_10129), .o(t_10138), .co(t_10139), .cout(t_10140));
compressor_4_2 u2_3500(.a(t_7313), .b(t_7310), .c(t_7307), .d(t_7304), .cin(t_10134), .o(t_10141), .co(t_10142), .cout(t_10143));
compressor_4_2 u2_3501(.a(t_7323), .b(t_7322), .c(t_7319), .d(t_7316), .cin(t_10137), .o(t_10144), .co(t_10145), .cout(t_10146));
compressor_4_2 u2_3502(.a(t_7335), .b(t_7332), .c(t_7329), .d(t_7326), .cin(t_10140), .o(t_10147), .co(t_10148), .cout(t_10149));
half_adder u0_3503(.a(t_7341), .b(t_7338), .o(t_10150), .cout(t_10151));
compressor_4_2 u2_3504(.a(t_7333), .b(t_7330), .c(t_7327), .d(t_7324), .cin(t_10143), .o(t_10152), .co(t_10153), .cout(t_10154));
compressor_4_2 u2_3505(.a(t_7343), .b(t_7342), .c(t_7339), .d(t_7336), .cin(t_10146), .o(t_10155), .co(t_10156), .cout(t_10157));
compressor_4_2 u2_3506(.a(t_7355), .b(t_7352), .c(t_7349), .d(t_7346), .cin(t_10149), .o(t_10158), .co(t_10159), .cout(t_10160));
half_adder u0_3507(.a(t_7361), .b(t_7358), .o(t_10161), .cout(t_10162));
compressor_4_2 u2_3508(.a(t_7353), .b(t_7350), .c(t_7347), .d(t_7344), .cin(t_10154), .o(t_10163), .co(t_10164), .cout(t_10165));
compressor_4_2 u2_3509(.a(t_7363), .b(t_7362), .c(t_7359), .d(t_7356), .cin(t_10157), .o(t_10166), .co(t_10167), .cout(t_10168));
compressor_4_2 u2_3510(.a(t_7375), .b(t_7372), .c(t_7369), .d(t_7366), .cin(t_10160), .o(t_10169), .co(t_10170), .cout(t_10171));
half_adder u0_3511(.a(t_7381), .b(t_7378), .o(t_10172), .cout(t_10173));
compressor_4_2 u2_3512(.a(t_7373), .b(t_7370), .c(t_7367), .d(t_7364), .cin(t_10165), .o(t_10174), .co(t_10175), .cout(t_10176));
compressor_4_2 u2_3513(.a(t_7383), .b(t_7382), .c(t_7379), .d(t_7376), .cin(t_10168), .o(t_10177), .co(t_10178), .cout(t_10179));
compressor_4_2 u2_3514(.a(t_7395), .b(t_7392), .c(t_7389), .d(t_7386), .cin(t_10171), .o(t_10180), .co(t_10181), .cout(t_10182));
half_adder u0_3515(.a(t_7401), .b(t_7398), .o(t_10183), .cout(t_10184));
compressor_4_2 u2_3516(.a(t_7393), .b(t_7390), .c(t_7387), .d(t_7384), .cin(t_10176), .o(t_10185), .co(t_10186), .cout(t_10187));
compressor_4_2 u2_3517(.a(t_7403), .b(t_7402), .c(t_7399), .d(t_7396), .cin(t_10179), .o(t_10188), .co(t_10189), .cout(t_10190));
compressor_4_2 u2_3518(.a(t_7415), .b(t_7412), .c(t_7409), .d(t_7406), .cin(t_10182), .o(t_10191), .co(t_10192), .cout(t_10193));
half_adder u0_3519(.a(t_7421), .b(t_7418), .o(t_10194), .cout(t_10195));
compressor_4_2 u2_3520(.a(t_7410), .b(t_7407), .c(t_7404), .d(t_2157), .cin(t_10187), .o(t_10196), .co(t_10197), .cout(t_10198));
compressor_4_2 u2_3521(.a(t_7422), .b(t_7419), .c(t_7416), .d(t_7413), .cin(t_10190), .o(t_10199), .co(t_10200), .cout(t_10201));
compressor_4_2 u2_3522(.a(t_7432), .b(t_7429), .c(t_7426), .d(t_7423), .cin(t_10193), .o(t_10202), .co(t_10203), .cout(t_10204));
compressor_3_2 u1_3523(.a(t_7441), .b(t_7438), .cin(t_7435), .o(t_10205), .cout(t_10206));
compressor_4_2 u2_3524(.a(t_7433), .b(t_7430), .c(t_7427), .d(t_7424), .cin(t_10198), .o(t_10207), .co(t_10208), .cout(t_10209));
compressor_4_2 u2_3525(.a(t_7443), .b(t_7442), .c(t_7439), .d(t_7436), .cin(t_10201), .o(t_10210), .co(t_10211), .cout(t_10212));
compressor_4_2 u2_3526(.a(t_7455), .b(t_7452), .c(t_7449), .d(t_7446), .cin(t_10204), .o(t_10213), .co(t_10214), .cout(t_10215));
half_adder u0_3527(.a(t_7461), .b(t_7458), .o(t_10216), .cout(t_10217));
compressor_4_2 u2_3528(.a(t_7450), .b(t_7447), .c(t_7444), .d(t_2240), .cin(t_10209), .o(t_10218), .co(t_10219), .cout(t_10220));
compressor_4_2 u2_3529(.a(t_7462), .b(t_7459), .c(t_7456), .d(t_7453), .cin(t_10212), .o(t_10221), .co(t_10222), .cout(t_10223));
compressor_4_2 u2_3530(.a(t_7472), .b(t_7469), .c(t_7466), .d(t_7463), .cin(t_10215), .o(t_10224), .co(t_10225), .cout(t_10226));
compressor_3_2 u1_3531(.a(t_7481), .b(t_7478), .cin(t_7475), .o(t_10227), .cout(t_10228));
compressor_4_2 u2_3532(.a(t_7473), .b(t_7470), .c(t_7467), .d(t_7464), .cin(t_10220), .o(t_10229), .co(t_10230), .cout(t_10231));
compressor_4_2 u2_3533(.a(t_7483), .b(t_7482), .c(t_7479), .d(t_7476), .cin(t_10223), .o(t_10232), .co(t_10233), .cout(t_10234));
compressor_4_2 u2_3534(.a(t_7495), .b(t_7492), .c(t_7489), .d(t_7486), .cin(t_10226), .o(t_10235), .co(t_10236), .cout(t_10237));
half_adder u0_3535(.a(t_7501), .b(t_7498), .o(t_10238), .cout(t_10239));
compressor_4_2 u2_3536(.a(t_7493), .b(t_7490), .c(t_7487), .d(t_7484), .cin(t_10231), .o(t_10240), .co(t_10241), .cout(t_10242));
compressor_4_2 u2_3537(.a(t_7504), .b(t_7502), .c(t_7499), .d(t_7496), .cin(t_10234), .o(t_10243), .co(t_10244), .cout(t_10245));
compressor_4_2 u2_3538(.a(t_7516), .b(t_7513), .c(t_7510), .d(t_7507), .cin(t_10237), .o(t_10246), .co(t_10247), .cout(t_10248));
half_adder u0_3539(.a(t_7522), .b(t_7519), .o(t_10249), .cout(t_10250));
compressor_4_2 u2_3540(.a(t_7514), .b(t_7511), .c(t_7508), .d(t_7505), .cin(t_10242), .o(t_10251), .co(t_10252), .cout(t_10253));
compressor_4_2 u2_3541(.a(t_7525), .b(t_7523), .c(t_7520), .d(t_7517), .cin(t_10245), .o(t_10254), .co(t_10255), .cout(t_10256));
compressor_4_2 u2_3542(.a(t_7537), .b(t_7534), .c(t_7531), .d(t_7528), .cin(t_10248), .o(t_10257), .co(t_10258), .cout(t_10259));
half_adder u0_3543(.a(t_7543), .b(t_7540), .o(t_10260), .cout(t_10261));
compressor_4_2 u2_3544(.a(t_7535), .b(t_7532), .c(t_7529), .d(t_7526), .cin(t_10253), .o(t_10262), .co(t_10263), .cout(t_10264));
compressor_4_2 u2_3545(.a(t_7546), .b(t_7544), .c(t_7541), .d(t_7538), .cin(t_10256), .o(t_10265), .co(t_10266), .cout(t_10267));
compressor_4_2 u2_3546(.a(t_7558), .b(t_7555), .c(t_7552), .d(t_7549), .cin(t_10259), .o(t_10268), .co(t_10269), .cout(t_10270));
half_adder u0_3547(.a(t_7564), .b(t_7561), .o(t_10271), .cout(t_10272));
compressor_4_2 u2_3548(.a(t_7553), .b(t_7550), .c(t_7547), .d(t_2450), .cin(t_10264), .o(t_10273), .co(t_10274), .cout(t_10275));
compressor_4_2 u2_3549(.a(t_7565), .b(t_7562), .c(t_7559), .d(t_7556), .cin(t_10267), .o(t_10276), .co(t_10277), .cout(t_10278));
compressor_4_2 u2_3550(.a(t_7576), .b(t_7573), .c(t_7570), .d(t_7567), .cin(t_10270), .o(t_10279), .co(t_10280), .cout(t_10281));
compressor_3_2 u1_3551(.a(t_7585), .b(t_7582), .cin(t_7579), .o(t_10282), .cout(t_10283));
compressor_4_2 u2_3552(.a(t_7577), .b(t_7574), .c(t_7571), .d(t_7568), .cin(t_10275), .o(t_10284), .co(t_10285), .cout(t_10286));
compressor_4_2 u2_3553(.a(t_7588), .b(t_7586), .c(t_7583), .d(t_7580), .cin(t_10278), .o(t_10287), .co(t_10288), .cout(t_10289));
compressor_4_2 u2_3554(.a(t_7600), .b(t_7597), .c(t_7594), .d(t_7591), .cin(t_10281), .o(t_10290), .co(t_10291), .cout(t_10292));
compressor_3_2 u1_3555(.a(t_7609), .b(t_7606), .cin(t_7603), .o(t_10293), .cout(t_10294));
compressor_4_2 u2_3556(.a(t_7595), .b(t_7592), .c(t_7589), .d(t_2536), .cin(t_10286), .o(t_10295), .co(t_10296), .cout(t_10297));
compressor_4_2 u2_3557(.a(t_7607), .b(t_7604), .c(t_7601), .d(t_7598), .cin(t_10289), .o(t_10298), .co(t_10299), .cout(t_10300));
compressor_4_2 u2_3558(.a(t_7617), .b(t_7614), .c(t_7611), .d(t_7610), .cin(t_10292), .o(t_10301), .co(t_10302), .cout(t_10303));
compressor_3_2 u1_3559(.a(t_7626), .b(t_7623), .cin(t_7620), .o(t_10304), .cout(t_10305));
compressor_4_2 u2_3560(.a(t_7621), .b(t_7618), .c(t_7615), .d(t_7612), .cin(t_10297), .o(t_10306), .co(t_10307), .cout(t_10308));
compressor_4_2 u2_3561(.a(t_7632), .b(t_7630), .c(t_7627), .d(t_7624), .cin(t_10300), .o(t_10309), .co(t_10310), .cout(t_10311));
compressor_4_2 u2_3562(.a(t_7644), .b(t_7641), .c(t_7638), .d(t_7635), .cin(t_10303), .o(t_10312), .co(t_10313), .cout(t_10314));
compressor_3_2 u1_3563(.a(t_7653), .b(t_7650), .cin(t_7647), .o(t_10315), .cout(t_10316));
compressor_4_2 u2_3564(.a(t_7642), .b(t_7639), .c(t_7636), .d(t_7633), .cin(t_10308), .o(t_10317), .co(t_10318), .cout(t_10319));
compressor_4_2 u2_3565(.a(t_7654), .b(t_7651), .c(t_7648), .d(t_7645), .cin(t_10311), .o(t_10320), .co(t_10321), .cout(t_10322));
compressor_4_2 u2_3566(.a(t_7664), .b(t_7661), .c(t_7658), .d(t_7655), .cin(t_10314), .o(t_10323), .co(t_10324), .cout(t_10325));
compressor_3_2 u1_3567(.a(t_7673), .b(t_7670), .cin(t_7667), .o(t_10326), .cout(t_10327));
compressor_4_2 u2_3568(.a(t_7665), .b(t_7662), .c(t_7659), .d(t_7656), .cin(t_10319), .o(t_10328), .co(t_10329), .cout(t_10330));
compressor_4_2 u2_3569(.a(t_7677), .b(t_7674), .c(t_7671), .d(t_7668), .cin(t_10322), .o(t_10331), .co(t_10332), .cout(t_10333));
compressor_4_2 u2_3570(.a(t_7687), .b(t_7684), .c(t_7681), .d(t_7678), .cin(t_10325), .o(t_10334), .co(t_10335), .cout(t_10336));
compressor_3_2 u1_3571(.a(t_7696), .b(t_7693), .cin(t_7690), .o(t_10337), .cout(t_10338));
compressor_4_2 u2_3572(.a(t_7688), .b(t_7685), .c(t_7682), .d(t_7679), .cin(t_10330), .o(t_10339), .co(t_10340), .cout(t_10341));
compressor_4_2 u2_3573(.a(t_7700), .b(t_7697), .c(t_7694), .d(t_7691), .cin(t_10333), .o(t_10342), .co(t_10343), .cout(t_10344));
compressor_4_2 u2_3574(.a(t_7710), .b(t_7707), .c(t_7704), .d(t_7701), .cin(t_10336), .o(t_10345), .co(t_10346), .cout(t_10347));
compressor_3_2 u1_3575(.a(t_7719), .b(t_7716), .cin(t_7713), .o(t_10348), .cout(t_10349));
compressor_4_2 u2_3576(.a(t_7711), .b(t_7708), .c(t_7705), .d(t_7702), .cin(t_10341), .o(t_10350), .co(t_10351), .cout(t_10352));
compressor_4_2 u2_3577(.a(t_7723), .b(t_7720), .c(t_7717), .d(t_7714), .cin(t_10344), .o(t_10353), .co(t_10354), .cout(t_10355));
compressor_4_2 u2_3578(.a(t_7733), .b(t_7730), .c(t_7727), .d(t_7724), .cin(t_10347), .o(t_10356), .co(t_10357), .cout(t_10358));
compressor_3_2 u1_3579(.a(t_7742), .b(t_7739), .cin(t_7736), .o(t_10359), .cout(t_10360));
compressor_4_2 u2_3580(.a(t_7734), .b(t_7731), .c(t_7728), .d(t_7725), .cin(t_10352), .o(t_10361), .co(t_10362), .cout(t_10363));
compressor_4_2 u2_3581(.a(t_7746), .b(t_7743), .c(t_7740), .d(t_7737), .cin(t_10355), .o(t_10364), .co(t_10365), .cout(t_10366));
compressor_4_2 u2_3582(.a(t_7756), .b(t_7753), .c(t_7750), .d(t_7747), .cin(t_10358), .o(t_10367), .co(t_10368), .cout(t_10369));
compressor_3_2 u1_3583(.a(t_7765), .b(t_7762), .cin(t_7759), .o(t_10370), .cout(t_10371));
compressor_4_2 u2_3584(.a(t_7754), .b(t_7751), .c(t_7748), .d(t_2849), .cin(t_10363), .o(t_10372), .co(t_10373), .cout(t_10374));
compressor_4_2 u2_3585(.a(t_7766), .b(t_7763), .c(t_7760), .d(t_7757), .cin(t_10366), .o(t_10375), .co(t_10376), .cout(t_10377));
compressor_4_2 u2_3586(.a(t_7776), .b(t_7773), .c(t_7770), .d(t_7769), .cin(t_10369), .o(t_10378), .co(t_10379), .cout(t_10380));
compressor_4_2 u2_3587(.a(t_7791), .b(t_7788), .c(t_7785), .d(t_7782), .cin(t_7779), .o(t_10381), .co(t_10382), .cout(t_10383));
compressor_4_2 u2_3588(.a(t_7780), .b(t_7777), .c(t_7774), .d(t_7771), .cin(t_10374), .o(t_10384), .co(t_10385), .cout(t_10386));
compressor_4_2 u2_3589(.a(t_7792), .b(t_7789), .c(t_7786), .d(t_7783), .cin(t_10377), .o(t_10387), .co(t_10388), .cout(t_10389));
compressor_4_2 u2_3590(.a(t_7802), .b(t_7799), .c(t_7796), .d(t_7793), .cin(t_10380), .o(t_10390), .co(t_10391), .cout(t_10392));
compressor_4_2 u2_3591(.a(t_7814), .b(t_7811), .c(t_7808), .d(t_7805), .cin(t_10383), .o(t_10393), .co(t_10394), .cout(t_10395));
compressor_4_2 u2_3592(.a(t_7800), .b(t_7797), .c(t_7794), .d(t_2944), .cin(t_10386), .o(t_10396), .co(t_10397), .cout(t_10398));
compressor_4_2 u2_3593(.a(t_7812), .b(t_7809), .c(t_7806), .d(t_7803), .cin(t_10389), .o(t_10399), .co(t_10400), .cout(t_10401));
compressor_4_2 u2_3594(.a(t_7822), .b(t_7819), .c(t_7816), .d(t_7815), .cin(t_10392), .o(t_10402), .co(t_10403), .cout(t_10404));
compressor_4_2 u2_3595(.a(t_7834), .b(t_7831), .c(t_7828), .d(t_7825), .cin(t_10395), .o(t_10405), .co(t_10406), .cout(t_10407));
compressor_4_2 u2_3596(.a(t_7826), .b(t_7823), .c(t_7820), .d(t_7817), .cin(t_10398), .o(t_10408), .co(t_10409), .cout(t_10410));
compressor_4_2 u2_3597(.a(t_7838), .b(t_7835), .c(t_7832), .d(t_7829), .cin(t_10401), .o(t_10411), .co(t_10412), .cout(t_10413));
compressor_4_2 u2_3598(.a(t_7848), .b(t_7845), .c(t_7842), .d(t_7839), .cin(t_10404), .o(t_10414), .co(t_10415), .cout(t_10416));
compressor_4_2 u2_3599(.a(t_7860), .b(t_7857), .c(t_7854), .d(t_7851), .cin(t_10407), .o(t_10417), .co(t_10418), .cout(t_10419));
compressor_4_2 u2_3600(.a(t_7849), .b(t_7846), .c(t_7843), .d(t_7840), .cin(t_10410), .o(t_10420), .co(t_10421), .cout(t_10422));
compressor_4_2 u2_3601(.a(t_7861), .b(t_7858), .c(t_7855), .d(t_7852), .cin(t_10413), .o(t_10423), .co(t_10424), .cout(t_10425));
compressor_4_2 u2_3602(.a(t_7872), .b(t_7869), .c(t_7866), .d(t_7863), .cin(t_10416), .o(t_10426), .co(t_10427), .cout(t_10428));
compressor_4_2 u2_3603(.a(t_7884), .b(t_7881), .c(t_7878), .d(t_7875), .cin(t_10419), .o(t_10429), .co(t_10430), .cout(t_10431));
compressor_4_2 u2_3604(.a(t_7873), .b(t_7870), .c(t_7867), .d(t_7864), .cin(t_10422), .o(t_10432), .co(t_10433), .cout(t_10434));
compressor_4_2 u2_3605(.a(t_7885), .b(t_7882), .c(t_7879), .d(t_7876), .cin(t_10425), .o(t_10435), .co(t_10436), .cout(t_10437));
compressor_4_2 u2_3606(.a(t_7896), .b(t_7893), .c(t_7890), .d(t_7887), .cin(t_10428), .o(t_10438), .co(t_10439), .cout(t_10440));
compressor_4_2 u2_3607(.a(t_7908), .b(t_7905), .c(t_7902), .d(t_7899), .cin(t_10431), .o(t_10441), .co(t_10442), .cout(t_10443));
compressor_4_2 u2_3608(.a(t_7897), .b(t_7894), .c(t_7891), .d(t_7888), .cin(t_10434), .o(t_10444), .co(t_10445), .cout(t_10446));
compressor_4_2 u2_3609(.a(t_7909), .b(t_7906), .c(t_7903), .d(t_7900), .cin(t_10437), .o(t_10447), .co(t_10448), .cout(t_10449));
compressor_4_2 u2_3610(.a(t_7920), .b(t_7917), .c(t_7914), .d(t_7911), .cin(t_10440), .o(t_10450), .co(t_10451), .cout(t_10452));
compressor_4_2 u2_3611(.a(t_7932), .b(t_7929), .c(t_7926), .d(t_7923), .cin(t_10443), .o(t_10453), .co(t_10454), .cout(t_10455));
compressor_4_2 u2_3612(.a(t_7918), .b(t_7915), .c(t_7912), .d(t_3181), .cin(t_10446), .o(t_10456), .co(t_10457), .cout(t_10458));
compressor_4_2 u2_3613(.a(t_7930), .b(t_7927), .c(t_7924), .d(t_7921), .cin(t_10449), .o(t_10459), .co(t_10460), .cout(t_10461));
compressor_4_2 u2_3614(.a(t_7941), .b(t_7938), .c(t_7935), .d(t_7933), .cin(t_10452), .o(t_10462), .co(t_10463), .cout(t_10464));
compressor_4_2 u2_3615(.a(t_7953), .b(t_7950), .c(t_7947), .d(t_7944), .cin(t_10455), .o(t_10465), .co(t_10466), .cout(t_10467));
compressor_4_2 u2_3616(.a(t_7942), .b(t_7939), .c(t_7936), .d(t_3229), .cin(t_10458), .o(t_10468), .co(t_10469), .cout(t_10470));
compressor_4_2 u2_3617(.a(t_7954), .b(t_7951), .c(t_7948), .d(t_7945), .cin(t_10461), .o(t_10471), .co(t_10472), .cout(t_10473));
compressor_4_2 u2_3618(.a(t_7965), .b(t_7962), .c(t_7959), .d(t_7957), .cin(t_10464), .o(t_10474), .co(t_10475), .cout(t_10476));
compressor_4_2 u2_3619(.a(t_7977), .b(t_7974), .c(t_7971), .d(t_7968), .cin(t_10467), .o(t_10477), .co(t_10478), .cout(t_10479));
compressor_4_2 u2_3620(.a(t_7969), .b(t_7966), .c(t_7963), .d(t_7960), .cin(t_10470), .o(t_10480), .co(t_10481), .cout(t_10482));
compressor_4_2 u2_3621(.a(t_7981), .b(t_7978), .c(t_7975), .d(t_7972), .cin(t_10473), .o(t_10483), .co(t_10484), .cout(t_10485));
compressor_4_2 u2_3622(.a(t_7992), .b(t_7989), .c(t_7986), .d(t_7983), .cin(t_10476), .o(t_10486), .co(t_10487), .cout(t_10488));
compressor_4_2 u2_3623(.a(t_8004), .b(t_8001), .c(t_7998), .d(t_7995), .cin(t_10479), .o(t_10489), .co(t_10490), .cout(t_10491));
compressor_4_2 u2_3624(.a(t_7993), .b(t_7990), .c(t_7987), .d(t_7984), .cin(t_10482), .o(t_10492), .co(t_10493), .cout(t_10494));
compressor_4_2 u2_3625(.a(t_8005), .b(t_8002), .c(t_7999), .d(t_7996), .cin(t_10485), .o(t_10495), .co(t_10496), .cout(t_10497));
compressor_4_2 u2_3626(.a(t_8016), .b(t_8013), .c(t_8010), .d(t_8007), .cin(t_10488), .o(t_10498), .co(t_10499), .cout(t_10500));
compressor_4_2 u2_3627(.a(t_8028), .b(t_8025), .c(t_8022), .d(t_8019), .cin(t_10491), .o(t_10501), .co(t_10502), .cout(t_10503));
compressor_4_2 u2_3628(.a(t_8014), .b(t_8011), .c(t_8008), .d(t_3373), .cin(t_10494), .o(t_10504), .co(t_10505), .cout(t_10506));
compressor_4_2 u2_3629(.a(t_8026), .b(t_8023), .c(t_8020), .d(t_8017), .cin(t_10497), .o(t_10507), .co(t_10508), .cout(t_10509));
compressor_4_2 u2_3630(.a(t_8037), .b(t_8034), .c(t_8031), .d(t_8029), .cin(t_10500), .o(t_10510), .co(t_10511), .cout(t_10512));
compressor_4_2 u2_3631(.a(t_8049), .b(t_8046), .c(t_8043), .d(t_8040), .cin(t_10503), .o(t_10513), .co(t_10514), .cout(t_10515));
compressor_4_2 u2_3632(.a(t_8041), .b(t_8038), .c(t_8035), .d(t_8032), .cin(t_10506), .o(t_10516), .co(t_10517), .cout(t_10518));
compressor_4_2 u2_3633(.a(t_8053), .b(t_8050), .c(t_8047), .d(t_8044), .cin(t_10509), .o(t_10519), .co(t_10520), .cout(t_10521));
compressor_4_2 u2_3634(.a(t_8064), .b(t_8061), .c(t_8058), .d(t_8055), .cin(t_10512), .o(t_10522), .co(t_10523), .cout(t_10524));
compressor_4_2 u2_3635(.a(t_8076), .b(t_8073), .c(t_8070), .d(t_8067), .cin(t_10515), .o(t_10525), .co(t_10526), .cout(t_10527));
compressor_4_2 u2_3636(.a(t_8065), .b(t_8062), .c(t_8059), .d(t_8056), .cin(t_10518), .o(t_10528), .co(t_10529), .cout(t_10530));
compressor_4_2 u2_3637(.a(t_8077), .b(t_8074), .c(t_8071), .d(t_8068), .cin(t_10521), .o(t_10531), .co(t_10532), .cout(t_10533));
compressor_4_2 u2_3638(.a(t_8088), .b(t_8085), .c(t_8082), .d(t_8079), .cin(t_10524), .o(t_10534), .co(t_10535), .cout(t_10536));
compressor_4_2 u2_3639(.a(t_8100), .b(t_8097), .c(t_8094), .d(t_8091), .cin(t_10527), .o(t_10537), .co(t_10538), .cout(t_10539));
compressor_4_2 u2_3640(.a(t_8089), .b(t_8086), .c(t_8083), .d(t_8080), .cin(t_10530), .o(t_10540), .co(t_10541), .cout(t_10542));
compressor_4_2 u2_3641(.a(t_8101), .b(t_8098), .c(t_8095), .d(t_8092), .cin(t_10533), .o(t_10543), .co(t_10544), .cout(t_10545));
compressor_4_2 u2_3642(.a(t_8112), .b(t_8109), .c(t_8106), .d(t_8103), .cin(t_10536), .o(t_10546), .co(t_10547), .cout(t_10548));
compressor_4_2 u2_3643(.a(t_8124), .b(t_8121), .c(t_8118), .d(t_8115), .cin(t_10539), .o(t_10549), .co(t_10550), .cout(t_10551));
compressor_4_2 u2_3644(.a(t_8113), .b(t_8110), .c(t_8107), .d(t_8104), .cin(t_10542), .o(t_10552), .co(t_10553), .cout(t_10554));
compressor_4_2 u2_3645(.a(t_8125), .b(t_8122), .c(t_8119), .d(t_8116), .cin(t_10545), .o(t_10555), .co(t_10556), .cout(t_10557));
compressor_4_2 u2_3646(.a(t_8136), .b(t_8133), .c(t_8130), .d(t_8127), .cin(t_10548), .o(t_10558), .co(t_10559), .cout(t_10560));
compressor_4_2 u2_3647(.a(t_8148), .b(t_8145), .c(t_8142), .d(t_8139), .cin(t_10551), .o(t_10561), .co(t_10562), .cout(t_10563));
compressor_4_2 u2_3648(.a(t_8134), .b(t_8131), .c(t_8128), .d(t_3603), .cin(t_10554), .o(t_10564), .co(t_10565), .cout(t_10566));
compressor_4_2 u2_3649(.a(t_8146), .b(t_8143), .c(t_8140), .d(t_8137), .cin(t_10557), .o(t_10567), .co(t_10568), .cout(t_10569));
compressor_4_2 u2_3650(.a(t_8157), .b(t_8154), .c(t_8151), .d(t_8149), .cin(t_10560), .o(t_10570), .co(t_10571), .cout(t_10572));
compressor_4_2 u2_3651(.a(t_8169), .b(t_8166), .c(t_8163), .d(t_8160), .cin(t_10563), .o(t_10573), .co(t_10574), .cout(t_10575));
compressor_4_2 u2_3652(.a(t_8161), .b(t_8158), .c(t_8155), .d(t_8152), .cin(t_10566), .o(t_10576), .co(t_10577), .cout(t_10578));
compressor_4_2 u2_3653(.a(t_8173), .b(t_8170), .c(t_8167), .d(t_8164), .cin(t_10569), .o(t_10579), .co(t_10580), .cout(t_10581));
compressor_4_2 u2_3654(.a(t_8183), .b(t_8180), .c(t_8177), .d(t_8174), .cin(t_10572), .o(t_10582), .co(t_10583), .cout(t_10584));
compressor_4_2 u2_3655(.a(t_8195), .b(t_8192), .c(t_8189), .d(t_8186), .cin(t_10575), .o(t_10585), .co(t_10586), .cout(t_10587));
compressor_4_2 u2_3656(.a(t_8184), .b(t_8181), .c(t_8178), .d(t_8175), .cin(t_10578), .o(t_10588), .co(t_10589), .cout(t_10590));
compressor_4_2 u2_3657(.a(t_8196), .b(t_8193), .c(t_8190), .d(t_8187), .cin(t_10581), .o(t_10591), .co(t_10592), .cout(t_10593));
compressor_4_2 u2_3658(.a(t_8206), .b(t_8203), .c(t_8200), .d(t_8197), .cin(t_10584), .o(t_10594), .co(t_10595), .cout(t_10596));
compressor_4_2 u2_3659(.a(t_8218), .b(t_8215), .c(t_8212), .d(t_8209), .cin(t_10587), .o(t_10597), .co(t_10598), .cout(t_10599));
compressor_4_2 u2_3660(.a(t_8207), .b(t_8204), .c(t_8201), .d(t_8198), .cin(t_10590), .o(t_10600), .co(t_10601), .cout(t_10602));
compressor_4_2 u2_3661(.a(t_8219), .b(t_8216), .c(t_8213), .d(t_8210), .cin(t_10593), .o(t_10603), .co(t_10604), .cout(t_10605));
compressor_4_2 u2_3662(.a(t_8229), .b(t_8226), .c(t_8223), .d(t_8220), .cin(t_10596), .o(t_10606), .co(t_10607), .cout(t_10608));
compressor_4_2 u2_3663(.a(t_8241), .b(t_8238), .c(t_8235), .d(t_8232), .cin(t_10599), .o(t_10609), .co(t_10610), .cout(t_10611));
compressor_4_2 u2_3664(.a(t_8230), .b(t_8227), .c(t_8224), .d(t_8221), .cin(t_10602), .o(t_10612), .co(t_10613), .cout(t_10614));
compressor_4_2 u2_3665(.a(t_8242), .b(t_8239), .c(t_8236), .d(t_8233), .cin(t_10605), .o(t_10615), .co(t_10616), .cout(t_10617));
compressor_4_2 u2_3666(.a(t_8252), .b(t_8249), .c(t_8246), .d(t_8243), .cin(t_10608), .o(t_10618), .co(t_10619), .cout(t_10620));
compressor_4_2 u2_3667(.a(t_8264), .b(t_8261), .c(t_8258), .d(t_8255), .cin(t_10611), .o(t_10621), .co(t_10622), .cout(t_10623));
compressor_4_2 u2_3668(.a(t_8253), .b(t_8250), .c(t_8247), .d(t_8244), .cin(t_10614), .o(t_10624), .co(t_10625), .cout(t_10626));
compressor_4_2 u2_3669(.a(t_8265), .b(t_8262), .c(t_8259), .d(t_8256), .cin(t_10617), .o(t_10627), .co(t_10628), .cout(t_10629));
compressor_4_2 u2_3670(.a(t_8275), .b(t_8272), .c(t_8269), .d(t_8266), .cin(t_10620), .o(t_10630), .co(t_10631), .cout(t_10632));
compressor_4_2 u2_3671(.a(t_8287), .b(t_8284), .c(t_8281), .d(t_8278), .cin(t_10623), .o(t_10633), .co(t_10634), .cout(t_10635));
compressor_4_2 u2_3672(.a(t_8276), .b(t_8273), .c(t_8270), .d(t_8267), .cin(t_10626), .o(t_10636), .co(t_10637), .cout(t_10638));
compressor_4_2 u2_3673(.a(t_8288), .b(t_8285), .c(t_8282), .d(t_8279), .cin(t_10629), .o(t_10639), .co(t_10640), .cout(t_10641));
compressor_4_2 u2_3674(.a(t_8298), .b(t_8295), .c(t_8292), .d(t_8289), .cin(t_10632), .o(t_10642), .co(t_10643), .cout(t_10644));
compressor_4_2 u2_3675(.a(t_8310), .b(t_8307), .c(t_8304), .d(t_8301), .cin(t_10635), .o(t_10645), .co(t_10646), .cout(t_10647));
compressor_4_2 u2_3676(.a(t_8299), .b(t_8296), .c(t_8293), .d(t_8290), .cin(t_10638), .o(t_10648), .co(t_10649), .cout(t_10650));
compressor_4_2 u2_3677(.a(t_8311), .b(t_8308), .c(t_8305), .d(t_8302), .cin(t_10641), .o(t_10651), .co(t_10652), .cout(t_10653));
compressor_4_2 u2_3678(.a(t_8321), .b(t_8318), .c(t_8315), .d(t_8312), .cin(t_10644), .o(t_10654), .co(t_10655), .cout(t_10656));
compressor_4_2 u2_3679(.a(t_8333), .b(t_8330), .c(t_8327), .d(t_8324), .cin(t_10647), .o(t_10657), .co(t_10658), .cout(t_10659));
compressor_4_2 u2_3680(.a(t_8319), .b(t_8316), .c(t_8313), .d(t_3953), .cin(t_10650), .o(t_10660), .co(t_10661), .cout(t_10662));
compressor_4_2 u2_3681(.a(t_8331), .b(t_8328), .c(t_8325), .d(t_8322), .cin(t_10653), .o(t_10663), .co(t_10664), .cout(t_10665));
compressor_4_2 u2_3682(.a(t_8341), .b(t_8338), .c(t_8335), .d(t_8334), .cin(t_10656), .o(t_10666), .co(t_10667), .cout(t_10668));
compressor_4_2 u2_3683(.a(t_8353), .b(t_8350), .c(t_8347), .d(t_8344), .cin(t_10659), .o(t_10669), .co(t_10670), .cout(t_10671));
compressor_4_2 u2_3684(.a(t_8345), .b(t_8342), .c(t_8339), .d(t_8336), .cin(t_10662), .o(t_10672), .co(t_10673), .cout(t_10674));
compressor_4_2 u2_3685(.a(t_8356), .b(t_8354), .c(t_8351), .d(t_8348), .cin(t_10665), .o(t_10675), .co(t_10676), .cout(t_10677));
compressor_4_2 u2_3686(.a(t_8368), .b(t_8365), .c(t_8362), .d(t_8359), .cin(t_10668), .o(t_10678), .co(t_10679), .cout(t_10680));
compressor_3_2 u1_3687(.a(t_8374), .b(t_8371), .cin(t_10671), .o(t_10681), .cout(t_10682));
compressor_4_2 u2_3688(.a(t_8366), .b(t_8363), .c(t_8360), .d(t_8357), .cin(t_10674), .o(t_10683), .co(t_10684), .cout(t_10685));
compressor_4_2 u2_3689(.a(t_8377), .b(t_8375), .c(t_8372), .d(t_8369), .cin(t_10677), .o(t_10686), .co(t_10687), .cout(t_10688));
compressor_4_2 u2_3690(.a(t_8389), .b(t_8386), .c(t_8383), .d(t_8380), .cin(t_10680), .o(t_10689), .co(t_10690), .cout(t_10691));
half_adder u0_3691(.a(t_8395), .b(t_8392), .o(t_10692), .cout(t_10693));
compressor_4_2 u2_3692(.a(t_8384), .b(t_8381), .c(t_8378), .d(t_4079), .cin(t_10685), .o(t_10694), .co(t_10695), .cout(t_10696));
compressor_4_2 u2_3693(.a(t_8396), .b(t_8393), .c(t_8390), .d(t_8387), .cin(t_10688), .o(t_10697), .co(t_10698), .cout(t_10699));
compressor_4_2 u2_3694(.a(t_8407), .b(t_8404), .c(t_8401), .d(t_8398), .cin(t_10691), .o(t_10700), .co(t_10701), .cout(t_10702));
compressor_3_2 u1_3695(.a(t_8416), .b(t_8413), .cin(t_8410), .o(t_10703), .cout(t_10704));
compressor_4_2 u2_3696(.a(t_8408), .b(t_8405), .c(t_8402), .d(t_8399), .cin(t_10696), .o(t_10705), .co(t_10706), .cout(t_10707));
compressor_4_2 u2_3697(.a(t_8419), .b(t_8417), .c(t_8414), .d(t_8411), .cin(t_10699), .o(t_10708), .co(t_10709), .cout(t_10710));
compressor_4_2 u2_3698(.a(t_8431), .b(t_8428), .c(t_8425), .d(t_8422), .cin(t_10702), .o(t_10711), .co(t_10712), .cout(t_10713));
half_adder u0_3699(.a(t_8437), .b(t_8434), .o(t_10714), .cout(t_10715));
compressor_4_2 u2_3700(.a(t_8429), .b(t_8426), .c(t_8423), .d(t_8420), .cin(t_10707), .o(t_10716), .co(t_10717), .cout(t_10718));
compressor_4_2 u2_3701(.a(t_8440), .b(t_8438), .c(t_8435), .d(t_8432), .cin(t_10710), .o(t_10719), .co(t_10720), .cout(t_10721));
compressor_4_2 u2_3702(.a(t_8452), .b(t_8449), .c(t_8446), .d(t_8443), .cin(t_10713), .o(t_10722), .co(t_10723), .cout(t_10724));
half_adder u0_3703(.a(t_8458), .b(t_8455), .o(t_10725), .cout(t_10726));
compressor_4_2 u2_3704(.a(t_8450), .b(t_8447), .c(t_8444), .d(t_8441), .cin(t_10718), .o(t_10727), .co(t_10728), .cout(t_10729));
compressor_4_2 u2_3705(.a(t_8461), .b(t_8459), .c(t_8456), .d(t_8453), .cin(t_10721), .o(t_10730), .co(t_10731), .cout(t_10732));
compressor_4_2 u2_3706(.a(t_8473), .b(t_8470), .c(t_8467), .d(t_8464), .cin(t_10724), .o(t_10733), .co(t_10734), .cout(t_10735));
half_adder u0_3707(.a(t_8479), .b(t_8476), .o(t_10736), .cout(t_10737));
compressor_4_2 u2_3708(.a(t_8471), .b(t_8468), .c(t_8465), .d(t_8462), .cin(t_10729), .o(t_10738), .co(t_10739), .cout(t_10740));
compressor_4_2 u2_3709(.a(t_8482), .b(t_8480), .c(t_8477), .d(t_8474), .cin(t_10732), .o(t_10741), .co(t_10742), .cout(t_10743));
compressor_4_2 u2_3710(.a(t_8494), .b(t_8491), .c(t_8488), .d(t_8485), .cin(t_10735), .o(t_10744), .co(t_10745), .cout(t_10746));
half_adder u0_3711(.a(t_8500), .b(t_8497), .o(t_10747), .cout(t_10748));
compressor_4_2 u2_3712(.a(t_8489), .b(t_8486), .c(t_8483), .d(t_4279), .cin(t_10740), .o(t_10749), .co(t_10750), .cout(t_10751));
compressor_4_2 u2_3713(.a(t_8501), .b(t_8498), .c(t_8495), .d(t_8492), .cin(t_10743), .o(t_10752), .co(t_10753), .cout(t_10754));
compressor_4_2 u2_3714(.a(t_8512), .b(t_8509), .c(t_8506), .d(t_8503), .cin(t_10746), .o(t_10755), .co(t_10756), .cout(t_10757));
compressor_3_2 u1_3715(.a(t_8521), .b(t_8518), .cin(t_8515), .o(t_10758), .cout(t_10759));
compressor_4_2 u2_3716(.a(t_8513), .b(t_8510), .c(t_8507), .d(t_8504), .cin(t_10751), .o(t_10760), .co(t_10761), .cout(t_10762));
compressor_4_2 u2_3717(.a(t_8523), .b(t_8522), .c(t_8519), .d(t_8516), .cin(t_10754), .o(t_10763), .co(t_10764), .cout(t_10765));
compressor_4_2 u2_3718(.a(t_8535), .b(t_8532), .c(t_8529), .d(t_8526), .cin(t_10757), .o(t_10766), .co(t_10767), .cout(t_10768));
half_adder u0_3719(.a(t_8541), .b(t_8538), .o(t_10769), .cout(t_10770));
compressor_4_2 u2_3720(.a(t_8533), .b(t_8530), .c(t_8527), .d(t_8524), .cin(t_10762), .o(t_10771), .co(t_10772), .cout(t_10773));
compressor_4_2 u2_3721(.a(t_8543), .b(t_8542), .c(t_8539), .d(t_8536), .cin(t_10765), .o(t_10774), .co(t_10775), .cout(t_10776));
compressor_4_2 u2_3722(.a(t_8555), .b(t_8552), .c(t_8549), .d(t_8546), .cin(t_10768), .o(t_10777), .co(t_10778), .cout(t_10779));
half_adder u0_3723(.a(t_8561), .b(t_8558), .o(t_10780), .cout(t_10781));
compressor_4_2 u2_3724(.a(t_8553), .b(t_8550), .c(t_8547), .d(t_8544), .cin(t_10773), .o(t_10782), .co(t_10783), .cout(t_10784));
compressor_4_2 u2_3725(.a(t_8563), .b(t_8562), .c(t_8559), .d(t_8556), .cin(t_10776), .o(t_10785), .co(t_10786), .cout(t_10787));
compressor_4_2 u2_3726(.a(t_8575), .b(t_8572), .c(t_8569), .d(t_8566), .cin(t_10779), .o(t_10788), .co(t_10789), .cout(t_10790));
half_adder u0_3727(.a(t_8581), .b(t_8578), .o(t_10791), .cout(t_10792));
compressor_4_2 u2_3728(.a(t_8573), .b(t_8570), .c(t_8567), .d(t_8564), .cin(t_10784), .o(t_10793), .co(t_10794), .cout(t_10795));
compressor_4_2 u2_3729(.a(t_8583), .b(t_8582), .c(t_8579), .d(t_8576), .cin(t_10787), .o(t_10796), .co(t_10797), .cout(t_10798));
compressor_4_2 u2_3730(.a(t_8595), .b(t_8592), .c(t_8589), .d(t_8586), .cin(t_10790), .o(t_10799), .co(t_10800), .cout(t_10801));
half_adder u0_3731(.a(t_8601), .b(t_8598), .o(t_10802), .cout(t_10803));
compressor_4_2 u2_3732(.a(t_8593), .b(t_8590), .c(t_8587), .d(t_8584), .cin(t_10795), .o(t_10804), .co(t_10805), .cout(t_10806));
compressor_4_2 u2_3733(.a(t_8603), .b(t_8602), .c(t_8599), .d(t_8596), .cin(t_10798), .o(t_10807), .co(t_10808), .cout(t_10809));
compressor_4_2 u2_3734(.a(t_8615), .b(t_8612), .c(t_8609), .d(t_8606), .cin(t_10801), .o(t_10810), .co(t_10811), .cout(t_10812));
half_adder u0_3735(.a(t_8621), .b(t_8618), .o(t_10813), .cout(t_10814));
compressor_4_2 u2_3736(.a(t_8613), .b(t_8610), .c(t_8607), .d(t_8604), .cin(t_10806), .o(t_10815), .co(t_10816), .cout(t_10817));
compressor_4_2 u2_3737(.a(t_8623), .b(t_8622), .c(t_8619), .d(t_8616), .cin(t_10809), .o(t_10818), .co(t_10819), .cout(t_10820));
compressor_4_2 u2_3738(.a(t_8635), .b(t_8632), .c(t_8629), .d(t_8626), .cin(t_10812), .o(t_10821), .co(t_10822), .cout(t_10823));
half_adder u0_3739(.a(t_8641), .b(t_8638), .o(t_10824), .cout(t_10825));
compressor_4_2 u2_3740(.a(t_8633), .b(t_8630), .c(t_8627), .d(t_8624), .cin(t_10817), .o(t_10826), .co(t_10827), .cout(t_10828));
compressor_4_2 u2_3741(.a(t_8643), .b(t_8642), .c(t_8639), .d(t_8636), .cin(t_10820), .o(t_10829), .co(t_10830), .cout(t_10831));
compressor_4_2 u2_3742(.a(t_8655), .b(t_8652), .c(t_8649), .d(t_8646), .cin(t_10823), .o(t_10832), .co(t_10833), .cout(t_10834));
half_adder u0_3743(.a(t_8661), .b(t_8658), .o(t_10835), .cout(t_10836));
compressor_4_2 u2_3744(.a(t_8650), .b(t_8647), .c(t_8644), .d(t_4581), .cin(t_10828), .o(t_10837), .co(t_10838), .cout(t_10839));
compressor_4_2 u2_3745(.a(t_8662), .b(t_8659), .c(t_8656), .d(t_8653), .cin(t_10831), .o(t_10840), .co(t_10841), .cout(t_10842));
compressor_4_2 u2_3746(.a(t_8672), .b(t_8669), .c(t_8666), .d(t_8663), .cin(t_10834), .o(t_10843), .co(t_10844), .cout(t_10845));
half_adder u0_3747(.a(t_8678), .b(t_8675), .o(t_10846), .cout(t_10847));
compressor_4_2 u2_3748(.a(t_8673), .b(t_8670), .c(t_8667), .d(t_8664), .cin(t_10839), .o(t_10848), .co(t_10849), .cout(t_10850));
compressor_4_2 u2_3749(.a(t_8684), .b(t_8681), .c(t_8679), .d(t_8676), .cin(t_10842), .o(t_10851), .co(t_10852), .cout(t_10853));
compressor_4_2 u2_3750(.a(t_8696), .b(t_8693), .c(t_8690), .d(t_8687), .cin(t_10845), .o(t_10854), .co(t_10855), .cout(t_10856));
compressor_4_2 u2_3751(.a(t_8691), .b(t_8688), .c(t_8685), .d(t_8682), .cin(t_10850), .o(t_10857), .co(t_10858), .cout(t_10859));
compressor_4_2 u2_3752(.a(t_8702), .b(t_8699), .c(t_8697), .d(t_8694), .cin(t_10853), .o(t_10860), .co(t_10861), .cout(t_10862));
compressor_4_2 u2_3753(.a(t_8714), .b(t_8711), .c(t_8708), .d(t_8705), .cin(t_10856), .o(t_10863), .co(t_10864), .cout(t_10865));
compressor_4_2 u2_3754(.a(t_8706), .b(t_8703), .c(t_8700), .d(t_4689), .cin(t_10859), .o(t_10866), .co(t_10867), .cout(t_10868));
compressor_4_2 u2_3755(.a(t_8717), .b(t_8715), .c(t_8712), .d(t_8709), .cin(t_10862), .o(t_10869), .co(t_10870), .cout(t_10871));
compressor_4_2 u2_3756(.a(t_8729), .b(t_8726), .c(t_8723), .d(t_8720), .cin(t_10865), .o(t_10872), .co(t_10873), .cout(t_10874));
compressor_4_2 u2_3757(.a(t_8727), .b(t_8724), .c(t_8721), .d(t_8718), .cin(t_10868), .o(t_10875), .co(t_10876), .cout(t_10877));
compressor_4_2 u2_3758(.a(t_8738), .b(t_8735), .c(t_8733), .d(t_8730), .cin(t_10871), .o(t_10878), .co(t_10879), .cout(t_10880));
compressor_4_2 u2_3759(.a(t_8750), .b(t_8747), .c(t_8744), .d(t_8741), .cin(t_10874), .o(t_10881), .co(t_10882), .cout(t_10883));
compressor_4_2 u2_3760(.a(t_8745), .b(t_8742), .c(t_8739), .d(t_8736), .cin(t_10877), .o(t_10884), .co(t_10885), .cout(t_10886));
compressor_4_2 u2_3761(.a(t_8756), .b(t_8753), .c(t_8751), .d(t_8748), .cin(t_10880), .o(t_10887), .co(t_10888), .cout(t_10889));
compressor_4_2 u2_3762(.a(t_8768), .b(t_8765), .c(t_8762), .d(t_8759), .cin(t_10883), .o(t_10890), .co(t_10891), .cout(t_10892));
compressor_4_2 u2_3763(.a(t_8763), .b(t_8760), .c(t_8757), .d(t_8754), .cin(t_10886), .o(t_10893), .co(t_10894), .cout(t_10895));
compressor_4_2 u2_3764(.a(t_8774), .b(t_8771), .c(t_8769), .d(t_8766), .cin(t_10889), .o(t_10896), .co(t_10897), .cout(t_10898));
compressor_4_2 u2_3765(.a(t_8786), .b(t_8783), .c(t_8780), .d(t_8777), .cin(t_10892), .o(t_10899), .co(t_10900), .cout(t_10901));
compressor_4_2 u2_3766(.a(t_8781), .b(t_8778), .c(t_8775), .d(t_8772), .cin(t_10895), .o(t_10902), .co(t_10903), .cout(t_10904));
compressor_4_2 u2_3767(.a(t_8792), .b(t_8789), .c(t_8787), .d(t_8784), .cin(t_10898), .o(t_10905), .co(t_10906), .cout(t_10907));
compressor_4_2 u2_3768(.a(t_8804), .b(t_8801), .c(t_8798), .d(t_8795), .cin(t_10901), .o(t_10908), .co(t_10909), .cout(t_10910));
compressor_4_2 u2_3769(.a(t_8796), .b(t_8793), .c(t_8790), .d(t_4859), .cin(t_10904), .o(t_10911), .co(t_10912), .cout(t_10913));
compressor_4_2 u2_3770(.a(t_8807), .b(t_8805), .c(t_8802), .d(t_8799), .cin(t_10907), .o(t_10914), .co(t_10915), .cout(t_10916));
compressor_4_2 u2_3771(.a(t_8819), .b(t_8816), .c(t_8813), .d(t_8810), .cin(t_10910), .o(t_10917), .co(t_10918), .cout(t_10919));
compressor_4_2 u2_3772(.a(t_8817), .b(t_8814), .c(t_8811), .d(t_8808), .cin(t_10913), .o(t_10920), .co(t_10921), .cout(t_10922));
compressor_4_2 u2_3773(.a(t_8827), .b(t_8824), .c(t_8823), .d(t_8820), .cin(t_10916), .o(t_10923), .co(t_10924), .cout(t_10925));
compressor_4_2 u2_3774(.a(t_8839), .b(t_8836), .c(t_8833), .d(t_8830), .cin(t_10919), .o(t_10926), .co(t_10927), .cout(t_10928));
compressor_4_2 u2_3775(.a(t_8834), .b(t_8831), .c(t_8828), .d(t_8825), .cin(t_10922), .o(t_10929), .co(t_10930), .cout(t_10931));
compressor_4_2 u2_3776(.a(t_8844), .b(t_8841), .c(t_8840), .d(t_8837), .cin(t_10925), .o(t_10932), .co(t_10933), .cout(t_10934));
compressor_4_2 u2_3777(.a(t_8856), .b(t_8853), .c(t_8850), .d(t_8847), .cin(t_10928), .o(t_10935), .co(t_10936), .cout(t_10937));
compressor_4_2 u2_3778(.a(t_8851), .b(t_8848), .c(t_8845), .d(t_8842), .cin(t_10931), .o(t_10938), .co(t_10939), .cout(t_10940));
compressor_4_2 u2_3779(.a(t_8861), .b(t_8858), .c(t_8857), .d(t_8854), .cin(t_10934), .o(t_10941), .co(t_10942), .cout(t_10943));
compressor_4_2 u2_3780(.a(t_8873), .b(t_8870), .c(t_8867), .d(t_8864), .cin(t_10937), .o(t_10944), .co(t_10945), .cout(t_10946));
compressor_4_2 u2_3781(.a(t_8868), .b(t_8865), .c(t_8862), .d(t_8859), .cin(t_10940), .o(t_10947), .co(t_10948), .cout(t_10949));
compressor_4_2 u2_3782(.a(t_8878), .b(t_8875), .c(t_8874), .d(t_8871), .cin(t_10943), .o(t_10950), .co(t_10951), .cout(t_10952));
compressor_4_2 u2_3783(.a(t_8890), .b(t_8887), .c(t_8884), .d(t_8881), .cin(t_10946), .o(t_10953), .co(t_10954), .cout(t_10955));
compressor_4_2 u2_3784(.a(t_8885), .b(t_8882), .c(t_8879), .d(t_8876), .cin(t_10949), .o(t_10956), .co(t_10957), .cout(t_10958));
compressor_4_2 u2_3785(.a(t_8895), .b(t_8892), .c(t_8891), .d(t_8888), .cin(t_10952), .o(t_10959), .co(t_10960), .cout(t_10961));
compressor_4_2 u2_3786(.a(t_8907), .b(t_8904), .c(t_8901), .d(t_8898), .cin(t_10955), .o(t_10962), .co(t_10963), .cout(t_10964));
compressor_4_2 u2_3787(.a(t_8902), .b(t_8899), .c(t_8896), .d(t_8893), .cin(t_10958), .o(t_10965), .co(t_10966), .cout(t_10967));
compressor_4_2 u2_3788(.a(t_8912), .b(t_8909), .c(t_8908), .d(t_8905), .cin(t_10961), .o(t_10968), .co(t_10969), .cout(t_10970));
compressor_4_2 u2_3789(.a(t_8924), .b(t_8921), .c(t_8918), .d(t_8915), .cin(t_10964), .o(t_10971), .co(t_10972), .cout(t_10973));
compressor_4_2 u2_3790(.a(t_8919), .b(t_8916), .c(t_8913), .d(t_8910), .cin(t_10967), .o(t_10974), .co(t_10975), .cout(t_10976));
compressor_4_2 u2_3791(.a(t_8929), .b(t_8926), .c(t_8925), .d(t_8922), .cin(t_10970), .o(t_10977), .co(t_10978), .cout(t_10979));
compressor_4_2 u2_3792(.a(t_8941), .b(t_8938), .c(t_8935), .d(t_8932), .cin(t_10973), .o(t_10980), .co(t_10981), .cout(t_10982));
compressor_4_2 u2_3793(.a(t_8933), .b(t_8930), .c(t_8927), .d(t_5113), .cin(t_10976), .o(t_10983), .co(t_10984), .cout(t_10985));
compressor_4_2 u2_3794(.a(t_8943), .b(t_8942), .c(t_8939), .d(t_8936), .cin(t_10979), .o(t_10986), .co(t_10987), .cout(t_10988));
compressor_4_2 u2_3795(.a(t_8955), .b(t_8952), .c(t_8949), .d(t_8946), .cin(t_10982), .o(t_10989), .co(t_10990), .cout(t_10991));
compressor_4_2 u2_3796(.a(t_8953), .b(t_8950), .c(t_8947), .d(t_8944), .cin(t_10985), .o(t_10992), .co(t_10993), .cout(t_10994));
compressor_4_2 u2_3797(.a(t_8964), .b(t_8961), .c(t_8958), .d(t_8956), .cin(t_10988), .o(t_10995), .co(t_10996), .cout(t_10997));
compressor_3_2 u1_3798(.a(t_8970), .b(t_8967), .cin(t_10991), .o(t_10998), .cout(t_10999));
compressor_4_2 u2_3799(.a(t_8968), .b(t_8965), .c(t_8962), .d(t_8959), .cin(t_10994), .o(t_11000), .co(t_11001), .cout(t_11002));
compressor_4_2 u2_3800(.a(t_8979), .b(t_8976), .c(t_8973), .d(t_8971), .cin(t_10997), .o(t_11003), .co(t_11004), .cout(t_11005));
half_adder u0_3801(.a(t_8985), .b(t_8982), .o(t_11006), .cout(t_11007));
compressor_4_2 u2_3802(.a(t_8980), .b(t_8977), .c(t_8974), .d(t_5203), .cin(t_11002), .o(t_11008), .co(t_11009), .cout(t_11010));
compressor_4_2 u2_3803(.a(t_8991), .b(t_8988), .c(t_8986), .d(t_8983), .cin(t_11005), .o(t_11011), .co(t_11012), .cout(t_11013));
compressor_3_2 u1_3804(.a(t_9000), .b(t_8997), .cin(t_8994), .o(t_11014), .cout(t_11015));
compressor_4_2 u2_3805(.a(t_8998), .b(t_8995), .c(t_8992), .d(t_8989), .cin(t_11010), .o(t_11016), .co(t_11017), .cout(t_11018));
compressor_4_2 u2_3806(.a(t_9009), .b(t_9006), .c(t_9003), .d(t_9001), .cin(t_11013), .o(t_11019), .co(t_11020), .cout(t_11021));
half_adder u0_3807(.a(t_9015), .b(t_9012), .o(t_11022), .cout(t_11023));
compressor_4_2 u2_3808(.a(t_9013), .b(t_9010), .c(t_9007), .d(t_9004), .cin(t_11018), .o(t_11024), .co(t_11025), .cout(t_11026));
compressor_4_2 u2_3809(.a(t_9024), .b(t_9021), .c(t_9018), .d(t_9016), .cin(t_11021), .o(t_11027), .co(t_11028), .cout(t_11029));
half_adder u0_3810(.a(t_9030), .b(t_9027), .o(t_11030), .cout(t_11031));
compressor_4_2 u2_3811(.a(t_9028), .b(t_9025), .c(t_9022), .d(t_9019), .cin(t_11026), .o(t_11032), .co(t_11033), .cout(t_11034));
compressor_4_2 u2_3812(.a(t_9039), .b(t_9036), .c(t_9033), .d(t_9031), .cin(t_11029), .o(t_11035), .co(t_11036), .cout(t_11037));
half_adder u0_3813(.a(t_9045), .b(t_9042), .o(t_11038), .cout(t_11039));
compressor_4_2 u2_3814(.a(t_9043), .b(t_9040), .c(t_9037), .d(t_9034), .cin(t_11034), .o(t_11040), .co(t_11041), .cout(t_11042));
compressor_4_2 u2_3815(.a(t_9054), .b(t_9051), .c(t_9048), .d(t_9046), .cin(t_11037), .o(t_11043), .co(t_11044), .cout(t_11045));
half_adder u0_3816(.a(t_9060), .b(t_9057), .o(t_11046), .cout(t_11047));
compressor_4_2 u2_3817(.a(t_9055), .b(t_9052), .c(t_9049), .d(t_5343), .cin(t_11042), .o(t_11048), .co(t_11049), .cout(t_11050));
compressor_4_2 u2_3818(.a(t_9066), .b(t_9063), .c(t_9061), .d(t_9058), .cin(t_11045), .o(t_11051), .co(t_11052), .cout(t_11053));
compressor_3_2 u1_3819(.a(t_9075), .b(t_9072), .cin(t_9069), .o(t_11054), .cout(t_11055));
compressor_4_2 u2_3820(.a(t_9073), .b(t_9070), .c(t_9067), .d(t_9064), .cin(t_11050), .o(t_11056), .co(t_11057), .cout(t_11058));
compressor_4_2 u2_3821(.a(t_9083), .b(t_9080), .c(t_9077), .d(t_9076), .cin(t_11053), .o(t_11059), .co(t_11060), .cout(t_11061));
half_adder u0_3822(.a(t_9089), .b(t_9086), .o(t_11062), .cout(t_11063));
compressor_4_2 u2_3823(.a(t_9087), .b(t_9084), .c(t_9081), .d(t_9078), .cin(t_11058), .o(t_11064), .co(t_11065), .cout(t_11066));
compressor_4_2 u2_3824(.a(t_9097), .b(t_9094), .c(t_9091), .d(t_9090), .cin(t_11061), .o(t_11067), .co(t_11068), .cout(t_11069));
half_adder u0_3825(.a(t_9103), .b(t_9100), .o(t_11070), .cout(t_11071));
compressor_4_2 u2_3826(.a(t_9101), .b(t_9098), .c(t_9095), .d(t_9092), .cin(t_11066), .o(t_11072), .co(t_11073), .cout(t_11074));
compressor_4_2 u2_3827(.a(t_9111), .b(t_9108), .c(t_9105), .d(t_9104), .cin(t_11069), .o(t_11075), .co(t_11076), .cout(t_11077));
half_adder u0_3828(.a(t_9117), .b(t_9114), .o(t_11078), .cout(t_11079));
compressor_4_2 u2_3829(.a(t_9115), .b(t_9112), .c(t_9109), .d(t_9106), .cin(t_11074), .o(t_11080), .co(t_11081), .cout(t_11082));
compressor_4_2 u2_3830(.a(t_9125), .b(t_9122), .c(t_9119), .d(t_9118), .cin(t_11077), .o(t_11083), .co(t_11084), .cout(t_11085));
half_adder u0_3831(.a(t_9131), .b(t_9128), .o(t_11086), .cout(t_11087));
compressor_4_2 u2_3832(.a(t_9129), .b(t_9126), .c(t_9123), .d(t_9120), .cin(t_11082), .o(t_11088), .co(t_11089), .cout(t_11090));
compressor_4_2 u2_3833(.a(t_9139), .b(t_9136), .c(t_9133), .d(t_9132), .cin(t_11085), .o(t_11091), .co(t_11092), .cout(t_11093));
half_adder u0_3834(.a(t_9145), .b(t_9142), .o(t_11094), .cout(t_11095));
compressor_4_2 u2_3835(.a(t_9143), .b(t_9140), .c(t_9137), .d(t_9134), .cin(t_11090), .o(t_11096), .co(t_11097), .cout(t_11098));
compressor_4_2 u2_3836(.a(t_9153), .b(t_9150), .c(t_9147), .d(t_9146), .cin(t_11093), .o(t_11099), .co(t_11100), .cout(t_11101));
half_adder u0_3837(.a(t_9159), .b(t_9156), .o(t_11102), .cout(t_11103));
compressor_4_2 u2_3838(.a(t_9157), .b(t_9154), .c(t_9151), .d(t_9148), .cin(t_11098), .o(t_11104), .co(t_11105), .cout(t_11106));
compressor_4_2 u2_3839(.a(t_9167), .b(t_9164), .c(t_9161), .d(t_9160), .cin(t_11101), .o(t_11107), .co(t_11108), .cout(t_11109));
half_adder u0_3840(.a(t_9173), .b(t_9170), .o(t_11110), .cout(t_11111));
compressor_4_2 u2_3841(.a(t_9168), .b(t_9165), .c(t_9162), .d(t_5549), .cin(t_11106), .o(t_11112), .co(t_11113), .cout(t_11114));
compressor_4_2 u2_3842(.a(t_9178), .b(t_9175), .c(t_9174), .d(t_9171), .cin(t_11109), .o(t_11115), .co(t_11116), .cout(t_11117));
half_adder u0_3843(.a(t_9184), .b(t_9181), .o(t_11118), .cout(t_11119));
compressor_4_2 u2_3844(.a(t_9185), .b(t_9182), .c(t_9179), .d(t_9176), .cin(t_11114), .o(t_11120), .co(t_11121), .cout(t_11122));
compressor_4_2 u2_3845(.a(t_9196), .b(t_9193), .c(t_9190), .d(t_9187), .cin(t_11117), .o(t_11123), .co(t_11124), .cout(t_11125));
compressor_4_2 u2_3846(.a(t_9197), .b(t_9194), .c(t_9191), .d(t_9188), .cin(t_11122), .o(t_11126), .co(t_11127), .cout(t_11128));
compressor_4_2 u2_3847(.a(t_9208), .b(t_9205), .c(t_9202), .d(t_9199), .cin(t_11125), .o(t_11129), .co(t_11130), .cout(t_11131));
compressor_4_2 u2_3848(.a(t_9206), .b(t_9203), .c(t_9200), .d(t_5621), .cin(t_11128), .o(t_11132), .co(t_11133), .cout(t_11134));
compressor_4_2 u2_3849(.a(t_9217), .b(t_9214), .c(t_9211), .d(t_9209), .cin(t_11131), .o(t_11135), .co(t_11136), .cout(t_11137));
compressor_4_2 u2_3850(.a(t_9221), .b(t_9218), .c(t_9215), .d(t_9212), .cin(t_11134), .o(t_11138), .co(t_11139), .cout(t_11140));
compressor_4_2 u2_3851(.a(t_9232), .b(t_9229), .c(t_9226), .d(t_9223), .cin(t_11137), .o(t_11141), .co(t_11142), .cout(t_11143));
compressor_4_2 u2_3852(.a(t_9233), .b(t_9230), .c(t_9227), .d(t_9224), .cin(t_11140), .o(t_11144), .co(t_11145), .cout(t_11146));
compressor_4_2 u2_3853(.a(t_9244), .b(t_9241), .c(t_9238), .d(t_9235), .cin(t_11143), .o(t_11147), .co(t_11148), .cout(t_11149));
compressor_4_2 u2_3854(.a(t_9245), .b(t_9242), .c(t_9239), .d(t_9236), .cin(t_11146), .o(t_11150), .co(t_11151), .cout(t_11152));
compressor_4_2 u2_3855(.a(t_9256), .b(t_9253), .c(t_9250), .d(t_9247), .cin(t_11149), .o(t_11153), .co(t_11154), .cout(t_11155));
compressor_4_2 u2_3856(.a(t_9257), .b(t_9254), .c(t_9251), .d(t_9248), .cin(t_11152), .o(t_11156), .co(t_11157), .cout(t_11158));
compressor_4_2 u2_3857(.a(t_9268), .b(t_9265), .c(t_9262), .d(t_9259), .cin(t_11155), .o(t_11159), .co(t_11160), .cout(t_11161));
compressor_4_2 u2_3858(.a(t_9266), .b(t_9263), .c(t_9260), .d(t_5731), .cin(t_11158), .o(t_11162), .co(t_11163), .cout(t_11164));
compressor_4_2 u2_3859(.a(t_9277), .b(t_9274), .c(t_9271), .d(t_9269), .cin(t_11161), .o(t_11165), .co(t_11166), .cout(t_11167));
compressor_4_2 u2_3860(.a(t_9281), .b(t_9278), .c(t_9275), .d(t_9272), .cin(t_11164), .o(t_11168), .co(t_11169), .cout(t_11170));
compressor_4_2 u2_3861(.a(t_9291), .b(t_9288), .c(t_9285), .d(t_9282), .cin(t_11167), .o(t_11171), .co(t_11172), .cout(t_11173));
compressor_4_2 u2_3862(.a(t_9292), .b(t_9289), .c(t_9286), .d(t_9283), .cin(t_11170), .o(t_11174), .co(t_11175), .cout(t_11176));
compressor_4_2 u2_3863(.a(t_9302), .b(t_9299), .c(t_9296), .d(t_9293), .cin(t_11173), .o(t_11177), .co(t_11178), .cout(t_11179));
compressor_4_2 u2_3864(.a(t_9303), .b(t_9300), .c(t_9297), .d(t_9294), .cin(t_11176), .o(t_11180), .co(t_11181), .cout(t_11182));
compressor_4_2 u2_3865(.a(t_9313), .b(t_9310), .c(t_9307), .d(t_9304), .cin(t_11179), .o(t_11183), .co(t_11184), .cout(t_11185));
compressor_4_2 u2_3866(.a(t_9314), .b(t_9311), .c(t_9308), .d(t_9305), .cin(t_11182), .o(t_11186), .co(t_11187), .cout(t_11188));
compressor_4_2 u2_3867(.a(t_9324), .b(t_9321), .c(t_9318), .d(t_9315), .cin(t_11185), .o(t_11189), .co(t_11190), .cout(t_11191));
compressor_4_2 u2_3868(.a(t_9325), .b(t_9322), .c(t_9319), .d(t_9316), .cin(t_11188), .o(t_11192), .co(t_11193), .cout(t_11194));
compressor_4_2 u2_3869(.a(t_9335), .b(t_9332), .c(t_9329), .d(t_9326), .cin(t_11191), .o(t_11195), .co(t_11196), .cout(t_11197));
compressor_4_2 u2_3870(.a(t_9336), .b(t_9333), .c(t_9330), .d(t_9327), .cin(t_11194), .o(t_11198), .co(t_11199), .cout(t_11200));
compressor_4_2 u2_3871(.a(t_9346), .b(t_9343), .c(t_9340), .d(t_9337), .cin(t_11197), .o(t_11201), .co(t_11202), .cout(t_11203));
compressor_4_2 u2_3872(.a(t_9347), .b(t_9344), .c(t_9341), .d(t_9338), .cin(t_11200), .o(t_11204), .co(t_11205), .cout(t_11206));
compressor_4_2 u2_3873(.a(t_9357), .b(t_9354), .c(t_9351), .d(t_9348), .cin(t_11203), .o(t_11207), .co(t_11208), .cout(t_11209));
compressor_4_2 u2_3874(.a(t_9355), .b(t_9352), .c(t_9349), .d(t_5889), .cin(t_11206), .o(t_11210), .co(t_11211), .cout(t_11212));
compressor_4_2 u2_3875(.a(t_9365), .b(t_9362), .c(t_9359), .d(t_9358), .cin(t_11209), .o(t_11213), .co(t_11214), .cout(t_11215));
compressor_4_2 u2_3876(.a(t_9368), .b(t_9366), .c(t_9363), .d(t_9360), .cin(t_11212), .o(t_11216), .co(t_11217), .cout(t_11218));
compressor_3_2 u1_3877(.a(t_9374), .b(t_9371), .cin(t_11215), .o(t_11219), .cout(t_11220));
compressor_4_2 u2_3878(.a(t_9377), .b(t_9375), .c(t_9372), .d(t_9369), .cin(t_11218), .o(t_11221), .co(t_11222), .cout(t_11223));
half_adder u0_3879(.a(t_9383), .b(t_9380), .o(t_11224), .cout(t_11225));
compressor_4_2 u2_3880(.a(t_9384), .b(t_9381), .c(t_9378), .d(t_5943), .cin(t_11223), .o(t_11226), .co(t_11227), .cout(t_11228));
compressor_3_2 u1_3881(.a(t_9392), .b(t_9389), .cin(t_9386), .o(t_11229), .cout(t_11230));
compressor_4_2 u2_3882(.a(t_9395), .b(t_9393), .c(t_9390), .d(t_9387), .cin(t_11228), .o(t_11231), .co(t_11232), .cout(t_11233));
half_adder u0_3883(.a(t_9401), .b(t_9398), .o(t_11234), .cout(t_11235));
compressor_4_2 u2_3884(.a(t_9404), .b(t_9402), .c(t_9399), .d(t_9396), .cin(t_11233), .o(t_11236), .co(t_11237), .cout(t_11238));
half_adder u0_3885(.a(t_9410), .b(t_9407), .o(t_11239), .cout(t_11240));
compressor_4_2 u2_3886(.a(t_9413), .b(t_9411), .c(t_9408), .d(t_9405), .cin(t_11238), .o(t_11241), .co(t_11242), .cout(t_11243));
half_adder u0_3887(.a(t_9419), .b(t_9416), .o(t_11244), .cout(t_11245));
compressor_4_2 u2_3888(.a(t_9422), .b(t_9420), .c(t_9417), .d(t_9414), .cin(t_11243), .o(t_11246), .co(t_11247), .cout(t_11248));
half_adder u0_3889(.a(t_9428), .b(t_9425), .o(t_11249), .cout(t_11250));
compressor_4_2 u2_3890(.a(t_9429), .b(t_9426), .c(t_9423), .d(t_6023), .cin(t_11248), .o(t_11251), .co(t_11252), .cout(t_11253));
compressor_3_2 u1_3891(.a(t_9437), .b(t_9434), .cin(t_9431), .o(t_11254), .cout(t_11255));
compressor_4_2 u2_3892(.a(t_9439), .b(t_9438), .c(t_9435), .d(t_9432), .cin(t_11253), .o(t_11256), .co(t_11257), .cout(t_11258));
half_adder u0_3893(.a(t_9445), .b(t_9442), .o(t_11259), .cout(t_11260));
compressor_4_2 u2_3894(.a(t_9447), .b(t_9446), .c(t_9443), .d(t_9440), .cin(t_11258), .o(t_11261), .co(t_11262), .cout(t_11263));
half_adder u0_3895(.a(t_9453), .b(t_9450), .o(t_11264), .cout(t_11265));
compressor_4_2 u2_3896(.a(t_9455), .b(t_9454), .c(t_9451), .d(t_9448), .cin(t_11263), .o(t_11266), .co(t_11267), .cout(t_11268));
half_adder u0_3897(.a(t_9461), .b(t_9458), .o(t_11269), .cout(t_11270));
compressor_4_2 u2_3898(.a(t_9463), .b(t_9462), .c(t_9459), .d(t_9456), .cin(t_11268), .o(t_11271), .co(t_11272), .cout(t_11273));
half_adder u0_3899(.a(t_9469), .b(t_9466), .o(t_11274), .cout(t_11275));
compressor_4_2 u2_3900(.a(t_9471), .b(t_9470), .c(t_9467), .d(t_9464), .cin(t_11273), .o(t_11276), .co(t_11277), .cout(t_11278));
half_adder u0_3901(.a(t_9477), .b(t_9474), .o(t_11279), .cout(t_11280));
compressor_4_2 u2_3902(.a(t_9479), .b(t_9478), .c(t_9475), .d(t_9472), .cin(t_11278), .o(t_11281), .co(t_11282), .cout(t_11283));
half_adder u0_3903(.a(t_9485), .b(t_9482), .o(t_11284), .cout(t_11285));
compressor_4_2 u2_3904(.a(t_9487), .b(t_9486), .c(t_9483), .d(t_9480), .cin(t_11283), .o(t_11286), .co(t_11287), .cout(t_11288));
half_adder u0_3905(.a(t_9493), .b(t_9490), .o(t_11289), .cout(t_11290));
compressor_4_2 u2_3906(.a(t_9494), .b(t_9491), .c(t_9488), .d(t_6133), .cin(t_11288), .o(t_11291), .co(t_11292), .cout(t_11293));
half_adder u0_3907(.a(t_9498), .b(t_9495), .o(t_11294), .cout(t_11295));
compressor_4_2 u2_3908(.a(t_9504), .b(t_9501), .c(t_9499), .d(t_9496), .cin(t_11293), .o(t_11296), .co(t_11297), .cout(t_11298));
compressor_4_2 u2_3909(.a(t_9510), .b(t_9507), .c(t_9505), .d(t_9502), .cin(t_11298), .o(t_11299), .co(t_11300), .cout(t_11301));
compressor_4_2 u2_3910(.a(t_9513), .b(t_9511), .c(t_9508), .d(t_6169), .cin(t_11301), .o(t_11302), .co(t_11303), .cout(t_11304));
compressor_4_2 u2_3911(.a(t_9522), .b(t_9519), .c(t_9517), .d(t_9514), .cin(t_11304), .o(t_11305), .co(t_11306), .cout(t_11307));
compressor_4_2 u2_3912(.a(t_9528), .b(t_9525), .c(t_9523), .d(t_9520), .cin(t_11307), .o(t_11308), .co(t_11309), .cout(t_11310));
compressor_4_2 u2_3913(.a(t_9534), .b(t_9531), .c(t_9529), .d(t_9526), .cin(t_11310), .o(t_11311), .co(t_11312), .cout(t_11313));
compressor_4_2 u2_3914(.a(t_9540), .b(t_9537), .c(t_9535), .d(t_9532), .cin(t_11313), .o(t_11314), .co(t_11315), .cout(t_11316));
compressor_4_2 u2_3915(.a(t_9543), .b(t_9541), .c(t_9538), .d(t_6219), .cin(t_11316), .o(t_11317), .co(t_11318), .cout(t_11319));
compressor_4_2 u2_3916(.a(t_9551), .b(t_9548), .c(t_9547), .d(t_9544), .cin(t_11319), .o(t_11320), .co(t_11321), .cout(t_11322));
compressor_4_2 u2_3917(.a(t_9556), .b(t_9553), .c(t_9552), .d(t_9549), .cin(t_11322), .o(t_11323), .co(t_11324), .cout(t_11325));
compressor_4_2 u2_3918(.a(t_9561), .b(t_9558), .c(t_9557), .d(t_9554), .cin(t_11325), .o(t_11326), .co(t_11327), .cout(t_11328));
compressor_4_2 u2_3919(.a(t_9566), .b(t_9563), .c(t_9562), .d(t_9559), .cin(t_11328), .o(t_11329), .co(t_11330), .cout(t_11331));
compressor_4_2 u2_3920(.a(t_9571), .b(t_9568), .c(t_9567), .d(t_9564), .cin(t_11331), .o(t_11332), .co(t_11333), .cout(t_11334));
compressor_4_2 u2_3921(.a(t_9576), .b(t_9573), .c(t_9572), .d(t_9569), .cin(t_11334), .o(t_11335), .co(t_11336), .cout(t_11337));
compressor_4_2 u2_3922(.a(t_9581), .b(t_9578), .c(t_9577), .d(t_9574), .cin(t_11337), .o(t_11338), .co(t_11339), .cout(t_11340));
compressor_4_2 u2_3923(.a(t_9583), .b(t_9582), .c(t_9579), .d(t_6281), .cin(t_11340), .o(t_11341), .co(t_11342), .cout(t_11343));
compressor_3_2 u1_3924(.a(t_9586), .b(t_9584), .cin(t_11343), .o(t_11344), .cout(t_11345));
half_adder u0_3925(.a(t_9589), .b(t_9587), .o(t_11346), .cout(t_11347));
compressor_3_2 u1_3926(.a(t_9592), .b(t_9590), .cin(t_6299), .o(t_11348), .cout(t_11349));
half_adder u0_3927(.a(t_9595), .b(t_9593), .o(t_11350), .cout(t_11351));
half_adder u0_3928(.a(t_9598), .b(t_9596), .o(t_11352), .cout(t_11353));
half_adder u0_3929(.a(t_9601), .b(t_9599), .o(t_11354), .cout(t_11355));
half_adder u0_3930(.a(t_9604), .b(t_9602), .o(t_11356), .cout(t_11357));
compressor_3_2 u1_3931(.a(t_9607), .b(t_9605), .cin(t_6319), .o(t_11358), .cout(t_11359));
half_adder u0_3932(.a(t_9609), .b(t_9608), .o(t_11360), .cout(t_11361));
half_adder u0_3933(.a(t_9611), .b(t_9610), .o(t_11362), .cout(t_11363));
half_adder u0_3934(.a(t_9613), .b(t_9612), .o(t_11364), .cout(t_11365));
half_adder u0_3935(.a(t_9615), .b(t_9614), .o(t_11366), .cout(t_11367));
half_adder u0_3936(.a(t_9617), .b(t_9616), .o(t_11368), .cout(t_11369));
half_adder u0_3937(.a(t_9619), .b(t_9618), .o(t_11370), .cout());

/* u0_3938 Output nets */
wire t_11371,  t_11372;
/* u0_3939 Output nets */
wire t_11373,  t_11374;
/* u0_3940 Output nets */
wire t_11375,  t_11376;
/* u0_3941 Output nets */
wire t_11377,  t_11378;
/* u0_3942 Output nets */
wire t_11379,  t_11380;
/* u0_3943 Output nets */
wire t_11381,  t_11382;
/* u0_3944 Output nets */
wire t_11383,  t_11384;
/* u0_3945 Output nets */
wire t_11385,  t_11386;
/* u0_3946 Output nets */
wire t_11387,  t_11388;
/* u0_3947 Output nets */
wire t_11389,  t_11390;
/* u0_3948 Output nets */
wire t_11391,  t_11392;
/* u0_3949 Output nets */
wire t_11393,  t_11394;
/* u0_3950 Output nets */
wire t_11395,  t_11396;
/* u0_3951 Output nets */
wire t_11397,  t_11398;
/* u1_3952 Output nets */
wire t_11399,  t_11400;
/* u0_3953 Output nets */
wire t_11401,  t_11402;
/* u1_3954 Output nets */
wire t_11403,  t_11404;
/* u1_3955 Output nets */
wire t_11405,  t_11406;
/* u1_3956 Output nets */
wire t_11407,  t_11408;
/* u1_3957 Output nets */
wire t_11409,  t_11410;
/* u1_3958 Output nets */
wire t_11411,  t_11412;
/* u0_3959 Output nets */
wire t_11413,  t_11414;
/* u0_3960 Output nets */
wire t_11415,  t_11416;
/* u1_3961 Output nets */
wire t_11417,  t_11418;
/* u0_3962 Output nets */
wire t_11419,  t_11420;
/* u0_3963 Output nets */
wire t_11421,  t_11422;
/* u0_3964 Output nets */
wire t_11423,  t_11424;
/* u0_3965 Output nets */
wire t_11425,  t_11426;
/* u1_3966 Output nets */
wire t_11427,  t_11428;
/* u1_3967 Output nets */
wire t_11429,  t_11430;
/* u1_3968 Output nets */
wire t_11431,  t_11432;
/* u1_3969 Output nets */
wire t_11433,  t_11434;
/* u1_3970 Output nets */
wire t_11435,  t_11436;
/* u1_3971 Output nets */
wire t_11437,  t_11438;
/* u1_3972 Output nets */
wire t_11439,  t_11440;
/* u1_3973 Output nets */
wire t_11441,  t_11442;
/* u1_3974 Output nets */
wire t_11443,  t_11444;
/* u1_3975 Output nets */
wire t_11445,  t_11446;
/* u1_3976 Output nets */
wire t_11447,  t_11448;
/* u1_3977 Output nets */
wire t_11449,  t_11450;
/* u1_3978 Output nets */
wire t_11451,  t_11452;
/* u1_3979 Output nets */
wire t_11453,  t_11454;
/* u1_3980 Output nets */
wire t_11455,  t_11456;
/* u1_3981 Output nets */
wire t_11457,  t_11458;
/* u1_3982 Output nets */
wire t_11459,  t_11460;
/* u1_3983 Output nets */
wire t_11461,  t_11462;
/* u2_3984 Output nets */
wire t_11463,  t_11464,  t_11465;
/* u2_3985 Output nets */
wire t_11466,  t_11467,  t_11468;
/* u2_3986 Output nets */
wire t_11469,  t_11470,  t_11471;
/* u2_3987 Output nets */
wire t_11472,  t_11473,  t_11474;
/* u2_3988 Output nets */
wire t_11475,  t_11476,  t_11477;
/* u2_3989 Output nets */
wire t_11478,  t_11479,  t_11480;
/* u2_3990 Output nets */
wire t_11481,  t_11482,  t_11483;
/* u2_3991 Output nets */
wire t_11484,  t_11485,  t_11486;
/* u2_3992 Output nets */
wire t_11487,  t_11488,  t_11489;
/* u2_3993 Output nets */
wire t_11490,  t_11491,  t_11492;
/* u2_3994 Output nets */
wire t_11493,  t_11494,  t_11495;
/* u2_3995 Output nets */
wire t_11496,  t_11497,  t_11498;
/* u2_3996 Output nets */
wire t_11499,  t_11500,  t_11501;
/* u2_3997 Output nets */
wire t_11502,  t_11503,  t_11504;
/* u2_3998 Output nets */
wire t_11505,  t_11506,  t_11507;
/* u2_3999 Output nets */
wire t_11508,  t_11509,  t_11510;
/* u2_4000 Output nets */
wire t_11511,  t_11512,  t_11513;
/* u2_4001 Output nets */
wire t_11514,  t_11515,  t_11516;
/* u0_4002 Output nets */
wire t_11517,  t_11518;
/* u2_4003 Output nets */
wire t_11519,  t_11520,  t_11521;
/* u2_4004 Output nets */
wire t_11522,  t_11523,  t_11524;
/* u0_4005 Output nets */
wire t_11525,  t_11526;
/* u2_4006 Output nets */
wire t_11527,  t_11528,  t_11529;
/* u0_4007 Output nets */
wire t_11530,  t_11531;
/* u2_4008 Output nets */
wire t_11532,  t_11533,  t_11534;
/* u0_4009 Output nets */
wire t_11535,  t_11536;
/* u2_4010 Output nets */
wire t_11537,  t_11538,  t_11539;
/* u0_4011 Output nets */
wire t_11540,  t_11541;
/* u2_4012 Output nets */
wire t_11542,  t_11543,  t_11544;
/* u0_4013 Output nets */
wire t_11545,  t_11546;
/* u2_4014 Output nets */
wire t_11547,  t_11548,  t_11549;
/* u0_4015 Output nets */
wire t_11550,  t_11551;
/* u2_4016 Output nets */
wire t_11552,  t_11553,  t_11554;
/* u0_4017 Output nets */
wire t_11555,  t_11556;
/* u2_4018 Output nets */
wire t_11557,  t_11558,  t_11559;
/* u0_4019 Output nets */
wire t_11560,  t_11561;
/* u2_4020 Output nets */
wire t_11562,  t_11563,  t_11564;
/* u0_4021 Output nets */
wire t_11565,  t_11566;
/* u2_4022 Output nets */
wire t_11567,  t_11568,  t_11569;
/* u0_4023 Output nets */
wire t_11570,  t_11571;
/* u2_4024 Output nets */
wire t_11572,  t_11573,  t_11574;
/* u0_4025 Output nets */
wire t_11575,  t_11576;
/* u2_4026 Output nets */
wire t_11577,  t_11578,  t_11579;
/* u0_4027 Output nets */
wire t_11580,  t_11581;
/* u2_4028 Output nets */
wire t_11582,  t_11583,  t_11584;
/* u0_4029 Output nets */
wire t_11585,  t_11586;
/* u2_4030 Output nets */
wire t_11587,  t_11588,  t_11589;
/* u1_4031 Output nets */
wire t_11590,  t_11591;
/* u2_4032 Output nets */
wire t_11592,  t_11593,  t_11594;
/* u0_4033 Output nets */
wire t_11595,  t_11596;
/* u2_4034 Output nets */
wire t_11597,  t_11598,  t_11599;
/* u1_4035 Output nets */
wire t_11600,  t_11601;
/* u2_4036 Output nets */
wire t_11602,  t_11603,  t_11604;
/* u1_4037 Output nets */
wire t_11605,  t_11606;
/* u2_4038 Output nets */
wire t_11607,  t_11608,  t_11609;
/* u1_4039 Output nets */
wire t_11610,  t_11611;
/* u2_4040 Output nets */
wire t_11612,  t_11613,  t_11614;
/* u1_4041 Output nets */
wire t_11615,  t_11616;
/* u2_4042 Output nets */
wire t_11617,  t_11618,  t_11619;
/* u1_4043 Output nets */
wire t_11620,  t_11621;
/* u2_4044 Output nets */
wire t_11622,  t_11623,  t_11624;
/* u0_4045 Output nets */
wire t_11625,  t_11626;
/* u2_4046 Output nets */
wire t_11627,  t_11628,  t_11629;
/* u0_4047 Output nets */
wire t_11630,  t_11631;
/* u2_4048 Output nets */
wire t_11632,  t_11633,  t_11634;
/* u1_4049 Output nets */
wire t_11635,  t_11636;
/* u2_4050 Output nets */
wire t_11637,  t_11638,  t_11639;
/* u0_4051 Output nets */
wire t_11640,  t_11641;
/* u2_4052 Output nets */
wire t_11642,  t_11643,  t_11644;
/* u0_4053 Output nets */
wire t_11645,  t_11646;
/* u2_4054 Output nets */
wire t_11647,  t_11648,  t_11649;
/* u0_4055 Output nets */
wire t_11650,  t_11651;
/* u2_4056 Output nets */
wire t_11652,  t_11653,  t_11654;
/* u0_4057 Output nets */
wire t_11655,  t_11656;
/* u2_4058 Output nets */
wire t_11657,  t_11658,  t_11659;
/* u1_4059 Output nets */
wire t_11660,  t_11661;
/* u2_4060 Output nets */
wire t_11662,  t_11663,  t_11664;
/* u1_4061 Output nets */
wire t_11665,  t_11666;
/* u2_4062 Output nets */
wire t_11667,  t_11668,  t_11669;
/* u1_4063 Output nets */
wire t_11670,  t_11671;
/* u2_4064 Output nets */
wire t_11672,  t_11673,  t_11674;
/* u1_4065 Output nets */
wire t_11675,  t_11676;
/* u2_4066 Output nets */
wire t_11677,  t_11678,  t_11679;
/* u1_4067 Output nets */
wire t_11680,  t_11681;
/* u2_4068 Output nets */
wire t_11682,  t_11683,  t_11684;
/* u1_4069 Output nets */
wire t_11685,  t_11686;
/* u2_4070 Output nets */
wire t_11687,  t_11688,  t_11689;
/* u1_4071 Output nets */
wire t_11690,  t_11691;
/* u2_4072 Output nets */
wire t_11692,  t_11693,  t_11694;
/* u1_4073 Output nets */
wire t_11695,  t_11696;
/* u2_4074 Output nets */
wire t_11697,  t_11698,  t_11699;
/* u1_4075 Output nets */
wire t_11700,  t_11701;
/* u2_4076 Output nets */
wire t_11702,  t_11703,  t_11704;
/* u1_4077 Output nets */
wire t_11705,  t_11706;
/* u2_4078 Output nets */
wire t_11707,  t_11708,  t_11709;
/* u1_4079 Output nets */
wire t_11710,  t_11711;
/* u2_4080 Output nets */
wire t_11712,  t_11713,  t_11714;
/* u1_4081 Output nets */
wire t_11715,  t_11716;
/* u2_4082 Output nets */
wire t_11717,  t_11718,  t_11719;
/* u1_4083 Output nets */
wire t_11720,  t_11721;
/* u2_4084 Output nets */
wire t_11722,  t_11723,  t_11724;
/* u1_4085 Output nets */
wire t_11725,  t_11726;
/* u2_4086 Output nets */
wire t_11727,  t_11728,  t_11729;
/* u1_4087 Output nets */
wire t_11730,  t_11731;
/* u2_4088 Output nets */
wire t_11732,  t_11733,  t_11734;
/* u1_4089 Output nets */
wire t_11735,  t_11736;
/* u2_4090 Output nets */
wire t_11737,  t_11738,  t_11739;
/* u1_4091 Output nets */
wire t_11740,  t_11741;
/* u2_4092 Output nets */
wire t_11742,  t_11743,  t_11744;
/* u1_4093 Output nets */
wire t_11745,  t_11746;
/* u2_4094 Output nets */
wire t_11747,  t_11748,  t_11749;
/* u2_4095 Output nets */
wire t_11750,  t_11751,  t_11752;
/* u2_4096 Output nets */
wire t_11753,  t_11754,  t_11755;
/* u2_4097 Output nets */
wire t_11756,  t_11757,  t_11758;
/* u2_4098 Output nets */
wire t_11759,  t_11760,  t_11761;
/* u2_4099 Output nets */
wire t_11762,  t_11763,  t_11764;
/* u2_4100 Output nets */
wire t_11765,  t_11766,  t_11767;
/* u2_4101 Output nets */
wire t_11768,  t_11769,  t_11770;
/* u2_4102 Output nets */
wire t_11771,  t_11772,  t_11773;
/* u2_4103 Output nets */
wire t_11774,  t_11775,  t_11776;
/* u2_4104 Output nets */
wire t_11777,  t_11778,  t_11779;
/* u2_4105 Output nets */
wire t_11780,  t_11781,  t_11782;
/* u2_4106 Output nets */
wire t_11783,  t_11784,  t_11785;
/* u2_4107 Output nets */
wire t_11786,  t_11787,  t_11788;
/* u2_4108 Output nets */
wire t_11789,  t_11790,  t_11791;
/* u2_4109 Output nets */
wire t_11792,  t_11793,  t_11794;
/* u2_4110 Output nets */
wire t_11795,  t_11796,  t_11797;
/* u2_4111 Output nets */
wire t_11798,  t_11799,  t_11800;
/* u2_4112 Output nets */
wire t_11801,  t_11802,  t_11803;
/* u2_4113 Output nets */
wire t_11804,  t_11805,  t_11806;
/* u2_4114 Output nets */
wire t_11807,  t_11808,  t_11809;
/* u2_4115 Output nets */
wire t_11810,  t_11811,  t_11812;
/* u2_4116 Output nets */
wire t_11813,  t_11814,  t_11815;
/* u2_4117 Output nets */
wire t_11816,  t_11817,  t_11818;
/* u2_4118 Output nets */
wire t_11819,  t_11820,  t_11821;
/* u2_4119 Output nets */
wire t_11822,  t_11823,  t_11824;
/* u2_4120 Output nets */
wire t_11825,  t_11826,  t_11827;
/* u2_4121 Output nets */
wire t_11828,  t_11829,  t_11830;
/* u2_4122 Output nets */
wire t_11831,  t_11832,  t_11833;
/* u2_4123 Output nets */
wire t_11834,  t_11835,  t_11836;
/* u2_4124 Output nets */
wire t_11837,  t_11838,  t_11839;
/* u2_4125 Output nets */
wire t_11840,  t_11841,  t_11842;
/* u2_4126 Output nets */
wire t_11843,  t_11844,  t_11845;
/* u2_4127 Output nets */
wire t_11846,  t_11847,  t_11848;
/* u2_4128 Output nets */
wire t_11849,  t_11850,  t_11851;
/* u2_4129 Output nets */
wire t_11852,  t_11853,  t_11854;
/* u2_4130 Output nets */
wire t_11855,  t_11856,  t_11857;
/* u2_4131 Output nets */
wire t_11858,  t_11859,  t_11860;
/* u2_4132 Output nets */
wire t_11861,  t_11862,  t_11863;
/* u2_4133 Output nets */
wire t_11864,  t_11865,  t_11866;
/* u2_4134 Output nets */
wire t_11867,  t_11868,  t_11869;
/* u2_4135 Output nets */
wire t_11870,  t_11871,  t_11872;
/* u2_4136 Output nets */
wire t_11873,  t_11874,  t_11875;
/* u2_4137 Output nets */
wire t_11876,  t_11877,  t_11878;
/* u2_4138 Output nets */
wire t_11879,  t_11880,  t_11881;
/* u2_4139 Output nets */
wire t_11882,  t_11883,  t_11884;
/* u2_4140 Output nets */
wire t_11885,  t_11886,  t_11887;
/* u2_4141 Output nets */
wire t_11888,  t_11889,  t_11890;
/* u2_4142 Output nets */
wire t_11891,  t_11892,  t_11893;
/* u2_4143 Output nets */
wire t_11894,  t_11895,  t_11896;
/* u2_4144 Output nets */
wire t_11897,  t_11898,  t_11899;
/* u2_4145 Output nets */
wire t_11900,  t_11901,  t_11902;
/* u2_4146 Output nets */
wire t_11903,  t_11904,  t_11905;
/* u2_4147 Output nets */
wire t_11906,  t_11907,  t_11908;
/* u2_4148 Output nets */
wire t_11909,  t_11910,  t_11911;
/* u2_4149 Output nets */
wire t_11912,  t_11913,  t_11914;
/* u2_4150 Output nets */
wire t_11915,  t_11916,  t_11917;
/* u2_4151 Output nets */
wire t_11918,  t_11919,  t_11920;
/* u2_4152 Output nets */
wire t_11921,  t_11922,  t_11923;
/* u2_4153 Output nets */
wire t_11924,  t_11925,  t_11926;
/* u2_4154 Output nets */
wire t_11927,  t_11928,  t_11929;
/* u2_4155 Output nets */
wire t_11930,  t_11931,  t_11932;
/* u2_4156 Output nets */
wire t_11933,  t_11934,  t_11935;
/* u2_4157 Output nets */
wire t_11936,  t_11937,  t_11938;
/* u2_4158 Output nets */
wire t_11939,  t_11940,  t_11941;
/* u2_4159 Output nets */
wire t_11942,  t_11943,  t_11944;
/* u2_4160 Output nets */
wire t_11945,  t_11946,  t_11947;
/* u2_4161 Output nets */
wire t_11948,  t_11949,  t_11950;
/* u2_4162 Output nets */
wire t_11951,  t_11952,  t_11953;
/* u2_4163 Output nets */
wire t_11954,  t_11955,  t_11956;
/* u2_4164 Output nets */
wire t_11957,  t_11958,  t_11959;
/* u2_4165 Output nets */
wire t_11960,  t_11961,  t_11962;
/* u2_4166 Output nets */
wire t_11963,  t_11964,  t_11965;
/* u2_4167 Output nets */
wire t_11966,  t_11967,  t_11968;
/* u2_4168 Output nets */
wire t_11969,  t_11970,  t_11971;
/* u2_4169 Output nets */
wire t_11972,  t_11973,  t_11974;
/* u2_4170 Output nets */
wire t_11975,  t_11976,  t_11977;
/* u2_4171 Output nets */
wire t_11978,  t_11979,  t_11980;
/* u2_4172 Output nets */
wire t_11981,  t_11982,  t_11983;
/* u2_4173 Output nets */
wire t_11984,  t_11985,  t_11986;
/* u2_4174 Output nets */
wire t_11987,  t_11988,  t_11989;
/* u2_4175 Output nets */
wire t_11990,  t_11991,  t_11992;
/* u2_4176 Output nets */
wire t_11993,  t_11994,  t_11995;
/* u2_4177 Output nets */
wire t_11996,  t_11997,  t_11998;
/* u2_4178 Output nets */
wire t_11999,  t_12000,  t_12001;
/* u2_4179 Output nets */
wire t_12002,  t_12003,  t_12004;
/* u2_4180 Output nets */
wire t_12005,  t_12006,  t_12007;
/* u2_4181 Output nets */
wire t_12008,  t_12009,  t_12010;
/* u2_4182 Output nets */
wire t_12011,  t_12012,  t_12013;
/* u2_4183 Output nets */
wire t_12014,  t_12015,  t_12016;
/* u2_4184 Output nets */
wire t_12017,  t_12018,  t_12019;
/* u2_4185 Output nets */
wire t_12020,  t_12021,  t_12022;
/* u2_4186 Output nets */
wire t_12023,  t_12024,  t_12025;
/* u2_4187 Output nets */
wire t_12026,  t_12027,  t_12028;
/* u2_4188 Output nets */
wire t_12029,  t_12030,  t_12031;
/* u2_4189 Output nets */
wire t_12032,  t_12033,  t_12034;
/* u2_4190 Output nets */
wire t_12035,  t_12036,  t_12037;
/* u1_4191 Output nets */
wire t_12038,  t_12039;
/* u2_4192 Output nets */
wire t_12040,  t_12041,  t_12042;
/* u0_4193 Output nets */
wire t_12043,  t_12044;
/* u2_4194 Output nets */
wire t_12045,  t_12046,  t_12047;
/* u1_4195 Output nets */
wire t_12048,  t_12049;
/* u2_4196 Output nets */
wire t_12050,  t_12051,  t_12052;
/* u0_4197 Output nets */
wire t_12053,  t_12054;
/* u2_4198 Output nets */
wire t_12055,  t_12056,  t_12057;
/* u0_4199 Output nets */
wire t_12058,  t_12059;
/* u2_4200 Output nets */
wire t_12060,  t_12061,  t_12062;
/* u0_4201 Output nets */
wire t_12063,  t_12064;
/* u2_4202 Output nets */
wire t_12065,  t_12066,  t_12067;
/* u0_4203 Output nets */
wire t_12068,  t_12069;
/* u2_4204 Output nets */
wire t_12070,  t_12071,  t_12072;
/* u1_4205 Output nets */
wire t_12073,  t_12074;
/* u2_4206 Output nets */
wire t_12075,  t_12076,  t_12077;
/* u0_4207 Output nets */
wire t_12078,  t_12079;
/* u2_4208 Output nets */
wire t_12080,  t_12081,  t_12082;
/* u0_4209 Output nets */
wire t_12083,  t_12084;
/* u2_4210 Output nets */
wire t_12085,  t_12086,  t_12087;
/* u0_4211 Output nets */
wire t_12088,  t_12089;
/* u2_4212 Output nets */
wire t_12090,  t_12091,  t_12092;
/* u0_4213 Output nets */
wire t_12093,  t_12094;
/* u2_4214 Output nets */
wire t_12095,  t_12096,  t_12097;
/* u0_4215 Output nets */
wire t_12098,  t_12099;
/* u2_4216 Output nets */
wire t_12100,  t_12101,  t_12102;
/* u0_4217 Output nets */
wire t_12103,  t_12104;
/* u2_4218 Output nets */
wire t_12105,  t_12106,  t_12107;
/* u0_4219 Output nets */
wire t_12108,  t_12109;
/* u2_4220 Output nets */
wire t_12110,  t_12111,  t_12112;
/* u0_4221 Output nets */
wire t_12113,  t_12114;
/* u2_4222 Output nets */
wire t_12115,  t_12116,  t_12117;
/* u0_4223 Output nets */
wire t_12118,  t_12119;
/* u2_4224 Output nets */
wire t_12120,  t_12121,  t_12122;
/* u0_4225 Output nets */
wire t_12123,  t_12124;
/* u2_4226 Output nets */
wire t_12125,  t_12126,  t_12127;
/* u0_4227 Output nets */
wire t_12128,  t_12129;
/* u2_4228 Output nets */
wire t_12130,  t_12131,  t_12132;
/* u0_4229 Output nets */
wire t_12133,  t_12134;
/* u2_4230 Output nets */
wire t_12135,  t_12136,  t_12137;
/* u0_4231 Output nets */
wire t_12138,  t_12139;
/* u2_4232 Output nets */
wire t_12140,  t_12141,  t_12142;
/* u0_4233 Output nets */
wire t_12143,  t_12144;
/* u2_4234 Output nets */
wire t_12145,  t_12146,  t_12147;
/* u0_4235 Output nets */
wire t_12148,  t_12149;
/* u2_4236 Output nets */
wire t_12150,  t_12151,  t_12152;
/* u0_4237 Output nets */
wire t_12153,  t_12154;
/* u2_4238 Output nets */
wire t_12155,  t_12156,  t_12157;
/* u0_4239 Output nets */
wire t_12158,  t_12159;
/* u2_4240 Output nets */
wire t_12160,  t_12161,  t_12162;
/* u0_4241 Output nets */
wire t_12163,  t_12164;
/* u2_4242 Output nets */
wire t_12165,  t_12166,  t_12167;
/* u0_4243 Output nets */
wire t_12168,  t_12169;
/* u2_4244 Output nets */
wire t_12170,  t_12171,  t_12172;
/* u0_4245 Output nets */
wire t_12173,  t_12174;
/* u2_4246 Output nets */
wire t_12175,  t_12176,  t_12177;
/* u0_4247 Output nets */
wire t_12178,  t_12179;
/* u2_4248 Output nets */
wire t_12180,  t_12181,  t_12182;
/* u0_4249 Output nets */
wire t_12183,  t_12184;
/* u2_4250 Output nets */
wire t_12185,  t_12186,  t_12187;
/* u0_4251 Output nets */
wire t_12188,  t_12189;
/* u2_4252 Output nets */
wire t_12190,  t_12191,  t_12192;
/* u0_4253 Output nets */
wire t_12193,  t_12194;
/* u2_4254 Output nets */
wire t_12195,  t_12196,  t_12197;
/* u2_4255 Output nets */
wire t_12198,  t_12199,  t_12200;
/* u2_4256 Output nets */
wire t_12201,  t_12202,  t_12203;
/* u2_4257 Output nets */
wire t_12204,  t_12205,  t_12206;
/* u2_4258 Output nets */
wire t_12207,  t_12208,  t_12209;
/* u2_4259 Output nets */
wire t_12210,  t_12211,  t_12212;
/* u2_4260 Output nets */
wire t_12213,  t_12214,  t_12215;
/* u2_4261 Output nets */
wire t_12216,  t_12217,  t_12218;
/* u2_4262 Output nets */
wire t_12219,  t_12220,  t_12221;
/* u2_4263 Output nets */
wire t_12222,  t_12223,  t_12224;
/* u2_4264 Output nets */
wire t_12225,  t_12226,  t_12227;
/* u2_4265 Output nets */
wire t_12228,  t_12229,  t_12230;
/* u2_4266 Output nets */
wire t_12231,  t_12232,  t_12233;
/* u2_4267 Output nets */
wire t_12234,  t_12235,  t_12236;
/* u2_4268 Output nets */
wire t_12237,  t_12238,  t_12239;
/* u2_4269 Output nets */
wire t_12240,  t_12241,  t_12242;
/* u2_4270 Output nets */
wire t_12243,  t_12244,  t_12245;
/* u2_4271 Output nets */
wire t_12246,  t_12247,  t_12248;
/* u2_4272 Output nets */
wire t_12249,  t_12250,  t_12251;
/* u2_4273 Output nets */
wire t_12252,  t_12253,  t_12254;
/* u2_4274 Output nets */
wire t_12255,  t_12256,  t_12257;
/* u2_4275 Output nets */
wire t_12258,  t_12259,  t_12260;
/* u2_4276 Output nets */
wire t_12261,  t_12262,  t_12263;
/* u2_4277 Output nets */
wire t_12264,  t_12265,  t_12266;
/* u2_4278 Output nets */
wire t_12267,  t_12268,  t_12269;
/* u2_4279 Output nets */
wire t_12270,  t_12271,  t_12272;
/* u2_4280 Output nets */
wire t_12273,  t_12274,  t_12275;
/* u2_4281 Output nets */
wire t_12276,  t_12277,  t_12278;
/* u2_4282 Output nets */
wire t_12279,  t_12280,  t_12281;
/* u2_4283 Output nets */
wire t_12282,  t_12283,  t_12284;
/* u2_4284 Output nets */
wire t_12285,  t_12286,  t_12287;
/* u2_4285 Output nets */
wire t_12288,  t_12289,  t_12290;
/* u1_4286 Output nets */
wire t_12291,  t_12292;
/* u0_4287 Output nets */
wire t_12293,  t_12294;
/* u1_4288 Output nets */
wire t_12295,  t_12296;
/* u0_4289 Output nets */
wire t_12297,  t_12298;
/* u0_4290 Output nets */
wire t_12299,  t_12300;
/* u0_4291 Output nets */
wire t_12301,  t_12302;
/* u0_4292 Output nets */
wire t_12303,  t_12304;
/* u1_4293 Output nets */
wire t_12305,  t_12306;
/* u0_4294 Output nets */
wire t_12307,  t_12308;
/* u0_4295 Output nets */
wire t_12309,  t_12310;
/* u0_4296 Output nets */
wire t_12311,  t_12312;
/* u0_4297 Output nets */
wire t_12313,  t_12314;
/* u0_4298 Output nets */
wire t_12315,  t_12316;
/* u0_4299 Output nets */
wire t_12317,  t_12318;
/* u0_4300 Output nets */
wire t_12319,  t_12320;
/* u0_4301 Output nets */
wire t_12321,  t_12322;
/* u0_4302 Output nets */
wire t_12323,  t_12324;
/* u0_4303 Output nets */
wire t_12325,  t_12326;
/* u0_4304 Output nets */
wire t_12327,  t_12328;
/* u0_4305 Output nets */
wire t_12329,  t_12330;
/* u0_4306 Output nets */
wire t_12331,  t_12332;
/* u0_4307 Output nets */
wire t_12333,  t_12334;
/* u0_4308 Output nets */
wire t_12335,  t_12336;
/* u0_4309 Output nets */
wire t_12337,  t_12338;
/* u0_4310 Output nets */
wire t_12339,  t_12340;
/* u0_4311 Output nets */
wire t_12341,  t_12342;
/* u0_4312 Output nets */
wire t_12343,  t_12344;
/* u0_4313 Output nets */
wire t_12345,  t_12346;
/* u0_4314 Output nets */
wire t_12347,  t_12348;
/* u0_4315 Output nets */
wire t_12349;

/* compress stage 4 */
half_adder u0_3938(.a(t_9621), .b(t_6337), .o(t_11371), .cout(t_11372));
half_adder u0_3939(.a(t_9624), .b(t_9623), .o(t_11373), .cout(t_11374));
half_adder u0_3940(.a(t_9626), .b(t_9625), .o(t_11375), .cout(t_11376));
half_adder u0_3941(.a(t_9628), .b(t_9627), .o(t_11377), .cout(t_11378));
half_adder u0_3942(.a(t_9630), .b(t_9629), .o(t_11379), .cout(t_11380));
half_adder u0_3943(.a(t_9632), .b(t_9631), .o(t_11381), .cout(t_11382));
half_adder u0_3944(.a(t_9634), .b(t_9633), .o(t_11383), .cout(t_11384));
half_adder u0_3945(.a(t_9636), .b(t_9635), .o(t_11385), .cout(t_11386));
half_adder u0_3946(.a(t_9638), .b(t_9637), .o(t_11387), .cout(t_11388));
half_adder u0_3947(.a(t_9640), .b(t_9639), .o(t_11389), .cout(t_11390));
half_adder u0_3948(.a(t_9642), .b(t_9641), .o(t_11391), .cout(t_11392));
half_adder u0_3949(.a(t_9644), .b(t_9643), .o(t_11393), .cout(t_11394));
half_adder u0_3950(.a(t_9646), .b(t_9645), .o(t_11395), .cout(t_11396));
half_adder u0_3951(.a(t_9648), .b(t_9647), .o(t_11397), .cout(t_11398));
compressor_3_2 u1_3952(.a(t_9650), .b(t_9649), .cin(t_6375), .o(t_11399), .cout(t_11400));
half_adder u0_3953(.a(t_9652), .b(t_9651), .o(t_11401), .cout(t_11402));
compressor_3_2 u1_3954(.a(t_9654), .b(t_9653), .cin(t_6386), .o(t_11403), .cout(t_11404));
compressor_3_2 u1_3955(.a(t_9656), .b(t_9655), .cin(t_6391), .o(t_11405), .cout(t_11406));
compressor_3_2 u1_3956(.a(t_9658), .b(t_9657), .cin(t_6396), .o(t_11407), .cout(t_11408));
compressor_3_2 u1_3957(.a(t_9660), .b(t_9659), .cin(t_6401), .o(t_11409), .cout(t_11410));
compressor_3_2 u1_3958(.a(t_9662), .b(t_9661), .cin(t_6406), .o(t_11411), .cout(t_11412));
half_adder u0_3959(.a(t_9664), .b(t_9663), .o(t_11413), .cout(t_11414));
half_adder u0_3960(.a(t_9667), .b(t_9665), .o(t_11415), .cout(t_11416));
compressor_3_2 u1_3961(.a(t_9670), .b(t_9668), .cin(t_6421), .o(t_11417), .cout(t_11418));
half_adder u0_3962(.a(t_9673), .b(t_9671), .o(t_11419), .cout(t_11420));
half_adder u0_3963(.a(t_9676), .b(t_9674), .o(t_11421), .cout(t_11422));
half_adder u0_3964(.a(t_9679), .b(t_9677), .o(t_11423), .cout(t_11424));
half_adder u0_3965(.a(t_9682), .b(t_9680), .o(t_11425), .cout(t_11426));
compressor_3_2 u1_3966(.a(t_9685), .b(t_9683), .cin(t_6450), .o(t_11427), .cout(t_11428));
compressor_3_2 u1_3967(.a(t_9688), .b(t_9686), .cin(t_6459), .o(t_11429), .cout(t_11430));
compressor_3_2 u1_3968(.a(t_9694), .b(t_9691), .cin(t_9689), .o(t_11431), .cout(t_11432));
compressor_3_2 u1_3969(.a(t_9695), .b(t_9692), .cin(t_6473), .o(t_11433), .cout(t_11434));
compressor_3_2 u1_3970(.a(t_9702), .b(t_9699), .cin(t_9697), .o(t_11435), .cout(t_11436));
compressor_3_2 u1_3971(.a(t_9704), .b(t_9703), .cin(t_9700), .o(t_11437), .cout(t_11438));
compressor_3_2 u1_3972(.a(t_9709), .b(t_9708), .cin(t_9705), .o(t_11439), .cout(t_11440));
compressor_3_2 u1_3973(.a(t_9714), .b(t_9713), .cin(t_9710), .o(t_11441), .cout(t_11442));
compressor_3_2 u1_3974(.a(t_9719), .b(t_9718), .cin(t_9715), .o(t_11443), .cout(t_11444));
compressor_3_2 u1_3975(.a(t_9724), .b(t_9723), .cin(t_9720), .o(t_11445), .cout(t_11446));
compressor_3_2 u1_3976(.a(t_9729), .b(t_9728), .cin(t_9725), .o(t_11447), .cout(t_11448));
compressor_3_2 u1_3977(.a(t_9734), .b(t_9733), .cin(t_9730), .o(t_11449), .cout(t_11450));
compressor_3_2 u1_3978(.a(t_9739), .b(t_9738), .cin(t_9735), .o(t_11451), .cout(t_11452));
compressor_3_2 u1_3979(.a(t_9744), .b(t_9743), .cin(t_9740), .o(t_11453), .cout(t_11454));
compressor_3_2 u1_3980(.a(t_9749), .b(t_9748), .cin(t_9745), .o(t_11455), .cout(t_11456));
compressor_3_2 u1_3981(.a(t_9754), .b(t_9753), .cin(t_9750), .o(t_11457), .cout(t_11458));
compressor_3_2 u1_3982(.a(t_9759), .b(t_9758), .cin(t_9755), .o(t_11459), .cout(t_11460));
compressor_3_2 u1_3983(.a(t_9764), .b(t_9763), .cin(t_9760), .o(t_11461), .cout(t_11462));
compressor_4_2 u2_3984(.a(t_9772), .b(t_9769), .c(t_9768), .d(t_9765), .cin(t_6601), .o(t_11463), .co(t_11464), .cout(t_11465));
compressor_4_2 u2_3985(.a(t_9777), .b(t_9774), .c(t_9773), .d(t_9770), .cin(t_11465), .o(t_11466), .co(t_11467), .cout(t_11468));
compressor_4_2 u2_3986(.a(t_9779), .b(t_9778), .c(t_9775), .d(t_6624), .cin(t_11468), .o(t_11469), .co(t_11470), .cout(t_11471));
compressor_4_2 u2_3987(.a(t_9784), .b(t_9783), .c(t_9780), .d(t_6635), .cin(t_11471), .o(t_11472), .co(t_11473), .cout(t_11474));
compressor_4_2 u2_3988(.a(t_9789), .b(t_9788), .c(t_9785), .d(t_6646), .cin(t_11474), .o(t_11475), .co(t_11476), .cout(t_11477));
compressor_4_2 u2_3989(.a(t_9794), .b(t_9793), .c(t_9790), .d(t_6657), .cin(t_11477), .o(t_11478), .co(t_11479), .cout(t_11480));
compressor_4_2 u2_3990(.a(t_9799), .b(t_9798), .c(t_9795), .d(t_6668), .cin(t_11480), .o(t_11481), .co(t_11482), .cout(t_11483));
compressor_4_2 u2_3991(.a(t_9807), .b(t_9804), .c(t_9803), .d(t_9800), .cin(t_11483), .o(t_11484), .co(t_11485), .cout(t_11486));
compressor_4_2 u2_3992(.a(t_9813), .b(t_9810), .c(t_9808), .d(t_9805), .cin(t_11486), .o(t_11487), .co(t_11488), .cout(t_11489));
compressor_4_2 u2_3993(.a(t_9816), .b(t_9814), .c(t_9811), .d(t_6701), .cin(t_11489), .o(t_11490), .co(t_11491), .cout(t_11492));
compressor_4_2 u2_3994(.a(t_9825), .b(t_9822), .c(t_9820), .d(t_9817), .cin(t_11492), .o(t_11493), .co(t_11494), .cout(t_11495));
compressor_4_2 u2_3995(.a(t_9831), .b(t_9828), .c(t_9826), .d(t_9823), .cin(t_11495), .o(t_11496), .co(t_11497), .cout(t_11498));
compressor_4_2 u2_3996(.a(t_9837), .b(t_9834), .c(t_9832), .d(t_9829), .cin(t_11498), .o(t_11499), .co(t_11500), .cout(t_11501));
compressor_4_2 u2_3997(.a(t_9843), .b(t_9840), .c(t_9838), .d(t_9835), .cin(t_11501), .o(t_11502), .co(t_11503), .cout(t_11504));
compressor_4_2 u2_3998(.a(t_9846), .b(t_9844), .c(t_9841), .d(t_6760), .cin(t_11504), .o(t_11505), .co(t_11506), .cout(t_11507));
compressor_4_2 u2_3999(.a(t_9852), .b(t_9850), .c(t_9847), .d(t_6775), .cin(t_11507), .o(t_11508), .co(t_11509), .cout(t_11510));
compressor_4_2 u2_4000(.a(t_9861), .b(t_9858), .c(t_9856), .d(t_9853), .cin(t_11510), .o(t_11511), .co(t_11512), .cout(t_11513));
compressor_4_2 u2_4001(.a(t_9865), .b(t_9862), .c(t_9859), .d(t_6801), .cin(t_11513), .o(t_11514), .co(t_11515), .cout(t_11516));
half_adder u0_4002(.a(t_9869), .b(t_9866), .o(t_11517), .cout(t_11518));
compressor_4_2 u2_4003(.a(t_9875), .b(t_9872), .c(t_9870), .d(t_9867), .cin(t_11516), .o(t_11519), .co(t_11520), .cout(t_11521));
compressor_4_2 u2_4004(.a(t_9880), .b(t_9879), .c(t_9876), .d(t_9873), .cin(t_11521), .o(t_11522), .co(t_11523), .cout(t_11524));
half_adder u0_4005(.a(t_9886), .b(t_9883), .o(t_11525), .cout(t_11526));
compressor_4_2 u2_4006(.a(t_9888), .b(t_9887), .c(t_9884), .d(t_9881), .cin(t_11524), .o(t_11527), .co(t_11528), .cout(t_11529));
half_adder u0_4007(.a(t_9894), .b(t_9891), .o(t_11530), .cout(t_11531));
compressor_4_2 u2_4008(.a(t_9896), .b(t_9895), .c(t_9892), .d(t_9889), .cin(t_11529), .o(t_11532), .co(t_11533), .cout(t_11534));
half_adder u0_4009(.a(t_9902), .b(t_9899), .o(t_11535), .cout(t_11536));
compressor_4_2 u2_4010(.a(t_9904), .b(t_9903), .c(t_9900), .d(t_9897), .cin(t_11534), .o(t_11537), .co(t_11538), .cout(t_11539));
half_adder u0_4011(.a(t_9910), .b(t_9907), .o(t_11540), .cout(t_11541));
compressor_4_2 u2_4012(.a(t_9912), .b(t_9911), .c(t_9908), .d(t_9905), .cin(t_11539), .o(t_11542), .co(t_11543), .cout(t_11544));
half_adder u0_4013(.a(t_9918), .b(t_9915), .o(t_11545), .cout(t_11546));
compressor_4_2 u2_4014(.a(t_9920), .b(t_9919), .c(t_9916), .d(t_9913), .cin(t_11544), .o(t_11547), .co(t_11548), .cout(t_11549));
half_adder u0_4015(.a(t_9926), .b(t_9923), .o(t_11550), .cout(t_11551));
compressor_4_2 u2_4016(.a(t_9928), .b(t_9927), .c(t_9924), .d(t_9921), .cin(t_11549), .o(t_11552), .co(t_11553), .cout(t_11554));
half_adder u0_4017(.a(t_9934), .b(t_9931), .o(t_11555), .cout(t_11556));
compressor_4_2 u2_4018(.a(t_9936), .b(t_9935), .c(t_9932), .d(t_9929), .cin(t_11554), .o(t_11557), .co(t_11558), .cout(t_11559));
half_adder u0_4019(.a(t_9942), .b(t_9939), .o(t_11560), .cout(t_11561));
compressor_4_2 u2_4020(.a(t_9944), .b(t_9943), .c(t_9940), .d(t_9937), .cin(t_11559), .o(t_11562), .co(t_11563), .cout(t_11564));
half_adder u0_4021(.a(t_9950), .b(t_9947), .o(t_11565), .cout(t_11566));
compressor_4_2 u2_4022(.a(t_9952), .b(t_9951), .c(t_9948), .d(t_9945), .cin(t_11564), .o(t_11567), .co(t_11568), .cout(t_11569));
half_adder u0_4023(.a(t_9958), .b(t_9955), .o(t_11570), .cout(t_11571));
compressor_4_2 u2_4024(.a(t_9960), .b(t_9959), .c(t_9956), .d(t_9953), .cin(t_11569), .o(t_11572), .co(t_11573), .cout(t_11574));
half_adder u0_4025(.a(t_9966), .b(t_9963), .o(t_11575), .cout(t_11576));
compressor_4_2 u2_4026(.a(t_9968), .b(t_9967), .c(t_9964), .d(t_9961), .cin(t_11574), .o(t_11577), .co(t_11578), .cout(t_11579));
half_adder u0_4027(.a(t_9974), .b(t_9971), .o(t_11580), .cout(t_11581));
compressor_4_2 u2_4028(.a(t_9976), .b(t_9975), .c(t_9972), .d(t_9969), .cin(t_11579), .o(t_11582), .co(t_11583), .cout(t_11584));
half_adder u0_4029(.a(t_9982), .b(t_9979), .o(t_11585), .cout(t_11586));
compressor_4_2 u2_4030(.a(t_9983), .b(t_9980), .c(t_9977), .d(t_7019), .cin(t_11584), .o(t_11587), .co(t_11588), .cout(t_11589));
compressor_3_2 u1_4031(.a(t_9990), .b(t_9987), .cin(t_9984), .o(t_11590), .cout(t_11591));
compressor_4_2 u2_4032(.a(t_9992), .b(t_9991), .c(t_9988), .d(t_9985), .cin(t_11589), .o(t_11592), .co(t_11593), .cout(t_11594));
half_adder u0_4033(.a(t_9998), .b(t_9995), .o(t_11595), .cout(t_11596));
compressor_4_2 u2_4034(.a(t_9999), .b(t_9996), .c(t_9993), .d(t_7054), .cin(t_11594), .o(t_11597), .co(t_11598), .cout(t_11599));
compressor_3_2 u1_4035(.a(t_10006), .b(t_10003), .cin(t_10000), .o(t_11600), .cout(t_11601));
compressor_4_2 u2_4036(.a(t_10007), .b(t_10004), .c(t_10001), .d(t_7071), .cin(t_11599), .o(t_11602), .co(t_11603), .cout(t_11604));
compressor_3_2 u1_4037(.a(t_10014), .b(t_10011), .cin(t_10008), .o(t_11605), .cout(t_11606));
compressor_4_2 u2_4038(.a(t_10015), .b(t_10012), .c(t_10009), .d(t_7088), .cin(t_11604), .o(t_11607), .co(t_11608), .cout(t_11609));
compressor_3_2 u1_4039(.a(t_10022), .b(t_10019), .cin(t_10016), .o(t_11610), .cout(t_11611));
compressor_4_2 u2_4040(.a(t_10023), .b(t_10020), .c(t_10017), .d(t_7105), .cin(t_11609), .o(t_11612), .co(t_11613), .cout(t_11614));
compressor_3_2 u1_4041(.a(t_10030), .b(t_10027), .cin(t_10024), .o(t_11615), .cout(t_11616));
compressor_4_2 u2_4042(.a(t_10031), .b(t_10028), .c(t_10025), .d(t_7122), .cin(t_11614), .o(t_11617), .co(t_11618), .cout(t_11619));
compressor_3_2 u1_4043(.a(t_10038), .b(t_10035), .cin(t_10032), .o(t_11620), .cout(t_11621));
compressor_4_2 u2_4044(.a(t_10040), .b(t_10039), .c(t_10036), .d(t_10033), .cin(t_11619), .o(t_11622), .co(t_11623), .cout(t_11624));
half_adder u0_4045(.a(t_10046), .b(t_10043), .o(t_11625), .cout(t_11626));
compressor_4_2 u2_4046(.a(t_10049), .b(t_10047), .c(t_10044), .d(t_10041), .cin(t_11624), .o(t_11627), .co(t_11628), .cout(t_11629));
half_adder u0_4047(.a(t_10055), .b(t_10052), .o(t_11630), .cout(t_11631));
compressor_4_2 u2_4048(.a(t_10056), .b(t_10053), .c(t_10050), .d(t_7173), .cin(t_11629), .o(t_11632), .co(t_11633), .cout(t_11634));
compressor_3_2 u1_4049(.a(t_10064), .b(t_10061), .cin(t_10058), .o(t_11635), .cout(t_11636));
compressor_4_2 u2_4050(.a(t_10067), .b(t_10065), .c(t_10062), .d(t_10059), .cin(t_11634), .o(t_11637), .co(t_11638), .cout(t_11639));
half_adder u0_4051(.a(t_10073), .b(t_10070), .o(t_11640), .cout(t_11641));
compressor_4_2 u2_4052(.a(t_10076), .b(t_10074), .c(t_10071), .d(t_10068), .cin(t_11639), .o(t_11642), .co(t_11643), .cout(t_11644));
half_adder u0_4053(.a(t_10082), .b(t_10079), .o(t_11645), .cout(t_11646));
compressor_4_2 u2_4054(.a(t_10085), .b(t_10083), .c(t_10080), .d(t_10077), .cin(t_11644), .o(t_11647), .co(t_11648), .cout(t_11649));
half_adder u0_4055(.a(t_10091), .b(t_10088), .o(t_11650), .cout(t_11651));
compressor_4_2 u2_4056(.a(t_10094), .b(t_10092), .c(t_10089), .d(t_10086), .cin(t_11649), .o(t_11652), .co(t_11653), .cout(t_11654));
half_adder u0_4057(.a(t_10100), .b(t_10097), .o(t_11655), .cout(t_11656));
compressor_4_2 u2_4058(.a(t_10101), .b(t_10098), .c(t_10095), .d(t_7262), .cin(t_11654), .o(t_11657), .co(t_11658), .cout(t_11659));
compressor_3_2 u1_4059(.a(t_10109), .b(t_10106), .cin(t_10103), .o(t_11660), .cout(t_11661));
compressor_4_2 u2_4060(.a(t_10110), .b(t_10107), .c(t_10104), .d(t_7283), .cin(t_11659), .o(t_11662), .co(t_11663), .cout(t_11664));
compressor_3_2 u1_4061(.a(t_10118), .b(t_10115), .cin(t_10112), .o(t_11665), .cout(t_11666));
compressor_4_2 u2_4062(.a(t_10121), .b(t_10119), .c(t_10116), .d(t_10113), .cin(t_11664), .o(t_11667), .co(t_11668), .cout(t_11669));
compressor_3_2 u1_4063(.a(t_10130), .b(t_10127), .cin(t_10124), .o(t_11670), .cout(t_11671));
compressor_4_2 u2_4064(.a(t_10128), .b(t_10125), .c(t_10122), .d(t_7321), .cin(t_11669), .o(t_11672), .co(t_11673), .cout(t_11674));
compressor_3_2 u1_4065(.a(t_10135), .b(t_10132), .cin(t_10131), .o(t_11675), .cout(t_11676));
compressor_4_2 u2_4066(.a(t_10141), .b(t_10139), .c(t_10136), .d(t_10133), .cin(t_11674), .o(t_11677), .co(t_11678), .cout(t_11679));
compressor_3_2 u1_4067(.a(t_10150), .b(t_10147), .cin(t_10144), .o(t_11680), .cout(t_11681));
compressor_4_2 u2_4068(.a(t_10151), .b(t_10148), .c(t_10145), .d(t_10142), .cin(t_11679), .o(t_11682), .co(t_11683), .cout(t_11684));
compressor_3_2 u1_4069(.a(t_10158), .b(t_10155), .cin(t_10152), .o(t_11685), .cout(t_11686));
compressor_4_2 u2_4070(.a(t_10162), .b(t_10159), .c(t_10156), .d(t_10153), .cin(t_11684), .o(t_11687), .co(t_11688), .cout(t_11689));
compressor_3_2 u1_4071(.a(t_10169), .b(t_10166), .cin(t_10163), .o(t_11690), .cout(t_11691));
compressor_4_2 u2_4072(.a(t_10173), .b(t_10170), .c(t_10167), .d(t_10164), .cin(t_11689), .o(t_11692), .co(t_11693), .cout(t_11694));
compressor_3_2 u1_4073(.a(t_10180), .b(t_10177), .cin(t_10174), .o(t_11695), .cout(t_11696));
compressor_4_2 u2_4074(.a(t_10184), .b(t_10181), .c(t_10178), .d(t_10175), .cin(t_11694), .o(t_11697), .co(t_11698), .cout(t_11699));
compressor_3_2 u1_4075(.a(t_10191), .b(t_10188), .cin(t_10185), .o(t_11700), .cout(t_11701));
compressor_4_2 u2_4076(.a(t_10195), .b(t_10192), .c(t_10189), .d(t_10186), .cin(t_11699), .o(t_11702), .co(t_11703), .cout(t_11704));
compressor_3_2 u1_4077(.a(t_10202), .b(t_10199), .cin(t_10196), .o(t_11705), .cout(t_11706));
compressor_4_2 u2_4078(.a(t_10206), .b(t_10203), .c(t_10200), .d(t_10197), .cin(t_11704), .o(t_11707), .co(t_11708), .cout(t_11709));
compressor_3_2 u1_4079(.a(t_10213), .b(t_10210), .cin(t_10207), .o(t_11710), .cout(t_11711));
compressor_4_2 u2_4080(.a(t_10217), .b(t_10214), .c(t_10211), .d(t_10208), .cin(t_11709), .o(t_11712), .co(t_11713), .cout(t_11714));
compressor_3_2 u1_4081(.a(t_10224), .b(t_10221), .cin(t_10218), .o(t_11715), .cout(t_11716));
compressor_4_2 u2_4082(.a(t_10228), .b(t_10225), .c(t_10222), .d(t_10219), .cin(t_11714), .o(t_11717), .co(t_11718), .cout(t_11719));
compressor_3_2 u1_4083(.a(t_10235), .b(t_10232), .cin(t_10229), .o(t_11720), .cout(t_11721));
compressor_4_2 u2_4084(.a(t_10239), .b(t_10236), .c(t_10233), .d(t_10230), .cin(t_11719), .o(t_11722), .co(t_11723), .cout(t_11724));
compressor_3_2 u1_4085(.a(t_10246), .b(t_10243), .cin(t_10240), .o(t_11725), .cout(t_11726));
compressor_4_2 u2_4086(.a(t_10250), .b(t_10247), .c(t_10244), .d(t_10241), .cin(t_11724), .o(t_11727), .co(t_11728), .cout(t_11729));
compressor_3_2 u1_4087(.a(t_10257), .b(t_10254), .cin(t_10251), .o(t_11730), .cout(t_11731));
compressor_4_2 u2_4088(.a(t_10261), .b(t_10258), .c(t_10255), .d(t_10252), .cin(t_11729), .o(t_11732), .co(t_11733), .cout(t_11734));
compressor_3_2 u1_4089(.a(t_10268), .b(t_10265), .cin(t_10262), .o(t_11735), .cout(t_11736));
compressor_4_2 u2_4090(.a(t_10272), .b(t_10269), .c(t_10266), .d(t_10263), .cin(t_11734), .o(t_11737), .co(t_11738), .cout(t_11739));
compressor_3_2 u1_4091(.a(t_10279), .b(t_10276), .cin(t_10273), .o(t_11740), .cout(t_11741));
compressor_4_2 u2_4092(.a(t_10283), .b(t_10280), .c(t_10277), .d(t_10274), .cin(t_11739), .o(t_11742), .co(t_11743), .cout(t_11744));
compressor_3_2 u1_4093(.a(t_10290), .b(t_10287), .cin(t_10284), .o(t_11745), .cout(t_11746));
compressor_4_2 u2_4094(.a(t_10291), .b(t_10288), .c(t_10285), .d(t_7629), .cin(t_11744), .o(t_11747), .co(t_11748), .cout(t_11749));
compressor_4_2 u2_4095(.a(t_10304), .b(t_10301), .c(t_10298), .d(t_10295), .cin(t_10294), .o(t_11750), .co(t_11751), .cout(t_11752));
compressor_4_2 u2_4096(.a(t_10305), .b(t_10302), .c(t_10299), .d(t_10296), .cin(t_11749), .o(t_11753), .co(t_11754), .cout(t_11755));
compressor_4_2 u2_4097(.a(t_10315), .b(t_10312), .c(t_10309), .d(t_10306), .cin(t_11752), .o(t_11756), .co(t_11757), .cout(t_11758));
compressor_4_2 u2_4098(.a(t_10313), .b(t_10310), .c(t_10307), .d(t_7676), .cin(t_11755), .o(t_11759), .co(t_11760), .cout(t_11761));
compressor_4_2 u2_4099(.a(t_10323), .b(t_10320), .c(t_10317), .d(t_10316), .cin(t_11758), .o(t_11762), .co(t_11763), .cout(t_11764));
compressor_4_2 u2_4100(.a(t_10324), .b(t_10321), .c(t_10318), .d(t_7699), .cin(t_11761), .o(t_11765), .co(t_11766), .cout(t_11767));
compressor_4_2 u2_4101(.a(t_10334), .b(t_10331), .c(t_10328), .d(t_10327), .cin(t_11764), .o(t_11768), .co(t_11769), .cout(t_11770));
compressor_4_2 u2_4102(.a(t_10335), .b(t_10332), .c(t_10329), .d(t_7722), .cin(t_11767), .o(t_11771), .co(t_11772), .cout(t_11773));
compressor_4_2 u2_4103(.a(t_10345), .b(t_10342), .c(t_10339), .d(t_10338), .cin(t_11770), .o(t_11774), .co(t_11775), .cout(t_11776));
compressor_4_2 u2_4104(.a(t_10346), .b(t_10343), .c(t_10340), .d(t_7745), .cin(t_11773), .o(t_11777), .co(t_11778), .cout(t_11779));
compressor_4_2 u2_4105(.a(t_10356), .b(t_10353), .c(t_10350), .d(t_10349), .cin(t_11776), .o(t_11780), .co(t_11781), .cout(t_11782));
compressor_4_2 u2_4106(.a(t_10357), .b(t_10354), .c(t_10351), .d(t_7768), .cin(t_11779), .o(t_11783), .co(t_11784), .cout(t_11785));
compressor_4_2 u2_4107(.a(t_10367), .b(t_10364), .c(t_10361), .d(t_10360), .cin(t_11782), .o(t_11786), .co(t_11787), .cout(t_11788));
compressor_4_2 u2_4108(.a(t_10371), .b(t_10368), .c(t_10365), .d(t_10362), .cin(t_11785), .o(t_11789), .co(t_11790), .cout(t_11791));
compressor_4_2 u2_4109(.a(t_10381), .b(t_10378), .c(t_10375), .d(t_10372), .cin(t_11788), .o(t_11792), .co(t_11793), .cout(t_11794));
compressor_4_2 u2_4110(.a(t_10382), .b(t_10379), .c(t_10376), .d(t_10373), .cin(t_11791), .o(t_11795), .co(t_11796), .cout(t_11797));
compressor_4_2 u2_4111(.a(t_10393), .b(t_10390), .c(t_10387), .d(t_10384), .cin(t_11794), .o(t_11798), .co(t_11799), .cout(t_11800));
compressor_4_2 u2_4112(.a(t_10391), .b(t_10388), .c(t_10385), .d(t_7837), .cin(t_11797), .o(t_11801), .co(t_11802), .cout(t_11803));
compressor_4_2 u2_4113(.a(t_10402), .b(t_10399), .c(t_10396), .d(t_10394), .cin(t_11800), .o(t_11804), .co(t_11805), .cout(t_11806));
compressor_4_2 u2_4114(.a(t_10406), .b(t_10403), .c(t_10400), .d(t_10397), .cin(t_11803), .o(t_11807), .co(t_11808), .cout(t_11809));
compressor_4_2 u2_4115(.a(t_10417), .b(t_10414), .c(t_10411), .d(t_10408), .cin(t_11806), .o(t_11810), .co(t_11811), .cout(t_11812));
compressor_4_2 u2_4116(.a(t_10418), .b(t_10415), .c(t_10412), .d(t_10409), .cin(t_11809), .o(t_11813), .co(t_11814), .cout(t_11815));
compressor_4_2 u2_4117(.a(t_10429), .b(t_10426), .c(t_10423), .d(t_10420), .cin(t_11812), .o(t_11816), .co(t_11817), .cout(t_11818));
compressor_4_2 u2_4118(.a(t_10430), .b(t_10427), .c(t_10424), .d(t_10421), .cin(t_11815), .o(t_11819), .co(t_11820), .cout(t_11821));
compressor_4_2 u2_4119(.a(t_10441), .b(t_10438), .c(t_10435), .d(t_10432), .cin(t_11818), .o(t_11822), .co(t_11823), .cout(t_11824));
compressor_4_2 u2_4120(.a(t_10442), .b(t_10439), .c(t_10436), .d(t_10433), .cin(t_11821), .o(t_11825), .co(t_11826), .cout(t_11827));
compressor_4_2 u2_4121(.a(t_10453), .b(t_10450), .c(t_10447), .d(t_10444), .cin(t_11824), .o(t_11828), .co(t_11829), .cout(t_11830));
compressor_4_2 u2_4122(.a(t_10451), .b(t_10448), .c(t_10445), .d(t_7956), .cin(t_11827), .o(t_11831), .co(t_11832), .cout(t_11833));
compressor_4_2 u2_4123(.a(t_10462), .b(t_10459), .c(t_10456), .d(t_10454), .cin(t_11830), .o(t_11834), .co(t_11835), .cout(t_11836));
compressor_4_2 u2_4124(.a(t_10463), .b(t_10460), .c(t_10457), .d(t_7980), .cin(t_11833), .o(t_11837), .co(t_11838), .cout(t_11839));
compressor_4_2 u2_4125(.a(t_10474), .b(t_10471), .c(t_10468), .d(t_10466), .cin(t_11836), .o(t_11840), .co(t_11841), .cout(t_11842));
compressor_4_2 u2_4126(.a(t_10478), .b(t_10475), .c(t_10472), .d(t_10469), .cin(t_11839), .o(t_11843), .co(t_11844), .cout(t_11845));
compressor_4_2 u2_4127(.a(t_10489), .b(t_10486), .c(t_10483), .d(t_10480), .cin(t_11842), .o(t_11846), .co(t_11847), .cout(t_11848));
compressor_4_2 u2_4128(.a(t_10490), .b(t_10487), .c(t_10484), .d(t_10481), .cin(t_11845), .o(t_11849), .co(t_11850), .cout(t_11851));
compressor_4_2 u2_4129(.a(t_10501), .b(t_10498), .c(t_10495), .d(t_10492), .cin(t_11848), .o(t_11852), .co(t_11853), .cout(t_11854));
compressor_4_2 u2_4130(.a(t_10499), .b(t_10496), .c(t_10493), .d(t_8052), .cin(t_11851), .o(t_11855), .co(t_11856), .cout(t_11857));
compressor_4_2 u2_4131(.a(t_10510), .b(t_10507), .c(t_10504), .d(t_10502), .cin(t_11854), .o(t_11858), .co(t_11859), .cout(t_11860));
compressor_4_2 u2_4132(.a(t_10514), .b(t_10511), .c(t_10508), .d(t_10505), .cin(t_11857), .o(t_11861), .co(t_11862), .cout(t_11863));
compressor_4_2 u2_4133(.a(t_10525), .b(t_10522), .c(t_10519), .d(t_10516), .cin(t_11860), .o(t_11864), .co(t_11865), .cout(t_11866));
compressor_4_2 u2_4134(.a(t_10526), .b(t_10523), .c(t_10520), .d(t_10517), .cin(t_11863), .o(t_11867), .co(t_11868), .cout(t_11869));
compressor_4_2 u2_4135(.a(t_10537), .b(t_10534), .c(t_10531), .d(t_10528), .cin(t_11866), .o(t_11870), .co(t_11871), .cout(t_11872));
compressor_4_2 u2_4136(.a(t_10538), .b(t_10535), .c(t_10532), .d(t_10529), .cin(t_11869), .o(t_11873), .co(t_11874), .cout(t_11875));
compressor_4_2 u2_4137(.a(t_10549), .b(t_10546), .c(t_10543), .d(t_10540), .cin(t_11872), .o(t_11876), .co(t_11877), .cout(t_11878));
compressor_4_2 u2_4138(.a(t_10550), .b(t_10547), .c(t_10544), .d(t_10541), .cin(t_11875), .o(t_11879), .co(t_11880), .cout(t_11881));
compressor_4_2 u2_4139(.a(t_10561), .b(t_10558), .c(t_10555), .d(t_10552), .cin(t_11878), .o(t_11882), .co(t_11883), .cout(t_11884));
compressor_4_2 u2_4140(.a(t_10559), .b(t_10556), .c(t_10553), .d(t_8172), .cin(t_11881), .o(t_11885), .co(t_11886), .cout(t_11887));
compressor_4_2 u2_4141(.a(t_10570), .b(t_10567), .c(t_10564), .d(t_10562), .cin(t_11884), .o(t_11888), .co(t_11889), .cout(t_11890));
compressor_4_2 u2_4142(.a(t_10574), .b(t_10571), .c(t_10568), .d(t_10565), .cin(t_11887), .o(t_11891), .co(t_11892), .cout(t_11893));
compressor_4_2 u2_4143(.a(t_10585), .b(t_10582), .c(t_10579), .d(t_10576), .cin(t_11890), .o(t_11894), .co(t_11895), .cout(t_11896));
compressor_4_2 u2_4144(.a(t_10586), .b(t_10583), .c(t_10580), .d(t_10577), .cin(t_11893), .o(t_11897), .co(t_11898), .cout(t_11899));
compressor_4_2 u2_4145(.a(t_10597), .b(t_10594), .c(t_10591), .d(t_10588), .cin(t_11896), .o(t_11900), .co(t_11901), .cout(t_11902));
compressor_4_2 u2_4146(.a(t_10598), .b(t_10595), .c(t_10592), .d(t_10589), .cin(t_11899), .o(t_11903), .co(t_11904), .cout(t_11905));
compressor_4_2 u2_4147(.a(t_10609), .b(t_10606), .c(t_10603), .d(t_10600), .cin(t_11902), .o(t_11906), .co(t_11907), .cout(t_11908));
compressor_4_2 u2_4148(.a(t_10610), .b(t_10607), .c(t_10604), .d(t_10601), .cin(t_11905), .o(t_11909), .co(t_11910), .cout(t_11911));
compressor_4_2 u2_4149(.a(t_10621), .b(t_10618), .c(t_10615), .d(t_10612), .cin(t_11908), .o(t_11912), .co(t_11913), .cout(t_11914));
compressor_4_2 u2_4150(.a(t_10622), .b(t_10619), .c(t_10616), .d(t_10613), .cin(t_11911), .o(t_11915), .co(t_11916), .cout(t_11917));
compressor_4_2 u2_4151(.a(t_10633), .b(t_10630), .c(t_10627), .d(t_10624), .cin(t_11914), .o(t_11918), .co(t_11919), .cout(t_11920));
compressor_4_2 u2_4152(.a(t_10634), .b(t_10631), .c(t_10628), .d(t_10625), .cin(t_11917), .o(t_11921), .co(t_11922), .cout(t_11923));
compressor_4_2 u2_4153(.a(t_10645), .b(t_10642), .c(t_10639), .d(t_10636), .cin(t_11920), .o(t_11924), .co(t_11925), .cout(t_11926));
compressor_4_2 u2_4154(.a(t_10646), .b(t_10643), .c(t_10640), .d(t_10637), .cin(t_11923), .o(t_11927), .co(t_11928), .cout(t_11929));
compressor_4_2 u2_4155(.a(t_10657), .b(t_10654), .c(t_10651), .d(t_10648), .cin(t_11926), .o(t_11930), .co(t_11931), .cout(t_11932));
compressor_4_2 u2_4156(.a(t_10658), .b(t_10655), .c(t_10652), .d(t_10649), .cin(t_11929), .o(t_11933), .co(t_11934), .cout(t_11935));
compressor_4_2 u2_4157(.a(t_10669), .b(t_10666), .c(t_10663), .d(t_10660), .cin(t_11932), .o(t_11936), .co(t_11937), .cout(t_11938));
compressor_4_2 u2_4158(.a(t_10670), .b(t_10667), .c(t_10664), .d(t_10661), .cin(t_11935), .o(t_11939), .co(t_11940), .cout(t_11941));
compressor_4_2 u2_4159(.a(t_10681), .b(t_10678), .c(t_10675), .d(t_10672), .cin(t_11938), .o(t_11942), .co(t_11943), .cout(t_11944));
compressor_4_2 u2_4160(.a(t_10682), .b(t_10679), .c(t_10676), .d(t_10673), .cin(t_11941), .o(t_11945), .co(t_11946), .cout(t_11947));
compressor_4_2 u2_4161(.a(t_10692), .b(t_10689), .c(t_10686), .d(t_10683), .cin(t_11944), .o(t_11948), .co(t_11949), .cout(t_11950));
compressor_4_2 u2_4162(.a(t_10693), .b(t_10690), .c(t_10687), .d(t_10684), .cin(t_11947), .o(t_11951), .co(t_11952), .cout(t_11953));
compressor_4_2 u2_4163(.a(t_10703), .b(t_10700), .c(t_10697), .d(t_10694), .cin(t_11950), .o(t_11954), .co(t_11955), .cout(t_11956));
compressor_4_2 u2_4164(.a(t_10704), .b(t_10701), .c(t_10698), .d(t_10695), .cin(t_11953), .o(t_11957), .co(t_11958), .cout(t_11959));
compressor_4_2 u2_4165(.a(t_10714), .b(t_10711), .c(t_10708), .d(t_10705), .cin(t_11956), .o(t_11960), .co(t_11961), .cout(t_11962));
compressor_4_2 u2_4166(.a(t_10715), .b(t_10712), .c(t_10709), .d(t_10706), .cin(t_11959), .o(t_11963), .co(t_11964), .cout(t_11965));
compressor_4_2 u2_4167(.a(t_10725), .b(t_10722), .c(t_10719), .d(t_10716), .cin(t_11962), .o(t_11966), .co(t_11967), .cout(t_11968));
compressor_4_2 u2_4168(.a(t_10726), .b(t_10723), .c(t_10720), .d(t_10717), .cin(t_11965), .o(t_11969), .co(t_11970), .cout(t_11971));
compressor_4_2 u2_4169(.a(t_10736), .b(t_10733), .c(t_10730), .d(t_10727), .cin(t_11968), .o(t_11972), .co(t_11973), .cout(t_11974));
compressor_4_2 u2_4170(.a(t_10737), .b(t_10734), .c(t_10731), .d(t_10728), .cin(t_11971), .o(t_11975), .co(t_11976), .cout(t_11977));
compressor_4_2 u2_4171(.a(t_10747), .b(t_10744), .c(t_10741), .d(t_10738), .cin(t_11974), .o(t_11978), .co(t_11979), .cout(t_11980));
compressor_4_2 u2_4172(.a(t_10748), .b(t_10745), .c(t_10742), .d(t_10739), .cin(t_11977), .o(t_11981), .co(t_11982), .cout(t_11983));
compressor_4_2 u2_4173(.a(t_10758), .b(t_10755), .c(t_10752), .d(t_10749), .cin(t_11980), .o(t_11984), .co(t_11985), .cout(t_11986));
compressor_4_2 u2_4174(.a(t_10759), .b(t_10756), .c(t_10753), .d(t_10750), .cin(t_11983), .o(t_11987), .co(t_11988), .cout(t_11989));
compressor_4_2 u2_4175(.a(t_10769), .b(t_10766), .c(t_10763), .d(t_10760), .cin(t_11986), .o(t_11990), .co(t_11991), .cout(t_11992));
compressor_4_2 u2_4176(.a(t_10770), .b(t_10767), .c(t_10764), .d(t_10761), .cin(t_11989), .o(t_11993), .co(t_11994), .cout(t_11995));
compressor_4_2 u2_4177(.a(t_10780), .b(t_10777), .c(t_10774), .d(t_10771), .cin(t_11992), .o(t_11996), .co(t_11997), .cout(t_11998));
compressor_4_2 u2_4178(.a(t_10781), .b(t_10778), .c(t_10775), .d(t_10772), .cin(t_11995), .o(t_11999), .co(t_12000), .cout(t_12001));
compressor_4_2 u2_4179(.a(t_10791), .b(t_10788), .c(t_10785), .d(t_10782), .cin(t_11998), .o(t_12002), .co(t_12003), .cout(t_12004));
compressor_4_2 u2_4180(.a(t_10792), .b(t_10789), .c(t_10786), .d(t_10783), .cin(t_12001), .o(t_12005), .co(t_12006), .cout(t_12007));
compressor_4_2 u2_4181(.a(t_10802), .b(t_10799), .c(t_10796), .d(t_10793), .cin(t_12004), .o(t_12008), .co(t_12009), .cout(t_12010));
compressor_4_2 u2_4182(.a(t_10803), .b(t_10800), .c(t_10797), .d(t_10794), .cin(t_12007), .o(t_12011), .co(t_12012), .cout(t_12013));
compressor_4_2 u2_4183(.a(t_10813), .b(t_10810), .c(t_10807), .d(t_10804), .cin(t_12010), .o(t_12014), .co(t_12015), .cout(t_12016));
compressor_4_2 u2_4184(.a(t_10814), .b(t_10811), .c(t_10808), .d(t_10805), .cin(t_12013), .o(t_12017), .co(t_12018), .cout(t_12019));
compressor_4_2 u2_4185(.a(t_10824), .b(t_10821), .c(t_10818), .d(t_10815), .cin(t_12016), .o(t_12020), .co(t_12021), .cout(t_12022));
compressor_4_2 u2_4186(.a(t_10825), .b(t_10822), .c(t_10819), .d(t_10816), .cin(t_12019), .o(t_12023), .co(t_12024), .cout(t_12025));
compressor_4_2 u2_4187(.a(t_10835), .b(t_10832), .c(t_10829), .d(t_10826), .cin(t_12022), .o(t_12026), .co(t_12027), .cout(t_12028));
compressor_4_2 u2_4188(.a(t_10836), .b(t_10833), .c(t_10830), .d(t_10827), .cin(t_12025), .o(t_12029), .co(t_12030), .cout(t_12031));
compressor_4_2 u2_4189(.a(t_10846), .b(t_10843), .c(t_10840), .d(t_10837), .cin(t_12028), .o(t_12032), .co(t_12033), .cout(t_12034));
compressor_4_2 u2_4190(.a(t_10847), .b(t_10844), .c(t_10841), .d(t_10838), .cin(t_12031), .o(t_12035), .co(t_12036), .cout(t_12037));
compressor_3_2 u1_4191(.a(t_10851), .b(t_10848), .cin(t_12034), .o(t_12038), .cout(t_12039));
compressor_4_2 u2_4192(.a(t_10857), .b(t_10855), .c(t_10852), .d(t_10849), .cin(t_12037), .o(t_12040), .co(t_12041), .cout(t_12042));
half_adder u0_4193(.a(t_10863), .b(t_10860), .o(t_12043), .cout(t_12044));
compressor_4_2 u2_4194(.a(t_10864), .b(t_10861), .c(t_10858), .d(t_8732), .cin(t_12042), .o(t_12045), .co(t_12046), .cout(t_12047));
compressor_3_2 u1_4195(.a(t_10872), .b(t_10869), .cin(t_10866), .o(t_12048), .cout(t_12049));
compressor_4_2 u2_4196(.a(t_10875), .b(t_10873), .c(t_10870), .d(t_10867), .cin(t_12047), .o(t_12050), .co(t_12051), .cout(t_12052));
half_adder u0_4197(.a(t_10881), .b(t_10878), .o(t_12053), .cout(t_12054));
compressor_4_2 u2_4198(.a(t_10884), .b(t_10882), .c(t_10879), .d(t_10876), .cin(t_12052), .o(t_12055), .co(t_12056), .cout(t_12057));
half_adder u0_4199(.a(t_10890), .b(t_10887), .o(t_12058), .cout(t_12059));
compressor_4_2 u2_4200(.a(t_10893), .b(t_10891), .c(t_10888), .d(t_10885), .cin(t_12057), .o(t_12060), .co(t_12061), .cout(t_12062));
half_adder u0_4201(.a(t_10899), .b(t_10896), .o(t_12063), .cout(t_12064));
compressor_4_2 u2_4202(.a(t_10902), .b(t_10900), .c(t_10897), .d(t_10894), .cin(t_12062), .o(t_12065), .co(t_12066), .cout(t_12067));
half_adder u0_4203(.a(t_10908), .b(t_10905), .o(t_12068), .cout(t_12069));
compressor_4_2 u2_4204(.a(t_10909), .b(t_10906), .c(t_10903), .d(t_8822), .cin(t_12067), .o(t_12070), .co(t_12071), .cout(t_12072));
compressor_3_2 u1_4205(.a(t_10917), .b(t_10914), .cin(t_10911), .o(t_12073), .cout(t_12074));
compressor_4_2 u2_4206(.a(t_10920), .b(t_10918), .c(t_10915), .d(t_10912), .cin(t_12072), .o(t_12075), .co(t_12076), .cout(t_12077));
half_adder u0_4207(.a(t_10926), .b(t_10923), .o(t_12078), .cout(t_12079));
compressor_4_2 u2_4208(.a(t_10929), .b(t_10927), .c(t_10924), .d(t_10921), .cin(t_12077), .o(t_12080), .co(t_12081), .cout(t_12082));
half_adder u0_4209(.a(t_10935), .b(t_10932), .o(t_12083), .cout(t_12084));
compressor_4_2 u2_4210(.a(t_10938), .b(t_10936), .c(t_10933), .d(t_10930), .cin(t_12082), .o(t_12085), .co(t_12086), .cout(t_12087));
half_adder u0_4211(.a(t_10944), .b(t_10941), .o(t_12088), .cout(t_12089));
compressor_4_2 u2_4212(.a(t_10947), .b(t_10945), .c(t_10942), .d(t_10939), .cin(t_12087), .o(t_12090), .co(t_12091), .cout(t_12092));
half_adder u0_4213(.a(t_10953), .b(t_10950), .o(t_12093), .cout(t_12094));
compressor_4_2 u2_4214(.a(t_10956), .b(t_10954), .c(t_10951), .d(t_10948), .cin(t_12092), .o(t_12095), .co(t_12096), .cout(t_12097));
half_adder u0_4215(.a(t_10962), .b(t_10959), .o(t_12098), .cout(t_12099));
compressor_4_2 u2_4216(.a(t_10965), .b(t_10963), .c(t_10960), .d(t_10957), .cin(t_12097), .o(t_12100), .co(t_12101), .cout(t_12102));
half_adder u0_4217(.a(t_10971), .b(t_10968), .o(t_12103), .cout(t_12104));
compressor_4_2 u2_4218(.a(t_10974), .b(t_10972), .c(t_10969), .d(t_10966), .cin(t_12102), .o(t_12105), .co(t_12106), .cout(t_12107));
half_adder u0_4219(.a(t_10980), .b(t_10977), .o(t_12108), .cout(t_12109));
compressor_4_2 u2_4220(.a(t_10983), .b(t_10981), .c(t_10978), .d(t_10975), .cin(t_12107), .o(t_12110), .co(t_12111), .cout(t_12112));
half_adder u0_4221(.a(t_10989), .b(t_10986), .o(t_12113), .cout(t_12114));
compressor_4_2 u2_4222(.a(t_10992), .b(t_10990), .c(t_10987), .d(t_10984), .cin(t_12112), .o(t_12115), .co(t_12116), .cout(t_12117));
half_adder u0_4223(.a(t_10998), .b(t_10995), .o(t_12118), .cout(t_12119));
compressor_4_2 u2_4224(.a(t_11000), .b(t_10999), .c(t_10996), .d(t_10993), .cin(t_12117), .o(t_12120), .co(t_12121), .cout(t_12122));
half_adder u0_4225(.a(t_11006), .b(t_11003), .o(t_12123), .cout(t_12124));
compressor_4_2 u2_4226(.a(t_11008), .b(t_11007), .c(t_11004), .d(t_11001), .cin(t_12122), .o(t_12125), .co(t_12126), .cout(t_12127));
half_adder u0_4227(.a(t_11014), .b(t_11011), .o(t_12128), .cout(t_12129));
compressor_4_2 u2_4228(.a(t_11016), .b(t_11015), .c(t_11012), .d(t_11009), .cin(t_12127), .o(t_12130), .co(t_12131), .cout(t_12132));
half_adder u0_4229(.a(t_11022), .b(t_11019), .o(t_12133), .cout(t_12134));
compressor_4_2 u2_4230(.a(t_11024), .b(t_11023), .c(t_11020), .d(t_11017), .cin(t_12132), .o(t_12135), .co(t_12136), .cout(t_12137));
half_adder u0_4231(.a(t_11030), .b(t_11027), .o(t_12138), .cout(t_12139));
compressor_4_2 u2_4232(.a(t_11032), .b(t_11031), .c(t_11028), .d(t_11025), .cin(t_12137), .o(t_12140), .co(t_12141), .cout(t_12142));
half_adder u0_4233(.a(t_11038), .b(t_11035), .o(t_12143), .cout(t_12144));
compressor_4_2 u2_4234(.a(t_11040), .b(t_11039), .c(t_11036), .d(t_11033), .cin(t_12142), .o(t_12145), .co(t_12146), .cout(t_12147));
half_adder u0_4235(.a(t_11046), .b(t_11043), .o(t_12148), .cout(t_12149));
compressor_4_2 u2_4236(.a(t_11048), .b(t_11047), .c(t_11044), .d(t_11041), .cin(t_12147), .o(t_12150), .co(t_12151), .cout(t_12152));
half_adder u0_4237(.a(t_11054), .b(t_11051), .o(t_12153), .cout(t_12154));
compressor_4_2 u2_4238(.a(t_11056), .b(t_11055), .c(t_11052), .d(t_11049), .cin(t_12152), .o(t_12155), .co(t_12156), .cout(t_12157));
half_adder u0_4239(.a(t_11062), .b(t_11059), .o(t_12158), .cout(t_12159));
compressor_4_2 u2_4240(.a(t_11064), .b(t_11063), .c(t_11060), .d(t_11057), .cin(t_12157), .o(t_12160), .co(t_12161), .cout(t_12162));
half_adder u0_4241(.a(t_11070), .b(t_11067), .o(t_12163), .cout(t_12164));
compressor_4_2 u2_4242(.a(t_11072), .b(t_11071), .c(t_11068), .d(t_11065), .cin(t_12162), .o(t_12165), .co(t_12166), .cout(t_12167));
half_adder u0_4243(.a(t_11078), .b(t_11075), .o(t_12168), .cout(t_12169));
compressor_4_2 u2_4244(.a(t_11080), .b(t_11079), .c(t_11076), .d(t_11073), .cin(t_12167), .o(t_12170), .co(t_12171), .cout(t_12172));
half_adder u0_4245(.a(t_11086), .b(t_11083), .o(t_12173), .cout(t_12174));
compressor_4_2 u2_4246(.a(t_11088), .b(t_11087), .c(t_11084), .d(t_11081), .cin(t_12172), .o(t_12175), .co(t_12176), .cout(t_12177));
half_adder u0_4247(.a(t_11094), .b(t_11091), .o(t_12178), .cout(t_12179));
compressor_4_2 u2_4248(.a(t_11096), .b(t_11095), .c(t_11092), .d(t_11089), .cin(t_12177), .o(t_12180), .co(t_12181), .cout(t_12182));
half_adder u0_4249(.a(t_11102), .b(t_11099), .o(t_12183), .cout(t_12184));
compressor_4_2 u2_4250(.a(t_11104), .b(t_11103), .c(t_11100), .d(t_11097), .cin(t_12182), .o(t_12185), .co(t_12186), .cout(t_12187));
half_adder u0_4251(.a(t_11110), .b(t_11107), .o(t_12188), .cout(t_12189));
compressor_4_2 u2_4252(.a(t_11112), .b(t_11111), .c(t_11108), .d(t_11105), .cin(t_12187), .o(t_12190), .co(t_12191), .cout(t_12192));
half_adder u0_4253(.a(t_11118), .b(t_11115), .o(t_12193), .cout(t_12194));
compressor_4_2 u2_4254(.a(t_11120), .b(t_11119), .c(t_11116), .d(t_11113), .cin(t_12192), .o(t_12195), .co(t_12196), .cout(t_12197));
compressor_4_2 u2_4255(.a(t_11129), .b(t_11126), .c(t_11124), .d(t_11121), .cin(t_12197), .o(t_12198), .co(t_12199), .cout(t_12200));
compressor_4_2 u2_4256(.a(t_11132), .b(t_11130), .c(t_11127), .d(t_9220), .cin(t_12200), .o(t_12201), .co(t_12202), .cout(t_12203));
compressor_4_2 u2_4257(.a(t_11141), .b(t_11138), .c(t_11136), .d(t_11133), .cin(t_12203), .o(t_12204), .co(t_12205), .cout(t_12206));
compressor_4_2 u2_4258(.a(t_11147), .b(t_11144), .c(t_11142), .d(t_11139), .cin(t_12206), .o(t_12207), .co(t_12208), .cout(t_12209));
compressor_4_2 u2_4259(.a(t_11153), .b(t_11150), .c(t_11148), .d(t_11145), .cin(t_12209), .o(t_12210), .co(t_12211), .cout(t_12212));
compressor_4_2 u2_4260(.a(t_11159), .b(t_11156), .c(t_11154), .d(t_11151), .cin(t_12212), .o(t_12213), .co(t_12214), .cout(t_12215));
compressor_4_2 u2_4261(.a(t_11162), .b(t_11160), .c(t_11157), .d(t_9280), .cin(t_12215), .o(t_12216), .co(t_12217), .cout(t_12218));
compressor_4_2 u2_4262(.a(t_11171), .b(t_11168), .c(t_11166), .d(t_11163), .cin(t_12218), .o(t_12219), .co(t_12220), .cout(t_12221));
compressor_4_2 u2_4263(.a(t_11177), .b(t_11174), .c(t_11172), .d(t_11169), .cin(t_12221), .o(t_12222), .co(t_12223), .cout(t_12224));
compressor_4_2 u2_4264(.a(t_11183), .b(t_11180), .c(t_11178), .d(t_11175), .cin(t_12224), .o(t_12225), .co(t_12226), .cout(t_12227));
compressor_4_2 u2_4265(.a(t_11189), .b(t_11186), .c(t_11184), .d(t_11181), .cin(t_12227), .o(t_12228), .co(t_12229), .cout(t_12230));
compressor_4_2 u2_4266(.a(t_11195), .b(t_11192), .c(t_11190), .d(t_11187), .cin(t_12230), .o(t_12231), .co(t_12232), .cout(t_12233));
compressor_4_2 u2_4267(.a(t_11201), .b(t_11198), .c(t_11196), .d(t_11193), .cin(t_12233), .o(t_12234), .co(t_12235), .cout(t_12236));
compressor_4_2 u2_4268(.a(t_11207), .b(t_11204), .c(t_11202), .d(t_11199), .cin(t_12236), .o(t_12237), .co(t_12238), .cout(t_12239));
compressor_4_2 u2_4269(.a(t_11213), .b(t_11210), .c(t_11208), .d(t_11205), .cin(t_12239), .o(t_12240), .co(t_12241), .cout(t_12242));
compressor_4_2 u2_4270(.a(t_11219), .b(t_11216), .c(t_11214), .d(t_11211), .cin(t_12242), .o(t_12243), .co(t_12244), .cout(t_12245));
compressor_4_2 u2_4271(.a(t_11224), .b(t_11221), .c(t_11220), .d(t_11217), .cin(t_12245), .o(t_12246), .co(t_12247), .cout(t_12248));
compressor_4_2 u2_4272(.a(t_11229), .b(t_11226), .c(t_11225), .d(t_11222), .cin(t_12248), .o(t_12249), .co(t_12250), .cout(t_12251));
compressor_4_2 u2_4273(.a(t_11234), .b(t_11231), .c(t_11230), .d(t_11227), .cin(t_12251), .o(t_12252), .co(t_12253), .cout(t_12254));
compressor_4_2 u2_4274(.a(t_11239), .b(t_11236), .c(t_11235), .d(t_11232), .cin(t_12254), .o(t_12255), .co(t_12256), .cout(t_12257));
compressor_4_2 u2_4275(.a(t_11244), .b(t_11241), .c(t_11240), .d(t_11237), .cin(t_12257), .o(t_12258), .co(t_12259), .cout(t_12260));
compressor_4_2 u2_4276(.a(t_11249), .b(t_11246), .c(t_11245), .d(t_11242), .cin(t_12260), .o(t_12261), .co(t_12262), .cout(t_12263));
compressor_4_2 u2_4277(.a(t_11254), .b(t_11251), .c(t_11250), .d(t_11247), .cin(t_12263), .o(t_12264), .co(t_12265), .cout(t_12266));
compressor_4_2 u2_4278(.a(t_11259), .b(t_11256), .c(t_11255), .d(t_11252), .cin(t_12266), .o(t_12267), .co(t_12268), .cout(t_12269));
compressor_4_2 u2_4279(.a(t_11264), .b(t_11261), .c(t_11260), .d(t_11257), .cin(t_12269), .o(t_12270), .co(t_12271), .cout(t_12272));
compressor_4_2 u2_4280(.a(t_11269), .b(t_11266), .c(t_11265), .d(t_11262), .cin(t_12272), .o(t_12273), .co(t_12274), .cout(t_12275));
compressor_4_2 u2_4281(.a(t_11274), .b(t_11271), .c(t_11270), .d(t_11267), .cin(t_12275), .o(t_12276), .co(t_12277), .cout(t_12278));
compressor_4_2 u2_4282(.a(t_11279), .b(t_11276), .c(t_11275), .d(t_11272), .cin(t_12278), .o(t_12279), .co(t_12280), .cout(t_12281));
compressor_4_2 u2_4283(.a(t_11284), .b(t_11281), .c(t_11280), .d(t_11277), .cin(t_12281), .o(t_12282), .co(t_12283), .cout(t_12284));
compressor_4_2 u2_4284(.a(t_11289), .b(t_11286), .c(t_11285), .d(t_11282), .cin(t_12284), .o(t_12285), .co(t_12286), .cout(t_12287));
compressor_4_2 u2_4285(.a(t_11294), .b(t_11291), .c(t_11290), .d(t_11287), .cin(t_12287), .o(t_12288), .co(t_12289), .cout(t_12290));
compressor_3_2 u1_4286(.a(t_11295), .b(t_11292), .cin(t_12290), .o(t_12291), .cout(t_12292));
half_adder u0_4287(.a(t_11299), .b(t_11297), .o(t_12293), .cout(t_12294));
compressor_3_2 u1_4288(.a(t_11302), .b(t_11300), .cin(t_9516), .o(t_12295), .cout(t_12296));
half_adder u0_4289(.a(t_11305), .b(t_11303), .o(t_12297), .cout(t_12298));
half_adder u0_4290(.a(t_11308), .b(t_11306), .o(t_12299), .cout(t_12300));
half_adder u0_4291(.a(t_11311), .b(t_11309), .o(t_12301), .cout(t_12302));
half_adder u0_4292(.a(t_11314), .b(t_11312), .o(t_12303), .cout(t_12304));
compressor_3_2 u1_4293(.a(t_11317), .b(t_11315), .cin(t_9546), .o(t_12305), .cout(t_12306));
half_adder u0_4294(.a(t_11320), .b(t_11318), .o(t_12307), .cout(t_12308));
half_adder u0_4295(.a(t_11323), .b(t_11321), .o(t_12309), .cout(t_12310));
half_adder u0_4296(.a(t_11326), .b(t_11324), .o(t_12311), .cout(t_12312));
half_adder u0_4297(.a(t_11329), .b(t_11327), .o(t_12313), .cout(t_12314));
half_adder u0_4298(.a(t_11332), .b(t_11330), .o(t_12315), .cout(t_12316));
half_adder u0_4299(.a(t_11335), .b(t_11333), .o(t_12317), .cout(t_12318));
half_adder u0_4300(.a(t_11338), .b(t_11336), .o(t_12319), .cout(t_12320));
half_adder u0_4301(.a(t_11341), .b(t_11339), .o(t_12321), .cout(t_12322));
half_adder u0_4302(.a(t_11344), .b(t_11342), .o(t_12323), .cout(t_12324));
half_adder u0_4303(.a(t_11346), .b(t_11345), .o(t_12325), .cout(t_12326));
half_adder u0_4304(.a(t_11348), .b(t_11347), .o(t_12327), .cout(t_12328));
half_adder u0_4305(.a(t_11350), .b(t_11349), .o(t_12329), .cout(t_12330));
half_adder u0_4306(.a(t_11352), .b(t_11351), .o(t_12331), .cout(t_12332));
half_adder u0_4307(.a(t_11354), .b(t_11353), .o(t_12333), .cout(t_12334));
half_adder u0_4308(.a(t_11356), .b(t_11355), .o(t_12335), .cout(t_12336));
half_adder u0_4309(.a(t_11358), .b(t_11357), .o(t_12337), .cout(t_12338));
half_adder u0_4310(.a(t_11360), .b(t_11359), .o(t_12339), .cout(t_12340));
half_adder u0_4311(.a(t_11362), .b(t_11361), .o(t_12341), .cout(t_12342));
half_adder u0_4312(.a(t_11364), .b(t_11363), .o(t_12343), .cout(t_12344));
half_adder u0_4313(.a(t_11366), .b(t_11365), .o(t_12345), .cout(t_12346));
half_adder u0_4314(.a(t_11368), .b(t_11367), .o(t_12347), .cout(t_12348));
half_adder u0_4315(.a(t_11370), .b(t_11369), .o(t_12349), .cout());

/* u0_4316 Output nets */
wire t_12350,  t_12351;
/* u0_4317 Output nets */
wire t_12352,  t_12353;
/* u0_4318 Output nets */
wire t_12354,  t_12355;
/* u0_4319 Output nets */
wire t_12356,  t_12357;
/* u0_4320 Output nets */
wire t_12358,  t_12359;
/* u0_4321 Output nets */
wire t_12360,  t_12361;
/* u0_4322 Output nets */
wire t_12362,  t_12363;
/* u0_4323 Output nets */
wire t_12364,  t_12365;
/* u0_4324 Output nets */
wire t_12366,  t_12367;
/* u0_4325 Output nets */
wire t_12368,  t_12369;
/* u0_4326 Output nets */
wire t_12370,  t_12371;
/* u0_4327 Output nets */
wire t_12372,  t_12373;
/* u0_4328 Output nets */
wire t_12374,  t_12375;
/* u0_4329 Output nets */
wire t_12376,  t_12377;
/* u0_4330 Output nets */
wire t_12378,  t_12379;
/* u0_4331 Output nets */
wire t_12380,  t_12381;
/* u0_4332 Output nets */
wire t_12382,  t_12383;
/* u0_4333 Output nets */
wire t_12384,  t_12385;
/* u0_4334 Output nets */
wire t_12386,  t_12387;
/* u0_4335 Output nets */
wire t_12388,  t_12389;
/* u0_4336 Output nets */
wire t_12390,  t_12391;
/* u0_4337 Output nets */
wire t_12392,  t_12393;
/* u0_4338 Output nets */
wire t_12394,  t_12395;
/* u0_4339 Output nets */
wire t_12396,  t_12397;
/* u0_4340 Output nets */
wire t_12398,  t_12399;
/* u0_4341 Output nets */
wire t_12400,  t_12401;
/* u0_4342 Output nets */
wire t_12402,  t_12403;
/* u0_4343 Output nets */
wire t_12404,  t_12405;
/* u0_4344 Output nets */
wire t_12406,  t_12407;
/* u0_4345 Output nets */
wire t_12408,  t_12409;
/* u1_4346 Output nets */
wire t_12410,  t_12411;
/* u0_4347 Output nets */
wire t_12412,  t_12413;
/* u1_4348 Output nets */
wire t_12414,  t_12415;
/* u1_4349 Output nets */
wire t_12416,  t_12417;
/* u1_4350 Output nets */
wire t_12418,  t_12419;
/* u1_4351 Output nets */
wire t_12420,  t_12421;
/* u1_4352 Output nets */
wire t_12422,  t_12423;
/* u1_4353 Output nets */
wire t_12424,  t_12425;
/* u1_4354 Output nets */
wire t_12426,  t_12427;
/* u1_4355 Output nets */
wire t_12428,  t_12429;
/* u1_4356 Output nets */
wire t_12430,  t_12431;
/* u1_4357 Output nets */
wire t_12432,  t_12433;
/* u1_4358 Output nets */
wire t_12434,  t_12435;
/* u1_4359 Output nets */
wire t_12436,  t_12437;
/* u1_4360 Output nets */
wire t_12438,  t_12439;
/* u0_4361 Output nets */
wire t_12440,  t_12441;
/* u0_4362 Output nets */
wire t_12442,  t_12443;
/* u1_4363 Output nets */
wire t_12444,  t_12445;
/* u1_4364 Output nets */
wire t_12446,  t_12447;
/* u1_4365 Output nets */
wire t_12448,  t_12449;
/* u1_4366 Output nets */
wire t_12450,  t_12451;
/* u1_4367 Output nets */
wire t_12452,  t_12453;
/* u0_4368 Output nets */
wire t_12454,  t_12455;
/* u0_4369 Output nets */
wire t_12456,  t_12457;
/* u1_4370 Output nets */
wire t_12458,  t_12459;
/* u0_4371 Output nets */
wire t_12460,  t_12461;
/* u0_4372 Output nets */
wire t_12462,  t_12463;
/* u0_4373 Output nets */
wire t_12464,  t_12465;
/* u0_4374 Output nets */
wire t_12466,  t_12467;
/* u1_4375 Output nets */
wire t_12468,  t_12469;
/* u1_4376 Output nets */
wire t_12470,  t_12471;
/* u1_4377 Output nets */
wire t_12472,  t_12473;
/* u1_4378 Output nets */
wire t_12474,  t_12475;
/* u1_4379 Output nets */
wire t_12476,  t_12477;
/* u1_4380 Output nets */
wire t_12478,  t_12479;
/* u1_4381 Output nets */
wire t_12480,  t_12481;
/* u1_4382 Output nets */
wire t_12482,  t_12483;
/* u1_4383 Output nets */
wire t_12484,  t_12485;
/* u1_4384 Output nets */
wire t_12486,  t_12487;
/* u1_4385 Output nets */
wire t_12488,  t_12489;
/* u1_4386 Output nets */
wire t_12490,  t_12491;
/* u1_4387 Output nets */
wire t_12492,  t_12493;
/* u1_4388 Output nets */
wire t_12494,  t_12495;
/* u1_4389 Output nets */
wire t_12496,  t_12497;
/* u1_4390 Output nets */
wire t_12498,  t_12499;
/* u1_4391 Output nets */
wire t_12500,  t_12501;
/* u1_4392 Output nets */
wire t_12502,  t_12503;
/* u1_4393 Output nets */
wire t_12504,  t_12505;
/* u1_4394 Output nets */
wire t_12506,  t_12507;
/* u1_4395 Output nets */
wire t_12508,  t_12509;
/* u1_4396 Output nets */
wire t_12510,  t_12511;
/* u1_4397 Output nets */
wire t_12512,  t_12513;
/* u1_4398 Output nets */
wire t_12514,  t_12515;
/* u1_4399 Output nets */
wire t_12516,  t_12517;
/* u1_4400 Output nets */
wire t_12518,  t_12519;
/* u1_4401 Output nets */
wire t_12520,  t_12521;
/* u1_4402 Output nets */
wire t_12522,  t_12523;
/* u1_4403 Output nets */
wire t_12524,  t_12525;
/* u1_4404 Output nets */
wire t_12526,  t_12527;
/* u1_4405 Output nets */
wire t_12528,  t_12529;
/* u1_4406 Output nets */
wire t_12530,  t_12531;
/* u1_4407 Output nets */
wire t_12532,  t_12533;
/* u1_4408 Output nets */
wire t_12534,  t_12535;
/* u1_4409 Output nets */
wire t_12536,  t_12537;
/* u2_4410 Output nets */
wire t_12538,  t_12539,  t_12540;
/* u2_4411 Output nets */
wire t_12541,  t_12542,  t_12543;
/* u2_4412 Output nets */
wire t_12544,  t_12545,  t_12546;
/* u2_4413 Output nets */
wire t_12547,  t_12548,  t_12549;
/* u2_4414 Output nets */
wire t_12550,  t_12551,  t_12552;
/* u2_4415 Output nets */
wire t_12553,  t_12554,  t_12555;
/* u2_4416 Output nets */
wire t_12556,  t_12557,  t_12558;
/* u2_4417 Output nets */
wire t_12559,  t_12560,  t_12561;
/* u2_4418 Output nets */
wire t_12562,  t_12563,  t_12564;
/* u2_4419 Output nets */
wire t_12565,  t_12566,  t_12567;
/* u2_4420 Output nets */
wire t_12568,  t_12569,  t_12570;
/* u2_4421 Output nets */
wire t_12571,  t_12572,  t_12573;
/* u2_4422 Output nets */
wire t_12574,  t_12575,  t_12576;
/* u2_4423 Output nets */
wire t_12577,  t_12578,  t_12579;
/* u2_4424 Output nets */
wire t_12580,  t_12581,  t_12582;
/* u2_4425 Output nets */
wire t_12583,  t_12584,  t_12585;
/* u2_4426 Output nets */
wire t_12586,  t_12587,  t_12588;
/* u2_4427 Output nets */
wire t_12589,  t_12590,  t_12591;
/* u2_4428 Output nets */
wire t_12592,  t_12593,  t_12594;
/* u2_4429 Output nets */
wire t_12595,  t_12596,  t_12597;
/* u2_4430 Output nets */
wire t_12598,  t_12599,  t_12600;
/* u2_4431 Output nets */
wire t_12601,  t_12602,  t_12603;
/* u2_4432 Output nets */
wire t_12604,  t_12605,  t_12606;
/* u2_4433 Output nets */
wire t_12607,  t_12608,  t_12609;
/* u2_4434 Output nets */
wire t_12610,  t_12611,  t_12612;
/* u2_4435 Output nets */
wire t_12613,  t_12614,  t_12615;
/* u2_4436 Output nets */
wire t_12616,  t_12617,  t_12618;
/* u2_4437 Output nets */
wire t_12619,  t_12620,  t_12621;
/* u2_4438 Output nets */
wire t_12622,  t_12623,  t_12624;
/* u2_4439 Output nets */
wire t_12625,  t_12626,  t_12627;
/* u2_4440 Output nets */
wire t_12628,  t_12629,  t_12630;
/* u2_4441 Output nets */
wire t_12631,  t_12632,  t_12633;
/* u2_4442 Output nets */
wire t_12634,  t_12635,  t_12636;
/* u2_4443 Output nets */
wire t_12637,  t_12638,  t_12639;
/* u2_4444 Output nets */
wire t_12640,  t_12641,  t_12642;
/* u2_4445 Output nets */
wire t_12643,  t_12644,  t_12645;
/* u2_4446 Output nets */
wire t_12646,  t_12647,  t_12648;
/* u2_4447 Output nets */
wire t_12649,  t_12650,  t_12651;
/* u2_4448 Output nets */
wire t_12652,  t_12653,  t_12654;
/* u2_4449 Output nets */
wire t_12655,  t_12656,  t_12657;
/* u2_4450 Output nets */
wire t_12658,  t_12659,  t_12660;
/* u2_4451 Output nets */
wire t_12661,  t_12662,  t_12663;
/* u2_4452 Output nets */
wire t_12664,  t_12665,  t_12666;
/* u2_4453 Output nets */
wire t_12667,  t_12668,  t_12669;
/* u2_4454 Output nets */
wire t_12670,  t_12671,  t_12672;
/* u2_4455 Output nets */
wire t_12673,  t_12674,  t_12675;
/* u2_4456 Output nets */
wire t_12676,  t_12677,  t_12678;
/* u2_4457 Output nets */
wire t_12679,  t_12680,  t_12681;
/* u2_4458 Output nets */
wire t_12682,  t_12683,  t_12684;
/* u2_4459 Output nets */
wire t_12685,  t_12686,  t_12687;
/* u2_4460 Output nets */
wire t_12688,  t_12689,  t_12690;
/* u2_4461 Output nets */
wire t_12691,  t_12692,  t_12693;
/* u2_4462 Output nets */
wire t_12694,  t_12695,  t_12696;
/* u2_4463 Output nets */
wire t_12697,  t_12698,  t_12699;
/* u2_4464 Output nets */
wire t_12700,  t_12701,  t_12702;
/* u2_4465 Output nets */
wire t_12703,  t_12704,  t_12705;
/* u2_4466 Output nets */
wire t_12706,  t_12707,  t_12708;
/* u2_4467 Output nets */
wire t_12709,  t_12710,  t_12711;
/* u2_4468 Output nets */
wire t_12712,  t_12713,  t_12714;
/* u2_4469 Output nets */
wire t_12715,  t_12716,  t_12717;
/* u2_4470 Output nets */
wire t_12718,  t_12719,  t_12720;
/* u2_4471 Output nets */
wire t_12721,  t_12722,  t_12723;
/* u2_4472 Output nets */
wire t_12724,  t_12725,  t_12726;
/* u2_4473 Output nets */
wire t_12727,  t_12728,  t_12729;
/* u2_4474 Output nets */
wire t_12730,  t_12731,  t_12732;
/* u2_4475 Output nets */
wire t_12733,  t_12734,  t_12735;
/* u2_4476 Output nets */
wire t_12736,  t_12737,  t_12738;
/* u2_4477 Output nets */
wire t_12739,  t_12740,  t_12741;
/* u2_4478 Output nets */
wire t_12742,  t_12743,  t_12744;
/* u2_4479 Output nets */
wire t_12745,  t_12746,  t_12747;
/* u2_4480 Output nets */
wire t_12748,  t_12749,  t_12750;
/* u2_4481 Output nets */
wire t_12751,  t_12752,  t_12753;
/* u2_4482 Output nets */
wire t_12754,  t_12755,  t_12756;
/* u2_4483 Output nets */
wire t_12757,  t_12758,  t_12759;
/* u2_4484 Output nets */
wire t_12760,  t_12761,  t_12762;
/* u2_4485 Output nets */
wire t_12763,  t_12764,  t_12765;
/* u2_4486 Output nets */
wire t_12766,  t_12767,  t_12768;
/* u2_4487 Output nets */
wire t_12769,  t_12770,  t_12771;
/* u2_4488 Output nets */
wire t_12772,  t_12773,  t_12774;
/* u2_4489 Output nets */
wire t_12775,  t_12776,  t_12777;
/* u2_4490 Output nets */
wire t_12778,  t_12779,  t_12780;
/* u2_4491 Output nets */
wire t_12781,  t_12782,  t_12783;
/* u2_4492 Output nets */
wire t_12784,  t_12785,  t_12786;
/* u2_4493 Output nets */
wire t_12787,  t_12788,  t_12789;
/* u2_4494 Output nets */
wire t_12790,  t_12791,  t_12792;
/* u2_4495 Output nets */
wire t_12793,  t_12794,  t_12795;
/* u2_4496 Output nets */
wire t_12796,  t_12797,  t_12798;
/* u2_4497 Output nets */
wire t_12799,  t_12800,  t_12801;
/* u2_4498 Output nets */
wire t_12802,  t_12803,  t_12804;
/* u2_4499 Output nets */
wire t_12805,  t_12806,  t_12807;
/* u2_4500 Output nets */
wire t_12808,  t_12809,  t_12810;
/* u2_4501 Output nets */
wire t_12811,  t_12812,  t_12813;
/* u2_4502 Output nets */
wire t_12814,  t_12815,  t_12816;
/* u2_4503 Output nets */
wire t_12817,  t_12818,  t_12819;
/* u2_4504 Output nets */
wire t_12820,  t_12821,  t_12822;
/* u2_4505 Output nets */
wire t_12823,  t_12824,  t_12825;
/* u1_4506 Output nets */
wire t_12826,  t_12827;
/* u1_4507 Output nets */
wire t_12828,  t_12829;
/* u0_4508 Output nets */
wire t_12830,  t_12831;
/* u0_4509 Output nets */
wire t_12832,  t_12833;
/* u0_4510 Output nets */
wire t_12834,  t_12835;
/* u0_4511 Output nets */
wire t_12836,  t_12837;
/* u1_4512 Output nets */
wire t_12838,  t_12839;
/* u0_4513 Output nets */
wire t_12840,  t_12841;
/* u0_4514 Output nets */
wire t_12842,  t_12843;
/* u0_4515 Output nets */
wire t_12844,  t_12845;
/* u0_4516 Output nets */
wire t_12846,  t_12847;
/* u0_4517 Output nets */
wire t_12848,  t_12849;
/* u0_4518 Output nets */
wire t_12850,  t_12851;
/* u0_4519 Output nets */
wire t_12852,  t_12853;
/* u0_4520 Output nets */
wire t_12854,  t_12855;
/* u0_4521 Output nets */
wire t_12856,  t_12857;
/* u0_4522 Output nets */
wire t_12858,  t_12859;
/* u0_4523 Output nets */
wire t_12860,  t_12861;
/* u0_4524 Output nets */
wire t_12862,  t_12863;
/* u0_4525 Output nets */
wire t_12864,  t_12865;
/* u0_4526 Output nets */
wire t_12866,  t_12867;
/* u0_4527 Output nets */
wire t_12868,  t_12869;
/* u0_4528 Output nets */
wire t_12870,  t_12871;
/* u0_4529 Output nets */
wire t_12872,  t_12873;
/* u0_4530 Output nets */
wire t_12874,  t_12875;
/* u0_4531 Output nets */
wire t_12876,  t_12877;
/* u0_4532 Output nets */
wire t_12878,  t_12879;
/* u0_4533 Output nets */
wire t_12880,  t_12881;
/* u0_4534 Output nets */
wire t_12882,  t_12883;
/* u0_4535 Output nets */
wire t_12884,  t_12885;
/* u0_4536 Output nets */
wire t_12886,  t_12887;
/* u1_4537 Output nets */
wire t_12888,  t_12889;
/* u0_4538 Output nets */
wire t_12890,  t_12891;
/* u0_4539 Output nets */
wire t_12892,  t_12893;
/* u0_4540 Output nets */
wire t_12894,  t_12895;
/* u0_4541 Output nets */
wire t_12896,  t_12897;
/* u0_4542 Output nets */
wire t_12898,  t_12899;
/* u0_4543 Output nets */
wire t_12900,  t_12901;
/* u0_4544 Output nets */
wire t_12902,  t_12903;
/* u0_4545 Output nets */
wire t_12904,  t_12905;
/* u0_4546 Output nets */
wire t_12906,  t_12907;
/* u0_4547 Output nets */
wire t_12908,  t_12909;
/* u0_4548 Output nets */
wire t_12910,  t_12911;
/* u0_4549 Output nets */
wire t_12912,  t_12913;
/* u0_4550 Output nets */
wire t_12914,  t_12915;
/* u0_4551 Output nets */
wire t_12916,  t_12917;
/* u0_4552 Output nets */
wire t_12918,  t_12919;
/* u0_4553 Output nets */
wire t_12920,  t_12921;
/* u0_4554 Output nets */
wire t_12922,  t_12923;
/* u0_4555 Output nets */
wire t_12924,  t_12925;
/* u0_4556 Output nets */
wire t_12926,  t_12927;
/* u0_4557 Output nets */
wire t_12928,  t_12929;
/* u0_4558 Output nets */
wire t_12930,  t_12931;
/* u0_4559 Output nets */
wire t_12932,  t_12933;
/* u0_4560 Output nets */
wire t_12934,  t_12935;
/* u0_4561 Output nets */
wire t_12936,  t_12937;
/* u0_4562 Output nets */
wire t_12938,  t_12939;
/* u0_4563 Output nets */
wire t_12940,  t_12941;
/* u0_4564 Output nets */
wire t_12942,  t_12943;
/* u0_4565 Output nets */
wire t_12944,  t_12945;
/* u0_4566 Output nets */
wire t_12946;

/* compress stage 5 */
half_adder u0_4316(.a(t_11372), .b(t_9622), .o(t_12350), .cout(t_12351));
half_adder u0_4317(.a(t_11375), .b(t_11374), .o(t_12352), .cout(t_12353));
half_adder u0_4318(.a(t_11377), .b(t_11376), .o(t_12354), .cout(t_12355));
half_adder u0_4319(.a(t_11379), .b(t_11378), .o(t_12356), .cout(t_12357));
half_adder u0_4320(.a(t_11381), .b(t_11380), .o(t_12358), .cout(t_12359));
half_adder u0_4321(.a(t_11383), .b(t_11382), .o(t_12360), .cout(t_12361));
half_adder u0_4322(.a(t_11385), .b(t_11384), .o(t_12362), .cout(t_12363));
half_adder u0_4323(.a(t_11387), .b(t_11386), .o(t_12364), .cout(t_12365));
half_adder u0_4324(.a(t_11389), .b(t_11388), .o(t_12366), .cout(t_12367));
half_adder u0_4325(.a(t_11391), .b(t_11390), .o(t_12368), .cout(t_12369));
half_adder u0_4326(.a(t_11393), .b(t_11392), .o(t_12370), .cout(t_12371));
half_adder u0_4327(.a(t_11395), .b(t_11394), .o(t_12372), .cout(t_12373));
half_adder u0_4328(.a(t_11397), .b(t_11396), .o(t_12374), .cout(t_12375));
half_adder u0_4329(.a(t_11399), .b(t_11398), .o(t_12376), .cout(t_12377));
half_adder u0_4330(.a(t_11401), .b(t_11400), .o(t_12378), .cout(t_12379));
half_adder u0_4331(.a(t_11403), .b(t_11402), .o(t_12380), .cout(t_12381));
half_adder u0_4332(.a(t_11405), .b(t_11404), .o(t_12382), .cout(t_12383));
half_adder u0_4333(.a(t_11407), .b(t_11406), .o(t_12384), .cout(t_12385));
half_adder u0_4334(.a(t_11409), .b(t_11408), .o(t_12386), .cout(t_12387));
half_adder u0_4335(.a(t_11411), .b(t_11410), .o(t_12388), .cout(t_12389));
half_adder u0_4336(.a(t_11413), .b(t_11412), .o(t_12390), .cout(t_12391));
half_adder u0_4337(.a(t_11415), .b(t_11414), .o(t_12392), .cout(t_12393));
half_adder u0_4338(.a(t_11417), .b(t_11416), .o(t_12394), .cout(t_12395));
half_adder u0_4339(.a(t_11419), .b(t_11418), .o(t_12396), .cout(t_12397));
half_adder u0_4340(.a(t_11421), .b(t_11420), .o(t_12398), .cout(t_12399));
half_adder u0_4341(.a(t_11423), .b(t_11422), .o(t_12400), .cout(t_12401));
half_adder u0_4342(.a(t_11425), .b(t_11424), .o(t_12402), .cout(t_12403));
half_adder u0_4343(.a(t_11427), .b(t_11426), .o(t_12404), .cout(t_12405));
half_adder u0_4344(.a(t_11429), .b(t_11428), .o(t_12406), .cout(t_12407));
half_adder u0_4345(.a(t_11431), .b(t_11430), .o(t_12408), .cout(t_12409));
compressor_3_2 u1_4346(.a(t_11433), .b(t_11432), .cin(t_9696), .o(t_12410), .cout(t_12411));
half_adder u0_4347(.a(t_11435), .b(t_11434), .o(t_12412), .cout(t_12413));
compressor_3_2 u1_4348(.a(t_11437), .b(t_11436), .cin(t_9707), .o(t_12414), .cout(t_12415));
compressor_3_2 u1_4349(.a(t_11439), .b(t_11438), .cin(t_9712), .o(t_12416), .cout(t_12417));
compressor_3_2 u1_4350(.a(t_11441), .b(t_11440), .cin(t_9717), .o(t_12418), .cout(t_12419));
compressor_3_2 u1_4351(.a(t_11443), .b(t_11442), .cin(t_9722), .o(t_12420), .cout(t_12421));
compressor_3_2 u1_4352(.a(t_11445), .b(t_11444), .cin(t_9727), .o(t_12422), .cout(t_12423));
compressor_3_2 u1_4353(.a(t_11447), .b(t_11446), .cin(t_9732), .o(t_12424), .cout(t_12425));
compressor_3_2 u1_4354(.a(t_11449), .b(t_11448), .cin(t_9737), .o(t_12426), .cout(t_12427));
compressor_3_2 u1_4355(.a(t_11451), .b(t_11450), .cin(t_9742), .o(t_12428), .cout(t_12429));
compressor_3_2 u1_4356(.a(t_11453), .b(t_11452), .cin(t_9747), .o(t_12430), .cout(t_12431));
compressor_3_2 u1_4357(.a(t_11455), .b(t_11454), .cin(t_9752), .o(t_12432), .cout(t_12433));
compressor_3_2 u1_4358(.a(t_11457), .b(t_11456), .cin(t_9757), .o(t_12434), .cout(t_12435));
compressor_3_2 u1_4359(.a(t_11459), .b(t_11458), .cin(t_9762), .o(t_12436), .cout(t_12437));
compressor_3_2 u1_4360(.a(t_11461), .b(t_11460), .cin(t_9767), .o(t_12438), .cout(t_12439));
half_adder u0_4361(.a(t_11463), .b(t_11462), .o(t_12440), .cout(t_12441));
half_adder u0_4362(.a(t_11466), .b(t_11464), .o(t_12442), .cout(t_12443));
compressor_3_2 u1_4363(.a(t_11469), .b(t_11467), .cin(t_9782), .o(t_12444), .cout(t_12445));
compressor_3_2 u1_4364(.a(t_11472), .b(t_11470), .cin(t_9787), .o(t_12446), .cout(t_12447));
compressor_3_2 u1_4365(.a(t_11475), .b(t_11473), .cin(t_9792), .o(t_12448), .cout(t_12449));
compressor_3_2 u1_4366(.a(t_11478), .b(t_11476), .cin(t_9797), .o(t_12450), .cout(t_12451));
compressor_3_2 u1_4367(.a(t_11481), .b(t_11479), .cin(t_9802), .o(t_12452), .cout(t_12453));
half_adder u0_4368(.a(t_11484), .b(t_11482), .o(t_12454), .cout(t_12455));
half_adder u0_4369(.a(t_11487), .b(t_11485), .o(t_12456), .cout(t_12457));
compressor_3_2 u1_4370(.a(t_11490), .b(t_11488), .cin(t_9819), .o(t_12458), .cout(t_12459));
half_adder u0_4371(.a(t_11493), .b(t_11491), .o(t_12460), .cout(t_12461));
half_adder u0_4372(.a(t_11496), .b(t_11494), .o(t_12462), .cout(t_12463));
half_adder u0_4373(.a(t_11499), .b(t_11497), .o(t_12464), .cout(t_12465));
half_adder u0_4374(.a(t_11502), .b(t_11500), .o(t_12466), .cout(t_12467));
compressor_3_2 u1_4375(.a(t_11505), .b(t_11503), .cin(t_9849), .o(t_12468), .cout(t_12469));
compressor_3_2 u1_4376(.a(t_11508), .b(t_11506), .cin(t_9855), .o(t_12470), .cout(t_12471));
compressor_3_2 u1_4377(.a(t_11511), .b(t_11509), .cin(t_9864), .o(t_12472), .cout(t_12473));
compressor_3_2 u1_4378(.a(t_11517), .b(t_11514), .cin(t_11512), .o(t_12474), .cout(t_12475));
compressor_3_2 u1_4379(.a(t_11518), .b(t_11515), .cin(t_9878), .o(t_12476), .cout(t_12477));
compressor_3_2 u1_4380(.a(t_11525), .b(t_11522), .cin(t_11520), .o(t_12478), .cout(t_12479));
compressor_3_2 u1_4381(.a(t_11527), .b(t_11526), .cin(t_11523), .o(t_12480), .cout(t_12481));
compressor_3_2 u1_4382(.a(t_11532), .b(t_11531), .cin(t_11528), .o(t_12482), .cout(t_12483));
compressor_3_2 u1_4383(.a(t_11537), .b(t_11536), .cin(t_11533), .o(t_12484), .cout(t_12485));
compressor_3_2 u1_4384(.a(t_11542), .b(t_11541), .cin(t_11538), .o(t_12486), .cout(t_12487));
compressor_3_2 u1_4385(.a(t_11547), .b(t_11546), .cin(t_11543), .o(t_12488), .cout(t_12489));
compressor_3_2 u1_4386(.a(t_11552), .b(t_11551), .cin(t_11548), .o(t_12490), .cout(t_12491));
compressor_3_2 u1_4387(.a(t_11557), .b(t_11556), .cin(t_11553), .o(t_12492), .cout(t_12493));
compressor_3_2 u1_4388(.a(t_11562), .b(t_11561), .cin(t_11558), .o(t_12494), .cout(t_12495));
compressor_3_2 u1_4389(.a(t_11567), .b(t_11566), .cin(t_11563), .o(t_12496), .cout(t_12497));
compressor_3_2 u1_4390(.a(t_11572), .b(t_11571), .cin(t_11568), .o(t_12498), .cout(t_12499));
compressor_3_2 u1_4391(.a(t_11577), .b(t_11576), .cin(t_11573), .o(t_12500), .cout(t_12501));
compressor_3_2 u1_4392(.a(t_11582), .b(t_11581), .cin(t_11578), .o(t_12502), .cout(t_12503));
compressor_3_2 u1_4393(.a(t_11587), .b(t_11586), .cin(t_11583), .o(t_12504), .cout(t_12505));
compressor_3_2 u1_4394(.a(t_11592), .b(t_11591), .cin(t_11588), .o(t_12506), .cout(t_12507));
compressor_3_2 u1_4395(.a(t_11597), .b(t_11596), .cin(t_11593), .o(t_12508), .cout(t_12509));
compressor_3_2 u1_4396(.a(t_11602), .b(t_11601), .cin(t_11598), .o(t_12510), .cout(t_12511));
compressor_3_2 u1_4397(.a(t_11607), .b(t_11606), .cin(t_11603), .o(t_12512), .cout(t_12513));
compressor_3_2 u1_4398(.a(t_11612), .b(t_11611), .cin(t_11608), .o(t_12514), .cout(t_12515));
compressor_3_2 u1_4399(.a(t_11617), .b(t_11616), .cin(t_11613), .o(t_12516), .cout(t_12517));
compressor_3_2 u1_4400(.a(t_11622), .b(t_11621), .cin(t_11618), .o(t_12518), .cout(t_12519));
compressor_3_2 u1_4401(.a(t_11627), .b(t_11626), .cin(t_11623), .o(t_12520), .cout(t_12521));
compressor_3_2 u1_4402(.a(t_11632), .b(t_11631), .cin(t_11628), .o(t_12522), .cout(t_12523));
compressor_3_2 u1_4403(.a(t_11637), .b(t_11636), .cin(t_11633), .o(t_12524), .cout(t_12525));
compressor_3_2 u1_4404(.a(t_11642), .b(t_11641), .cin(t_11638), .o(t_12526), .cout(t_12527));
compressor_3_2 u1_4405(.a(t_11647), .b(t_11646), .cin(t_11643), .o(t_12528), .cout(t_12529));
compressor_3_2 u1_4406(.a(t_11652), .b(t_11651), .cin(t_11648), .o(t_12530), .cout(t_12531));
compressor_3_2 u1_4407(.a(t_11657), .b(t_11656), .cin(t_11653), .o(t_12532), .cout(t_12533));
compressor_3_2 u1_4408(.a(t_11662), .b(t_11661), .cin(t_11658), .o(t_12534), .cout(t_12535));
compressor_3_2 u1_4409(.a(t_11667), .b(t_11666), .cin(t_11663), .o(t_12536), .cout(t_12537));
compressor_4_2 u2_4410(.a(t_11675), .b(t_11672), .c(t_11671), .d(t_11668), .cin(t_10138), .o(t_12538), .co(t_12539), .cout(t_12540));
compressor_4_2 u2_4411(.a(t_11680), .b(t_11677), .c(t_11676), .d(t_11673), .cin(t_12540), .o(t_12541), .co(t_12542), .cout(t_12543));
compressor_4_2 u2_4412(.a(t_11682), .b(t_11681), .c(t_11678), .d(t_10161), .cin(t_12543), .o(t_12544), .co(t_12545), .cout(t_12546));
compressor_4_2 u2_4413(.a(t_11687), .b(t_11686), .c(t_11683), .d(t_10172), .cin(t_12546), .o(t_12547), .co(t_12548), .cout(t_12549));
compressor_4_2 u2_4414(.a(t_11692), .b(t_11691), .c(t_11688), .d(t_10183), .cin(t_12549), .o(t_12550), .co(t_12551), .cout(t_12552));
compressor_4_2 u2_4415(.a(t_11697), .b(t_11696), .c(t_11693), .d(t_10194), .cin(t_12552), .o(t_12553), .co(t_12554), .cout(t_12555));
compressor_4_2 u2_4416(.a(t_11702), .b(t_11701), .c(t_11698), .d(t_10205), .cin(t_12555), .o(t_12556), .co(t_12557), .cout(t_12558));
compressor_4_2 u2_4417(.a(t_11707), .b(t_11706), .c(t_11703), .d(t_10216), .cin(t_12558), .o(t_12559), .co(t_12560), .cout(t_12561));
compressor_4_2 u2_4418(.a(t_11712), .b(t_11711), .c(t_11708), .d(t_10227), .cin(t_12561), .o(t_12562), .co(t_12563), .cout(t_12564));
compressor_4_2 u2_4419(.a(t_11717), .b(t_11716), .c(t_11713), .d(t_10238), .cin(t_12564), .o(t_12565), .co(t_12566), .cout(t_12567));
compressor_4_2 u2_4420(.a(t_11722), .b(t_11721), .c(t_11718), .d(t_10249), .cin(t_12567), .o(t_12568), .co(t_12569), .cout(t_12570));
compressor_4_2 u2_4421(.a(t_11727), .b(t_11726), .c(t_11723), .d(t_10260), .cin(t_12570), .o(t_12571), .co(t_12572), .cout(t_12573));
compressor_4_2 u2_4422(.a(t_11732), .b(t_11731), .c(t_11728), .d(t_10271), .cin(t_12573), .o(t_12574), .co(t_12575), .cout(t_12576));
compressor_4_2 u2_4423(.a(t_11737), .b(t_11736), .c(t_11733), .d(t_10282), .cin(t_12576), .o(t_12577), .co(t_12578), .cout(t_12579));
compressor_4_2 u2_4424(.a(t_11742), .b(t_11741), .c(t_11738), .d(t_10293), .cin(t_12579), .o(t_12580), .co(t_12581), .cout(t_12582));
compressor_4_2 u2_4425(.a(t_11750), .b(t_11747), .c(t_11746), .d(t_11743), .cin(t_12582), .o(t_12583), .co(t_12584), .cout(t_12585));
compressor_4_2 u2_4426(.a(t_11756), .b(t_11753), .c(t_11751), .d(t_11748), .cin(t_12585), .o(t_12586), .co(t_12587), .cout(t_12588));
compressor_4_2 u2_4427(.a(t_11759), .b(t_11757), .c(t_11754), .d(t_10326), .cin(t_12588), .o(t_12589), .co(t_12590), .cout(t_12591));
compressor_4_2 u2_4428(.a(t_11765), .b(t_11763), .c(t_11760), .d(t_10337), .cin(t_12591), .o(t_12592), .co(t_12593), .cout(t_12594));
compressor_4_2 u2_4429(.a(t_11771), .b(t_11769), .c(t_11766), .d(t_10348), .cin(t_12594), .o(t_12595), .co(t_12596), .cout(t_12597));
compressor_4_2 u2_4430(.a(t_11777), .b(t_11775), .c(t_11772), .d(t_10359), .cin(t_12597), .o(t_12598), .co(t_12599), .cout(t_12600));
compressor_4_2 u2_4431(.a(t_11783), .b(t_11781), .c(t_11778), .d(t_10370), .cin(t_12600), .o(t_12601), .co(t_12602), .cout(t_12603));
compressor_4_2 u2_4432(.a(t_11792), .b(t_11789), .c(t_11787), .d(t_11784), .cin(t_12603), .o(t_12604), .co(t_12605), .cout(t_12606));
compressor_4_2 u2_4433(.a(t_11798), .b(t_11795), .c(t_11793), .d(t_11790), .cin(t_12606), .o(t_12607), .co(t_12608), .cout(t_12609));
compressor_4_2 u2_4434(.a(t_11801), .b(t_11799), .c(t_11796), .d(t_10405), .cin(t_12609), .o(t_12610), .co(t_12611), .cout(t_12612));
compressor_4_2 u2_4435(.a(t_11810), .b(t_11807), .c(t_11805), .d(t_11802), .cin(t_12612), .o(t_12613), .co(t_12614), .cout(t_12615));
compressor_4_2 u2_4436(.a(t_11816), .b(t_11813), .c(t_11811), .d(t_11808), .cin(t_12615), .o(t_12616), .co(t_12617), .cout(t_12618));
compressor_4_2 u2_4437(.a(t_11822), .b(t_11819), .c(t_11817), .d(t_11814), .cin(t_12618), .o(t_12619), .co(t_12620), .cout(t_12621));
compressor_4_2 u2_4438(.a(t_11828), .b(t_11825), .c(t_11823), .d(t_11820), .cin(t_12621), .o(t_12622), .co(t_12623), .cout(t_12624));
compressor_4_2 u2_4439(.a(t_11831), .b(t_11829), .c(t_11826), .d(t_10465), .cin(t_12624), .o(t_12625), .co(t_12626), .cout(t_12627));
compressor_4_2 u2_4440(.a(t_11837), .b(t_11835), .c(t_11832), .d(t_10477), .cin(t_12627), .o(t_12628), .co(t_12629), .cout(t_12630));
compressor_4_2 u2_4441(.a(t_11846), .b(t_11843), .c(t_11841), .d(t_11838), .cin(t_12630), .o(t_12631), .co(t_12632), .cout(t_12633));
compressor_4_2 u2_4442(.a(t_11852), .b(t_11849), .c(t_11847), .d(t_11844), .cin(t_12633), .o(t_12634), .co(t_12635), .cout(t_12636));
compressor_4_2 u2_4443(.a(t_11855), .b(t_11853), .c(t_11850), .d(t_10513), .cin(t_12636), .o(t_12637), .co(t_12638), .cout(t_12639));
compressor_4_2 u2_4444(.a(t_11864), .b(t_11861), .c(t_11859), .d(t_11856), .cin(t_12639), .o(t_12640), .co(t_12641), .cout(t_12642));
compressor_4_2 u2_4445(.a(t_11870), .b(t_11867), .c(t_11865), .d(t_11862), .cin(t_12642), .o(t_12643), .co(t_12644), .cout(t_12645));
compressor_4_2 u2_4446(.a(t_11876), .b(t_11873), .c(t_11871), .d(t_11868), .cin(t_12645), .o(t_12646), .co(t_12647), .cout(t_12648));
compressor_4_2 u2_4447(.a(t_11882), .b(t_11879), .c(t_11877), .d(t_11874), .cin(t_12648), .o(t_12649), .co(t_12650), .cout(t_12651));
compressor_4_2 u2_4448(.a(t_11885), .b(t_11883), .c(t_11880), .d(t_10573), .cin(t_12651), .o(t_12652), .co(t_12653), .cout(t_12654));
compressor_4_2 u2_4449(.a(t_11894), .b(t_11891), .c(t_11889), .d(t_11886), .cin(t_12654), .o(t_12655), .co(t_12656), .cout(t_12657));
compressor_4_2 u2_4450(.a(t_11900), .b(t_11897), .c(t_11895), .d(t_11892), .cin(t_12657), .o(t_12658), .co(t_12659), .cout(t_12660));
compressor_4_2 u2_4451(.a(t_11906), .b(t_11903), .c(t_11901), .d(t_11898), .cin(t_12660), .o(t_12661), .co(t_12662), .cout(t_12663));
compressor_4_2 u2_4452(.a(t_11912), .b(t_11909), .c(t_11907), .d(t_11904), .cin(t_12663), .o(t_12664), .co(t_12665), .cout(t_12666));
compressor_4_2 u2_4453(.a(t_11918), .b(t_11915), .c(t_11913), .d(t_11910), .cin(t_12666), .o(t_12667), .co(t_12668), .cout(t_12669));
compressor_4_2 u2_4454(.a(t_11924), .b(t_11921), .c(t_11919), .d(t_11916), .cin(t_12669), .o(t_12670), .co(t_12671), .cout(t_12672));
compressor_4_2 u2_4455(.a(t_11930), .b(t_11927), .c(t_11925), .d(t_11922), .cin(t_12672), .o(t_12673), .co(t_12674), .cout(t_12675));
compressor_4_2 u2_4456(.a(t_11936), .b(t_11933), .c(t_11931), .d(t_11928), .cin(t_12675), .o(t_12676), .co(t_12677), .cout(t_12678));
compressor_4_2 u2_4457(.a(t_11942), .b(t_11939), .c(t_11937), .d(t_11934), .cin(t_12678), .o(t_12679), .co(t_12680), .cout(t_12681));
compressor_4_2 u2_4458(.a(t_11948), .b(t_11945), .c(t_11943), .d(t_11940), .cin(t_12681), .o(t_12682), .co(t_12683), .cout(t_12684));
compressor_4_2 u2_4459(.a(t_11954), .b(t_11951), .c(t_11949), .d(t_11946), .cin(t_12684), .o(t_12685), .co(t_12686), .cout(t_12687));
compressor_4_2 u2_4460(.a(t_11960), .b(t_11957), .c(t_11955), .d(t_11952), .cin(t_12687), .o(t_12688), .co(t_12689), .cout(t_12690));
compressor_4_2 u2_4461(.a(t_11966), .b(t_11963), .c(t_11961), .d(t_11958), .cin(t_12690), .o(t_12691), .co(t_12692), .cout(t_12693));
compressor_4_2 u2_4462(.a(t_11972), .b(t_11969), .c(t_11967), .d(t_11964), .cin(t_12693), .o(t_12694), .co(t_12695), .cout(t_12696));
compressor_4_2 u2_4463(.a(t_11978), .b(t_11975), .c(t_11973), .d(t_11970), .cin(t_12696), .o(t_12697), .co(t_12698), .cout(t_12699));
compressor_4_2 u2_4464(.a(t_11984), .b(t_11981), .c(t_11979), .d(t_11976), .cin(t_12699), .o(t_12700), .co(t_12701), .cout(t_12702));
compressor_4_2 u2_4465(.a(t_11990), .b(t_11987), .c(t_11985), .d(t_11982), .cin(t_12702), .o(t_12703), .co(t_12704), .cout(t_12705));
compressor_4_2 u2_4466(.a(t_11996), .b(t_11993), .c(t_11991), .d(t_11988), .cin(t_12705), .o(t_12706), .co(t_12707), .cout(t_12708));
compressor_4_2 u2_4467(.a(t_12002), .b(t_11999), .c(t_11997), .d(t_11994), .cin(t_12708), .o(t_12709), .co(t_12710), .cout(t_12711));
compressor_4_2 u2_4468(.a(t_12008), .b(t_12005), .c(t_12003), .d(t_12000), .cin(t_12711), .o(t_12712), .co(t_12713), .cout(t_12714));
compressor_4_2 u2_4469(.a(t_12014), .b(t_12011), .c(t_12009), .d(t_12006), .cin(t_12714), .o(t_12715), .co(t_12716), .cout(t_12717));
compressor_4_2 u2_4470(.a(t_12020), .b(t_12017), .c(t_12015), .d(t_12012), .cin(t_12717), .o(t_12718), .co(t_12719), .cout(t_12720));
compressor_4_2 u2_4471(.a(t_12026), .b(t_12023), .c(t_12021), .d(t_12018), .cin(t_12720), .o(t_12721), .co(t_12722), .cout(t_12723));
compressor_4_2 u2_4472(.a(t_12032), .b(t_12029), .c(t_12027), .d(t_12024), .cin(t_12723), .o(t_12724), .co(t_12725), .cout(t_12726));
compressor_4_2 u2_4473(.a(t_12035), .b(t_12033), .c(t_12030), .d(t_10854), .cin(t_12726), .o(t_12727), .co(t_12728), .cout(t_12729));
compressor_4_2 u2_4474(.a(t_12043), .b(t_12040), .c(t_12039), .d(t_12036), .cin(t_12729), .o(t_12730), .co(t_12731), .cout(t_12732));
compressor_4_2 u2_4475(.a(t_12048), .b(t_12045), .c(t_12044), .d(t_12041), .cin(t_12732), .o(t_12733), .co(t_12734), .cout(t_12735));
compressor_4_2 u2_4476(.a(t_12053), .b(t_12050), .c(t_12049), .d(t_12046), .cin(t_12735), .o(t_12736), .co(t_12737), .cout(t_12738));
compressor_4_2 u2_4477(.a(t_12058), .b(t_12055), .c(t_12054), .d(t_12051), .cin(t_12738), .o(t_12739), .co(t_12740), .cout(t_12741));
compressor_4_2 u2_4478(.a(t_12063), .b(t_12060), .c(t_12059), .d(t_12056), .cin(t_12741), .o(t_12742), .co(t_12743), .cout(t_12744));
compressor_4_2 u2_4479(.a(t_12068), .b(t_12065), .c(t_12064), .d(t_12061), .cin(t_12744), .o(t_12745), .co(t_12746), .cout(t_12747));
compressor_4_2 u2_4480(.a(t_12073), .b(t_12070), .c(t_12069), .d(t_12066), .cin(t_12747), .o(t_12748), .co(t_12749), .cout(t_12750));
compressor_4_2 u2_4481(.a(t_12078), .b(t_12075), .c(t_12074), .d(t_12071), .cin(t_12750), .o(t_12751), .co(t_12752), .cout(t_12753));
compressor_4_2 u2_4482(.a(t_12083), .b(t_12080), .c(t_12079), .d(t_12076), .cin(t_12753), .o(t_12754), .co(t_12755), .cout(t_12756));
compressor_4_2 u2_4483(.a(t_12088), .b(t_12085), .c(t_12084), .d(t_12081), .cin(t_12756), .o(t_12757), .co(t_12758), .cout(t_12759));
compressor_4_2 u2_4484(.a(t_12093), .b(t_12090), .c(t_12089), .d(t_12086), .cin(t_12759), .o(t_12760), .co(t_12761), .cout(t_12762));
compressor_4_2 u2_4485(.a(t_12098), .b(t_12095), .c(t_12094), .d(t_12091), .cin(t_12762), .o(t_12763), .co(t_12764), .cout(t_12765));
compressor_4_2 u2_4486(.a(t_12103), .b(t_12100), .c(t_12099), .d(t_12096), .cin(t_12765), .o(t_12766), .co(t_12767), .cout(t_12768));
compressor_4_2 u2_4487(.a(t_12108), .b(t_12105), .c(t_12104), .d(t_12101), .cin(t_12768), .o(t_12769), .co(t_12770), .cout(t_12771));
compressor_4_2 u2_4488(.a(t_12113), .b(t_12110), .c(t_12109), .d(t_12106), .cin(t_12771), .o(t_12772), .co(t_12773), .cout(t_12774));
compressor_4_2 u2_4489(.a(t_12118), .b(t_12115), .c(t_12114), .d(t_12111), .cin(t_12774), .o(t_12775), .co(t_12776), .cout(t_12777));
compressor_4_2 u2_4490(.a(t_12123), .b(t_12120), .c(t_12119), .d(t_12116), .cin(t_12777), .o(t_12778), .co(t_12779), .cout(t_12780));
compressor_4_2 u2_4491(.a(t_12128), .b(t_12125), .c(t_12124), .d(t_12121), .cin(t_12780), .o(t_12781), .co(t_12782), .cout(t_12783));
compressor_4_2 u2_4492(.a(t_12133), .b(t_12130), .c(t_12129), .d(t_12126), .cin(t_12783), .o(t_12784), .co(t_12785), .cout(t_12786));
compressor_4_2 u2_4493(.a(t_12138), .b(t_12135), .c(t_12134), .d(t_12131), .cin(t_12786), .o(t_12787), .co(t_12788), .cout(t_12789));
compressor_4_2 u2_4494(.a(t_12143), .b(t_12140), .c(t_12139), .d(t_12136), .cin(t_12789), .o(t_12790), .co(t_12791), .cout(t_12792));
compressor_4_2 u2_4495(.a(t_12148), .b(t_12145), .c(t_12144), .d(t_12141), .cin(t_12792), .o(t_12793), .co(t_12794), .cout(t_12795));
compressor_4_2 u2_4496(.a(t_12153), .b(t_12150), .c(t_12149), .d(t_12146), .cin(t_12795), .o(t_12796), .co(t_12797), .cout(t_12798));
compressor_4_2 u2_4497(.a(t_12158), .b(t_12155), .c(t_12154), .d(t_12151), .cin(t_12798), .o(t_12799), .co(t_12800), .cout(t_12801));
compressor_4_2 u2_4498(.a(t_12163), .b(t_12160), .c(t_12159), .d(t_12156), .cin(t_12801), .o(t_12802), .co(t_12803), .cout(t_12804));
compressor_4_2 u2_4499(.a(t_12168), .b(t_12165), .c(t_12164), .d(t_12161), .cin(t_12804), .o(t_12805), .co(t_12806), .cout(t_12807));
compressor_4_2 u2_4500(.a(t_12173), .b(t_12170), .c(t_12169), .d(t_12166), .cin(t_12807), .o(t_12808), .co(t_12809), .cout(t_12810));
compressor_4_2 u2_4501(.a(t_12178), .b(t_12175), .c(t_12174), .d(t_12171), .cin(t_12810), .o(t_12811), .co(t_12812), .cout(t_12813));
compressor_4_2 u2_4502(.a(t_12183), .b(t_12180), .c(t_12179), .d(t_12176), .cin(t_12813), .o(t_12814), .co(t_12815), .cout(t_12816));
compressor_4_2 u2_4503(.a(t_12188), .b(t_12185), .c(t_12184), .d(t_12181), .cin(t_12816), .o(t_12817), .co(t_12818), .cout(t_12819));
compressor_4_2 u2_4504(.a(t_12193), .b(t_12190), .c(t_12189), .d(t_12186), .cin(t_12819), .o(t_12820), .co(t_12821), .cout(t_12822));
compressor_4_2 u2_4505(.a(t_12195), .b(t_12194), .c(t_12191), .d(t_11123), .cin(t_12822), .o(t_12823), .co(t_12824), .cout(t_12825));
compressor_3_2 u1_4506(.a(t_12198), .b(t_12196), .cin(t_12825), .o(t_12826), .cout(t_12827));
compressor_3_2 u1_4507(.a(t_12201), .b(t_12199), .cin(t_11135), .o(t_12828), .cout(t_12829));
half_adder u0_4508(.a(t_12204), .b(t_12202), .o(t_12830), .cout(t_12831));
half_adder u0_4509(.a(t_12207), .b(t_12205), .o(t_12832), .cout(t_12833));
half_adder u0_4510(.a(t_12210), .b(t_12208), .o(t_12834), .cout(t_12835));
half_adder u0_4511(.a(t_12213), .b(t_12211), .o(t_12836), .cout(t_12837));
compressor_3_2 u1_4512(.a(t_12216), .b(t_12214), .cin(t_11165), .o(t_12838), .cout(t_12839));
half_adder u0_4513(.a(t_12219), .b(t_12217), .o(t_12840), .cout(t_12841));
half_adder u0_4514(.a(t_12222), .b(t_12220), .o(t_12842), .cout(t_12843));
half_adder u0_4515(.a(t_12225), .b(t_12223), .o(t_12844), .cout(t_12845));
half_adder u0_4516(.a(t_12228), .b(t_12226), .o(t_12846), .cout(t_12847));
half_adder u0_4517(.a(t_12231), .b(t_12229), .o(t_12848), .cout(t_12849));
half_adder u0_4518(.a(t_12234), .b(t_12232), .o(t_12850), .cout(t_12851));
half_adder u0_4519(.a(t_12237), .b(t_12235), .o(t_12852), .cout(t_12853));
half_adder u0_4520(.a(t_12240), .b(t_12238), .o(t_12854), .cout(t_12855));
half_adder u0_4521(.a(t_12243), .b(t_12241), .o(t_12856), .cout(t_12857));
half_adder u0_4522(.a(t_12246), .b(t_12244), .o(t_12858), .cout(t_12859));
half_adder u0_4523(.a(t_12249), .b(t_12247), .o(t_12860), .cout(t_12861));
half_adder u0_4524(.a(t_12252), .b(t_12250), .o(t_12862), .cout(t_12863));
half_adder u0_4525(.a(t_12255), .b(t_12253), .o(t_12864), .cout(t_12865));
half_adder u0_4526(.a(t_12258), .b(t_12256), .o(t_12866), .cout(t_12867));
half_adder u0_4527(.a(t_12261), .b(t_12259), .o(t_12868), .cout(t_12869));
half_adder u0_4528(.a(t_12264), .b(t_12262), .o(t_12870), .cout(t_12871));
half_adder u0_4529(.a(t_12267), .b(t_12265), .o(t_12872), .cout(t_12873));
half_adder u0_4530(.a(t_12270), .b(t_12268), .o(t_12874), .cout(t_12875));
half_adder u0_4531(.a(t_12273), .b(t_12271), .o(t_12876), .cout(t_12877));
half_adder u0_4532(.a(t_12276), .b(t_12274), .o(t_12878), .cout(t_12879));
half_adder u0_4533(.a(t_12279), .b(t_12277), .o(t_12880), .cout(t_12881));
half_adder u0_4534(.a(t_12282), .b(t_12280), .o(t_12882), .cout(t_12883));
half_adder u0_4535(.a(t_12285), .b(t_12283), .o(t_12884), .cout(t_12885));
half_adder u0_4536(.a(t_12288), .b(t_12286), .o(t_12886), .cout(t_12887));
compressor_3_2 u1_4537(.a(t_12291), .b(t_12289), .cin(t_11296), .o(t_12888), .cout(t_12889));
half_adder u0_4538(.a(t_12293), .b(t_12292), .o(t_12890), .cout(t_12891));
half_adder u0_4539(.a(t_12295), .b(t_12294), .o(t_12892), .cout(t_12893));
half_adder u0_4540(.a(t_12297), .b(t_12296), .o(t_12894), .cout(t_12895));
half_adder u0_4541(.a(t_12299), .b(t_12298), .o(t_12896), .cout(t_12897));
half_adder u0_4542(.a(t_12301), .b(t_12300), .o(t_12898), .cout(t_12899));
half_adder u0_4543(.a(t_12303), .b(t_12302), .o(t_12900), .cout(t_12901));
half_adder u0_4544(.a(t_12305), .b(t_12304), .o(t_12902), .cout(t_12903));
half_adder u0_4545(.a(t_12307), .b(t_12306), .o(t_12904), .cout(t_12905));
half_adder u0_4546(.a(t_12309), .b(t_12308), .o(t_12906), .cout(t_12907));
half_adder u0_4547(.a(t_12311), .b(t_12310), .o(t_12908), .cout(t_12909));
half_adder u0_4548(.a(t_12313), .b(t_12312), .o(t_12910), .cout(t_12911));
half_adder u0_4549(.a(t_12315), .b(t_12314), .o(t_12912), .cout(t_12913));
half_adder u0_4550(.a(t_12317), .b(t_12316), .o(t_12914), .cout(t_12915));
half_adder u0_4551(.a(t_12319), .b(t_12318), .o(t_12916), .cout(t_12917));
half_adder u0_4552(.a(t_12321), .b(t_12320), .o(t_12918), .cout(t_12919));
half_adder u0_4553(.a(t_12323), .b(t_12322), .o(t_12920), .cout(t_12921));
half_adder u0_4554(.a(t_12325), .b(t_12324), .o(t_12922), .cout(t_12923));
half_adder u0_4555(.a(t_12327), .b(t_12326), .o(t_12924), .cout(t_12925));
half_adder u0_4556(.a(t_12329), .b(t_12328), .o(t_12926), .cout(t_12927));
half_adder u0_4557(.a(t_12331), .b(t_12330), .o(t_12928), .cout(t_12929));
half_adder u0_4558(.a(t_12333), .b(t_12332), .o(t_12930), .cout(t_12931));
half_adder u0_4559(.a(t_12335), .b(t_12334), .o(t_12932), .cout(t_12933));
half_adder u0_4560(.a(t_12337), .b(t_12336), .o(t_12934), .cout(t_12935));
half_adder u0_4561(.a(t_12339), .b(t_12338), .o(t_12936), .cout(t_12937));
half_adder u0_4562(.a(t_12341), .b(t_12340), .o(t_12938), .cout(t_12939));
half_adder u0_4563(.a(t_12343), .b(t_12342), .o(t_12940), .cout(t_12941));
half_adder u0_4564(.a(t_12345), .b(t_12344), .o(t_12942), .cout(t_12943));
half_adder u0_4565(.a(t_12347), .b(t_12346), .o(t_12944), .cout(t_12945));
half_adder u0_4566(.a(t_12349), .b(t_12348), .o(t_12946), .cout());

/* u0_4567 Output nets */
wire t_12947,  t_12948;
/* u0_4568 Output nets */
wire t_12949,  t_12950;
/* u0_4569 Output nets */
wire t_12951,  t_12952;
/* u0_4570 Output nets */
wire t_12953,  t_12954;
/* u0_4571 Output nets */
wire t_12955,  t_12956;
/* u0_4572 Output nets */
wire t_12957,  t_12958;
/* u0_4573 Output nets */
wire t_12959,  t_12960;
/* u0_4574 Output nets */
wire t_12961,  t_12962;
/* u0_4575 Output nets */
wire t_12963,  t_12964;
/* u0_4576 Output nets */
wire t_12965,  t_12966;
/* u0_4577 Output nets */
wire t_12967,  t_12968;
/* u0_4578 Output nets */
wire t_12969,  t_12970;
/* u0_4579 Output nets */
wire t_12971,  t_12972;
/* u0_4580 Output nets */
wire t_12973,  t_12974;
/* u0_4581 Output nets */
wire t_12975,  t_12976;
/* u0_4582 Output nets */
wire t_12977,  t_12978;
/* u0_4583 Output nets */
wire t_12979,  t_12980;
/* u0_4584 Output nets */
wire t_12981,  t_12982;
/* u0_4585 Output nets */
wire t_12983,  t_12984;
/* u0_4586 Output nets */
wire t_12985,  t_12986;
/* u0_4587 Output nets */
wire t_12987,  t_12988;
/* u0_4588 Output nets */
wire t_12989,  t_12990;
/* u0_4589 Output nets */
wire t_12991,  t_12992;
/* u0_4590 Output nets */
wire t_12993,  t_12994;
/* u0_4591 Output nets */
wire t_12995,  t_12996;
/* u0_4592 Output nets */
wire t_12997,  t_12998;
/* u0_4593 Output nets */
wire t_12999,  t_13000;
/* u0_4594 Output nets */
wire t_13001,  t_13002;
/* u0_4595 Output nets */
wire t_13003,  t_13004;
/* u0_4596 Output nets */
wire t_13005,  t_13006;
/* u0_4597 Output nets */
wire t_13007,  t_13008;
/* u0_4598 Output nets */
wire t_13009,  t_13010;
/* u0_4599 Output nets */
wire t_13011,  t_13012;
/* u0_4600 Output nets */
wire t_13013,  t_13014;
/* u0_4601 Output nets */
wire t_13015,  t_13016;
/* u0_4602 Output nets */
wire t_13017,  t_13018;
/* u0_4603 Output nets */
wire t_13019,  t_13020;
/* u0_4604 Output nets */
wire t_13021,  t_13022;
/* u0_4605 Output nets */
wire t_13023,  t_13024;
/* u0_4606 Output nets */
wire t_13025,  t_13026;
/* u0_4607 Output nets */
wire t_13027,  t_13028;
/* u0_4608 Output nets */
wire t_13029,  t_13030;
/* u0_4609 Output nets */
wire t_13031,  t_13032;
/* u0_4610 Output nets */
wire t_13033,  t_13034;
/* u0_4611 Output nets */
wire t_13035,  t_13036;
/* u0_4612 Output nets */
wire t_13037,  t_13038;
/* u0_4613 Output nets */
wire t_13039,  t_13040;
/* u0_4614 Output nets */
wire t_13041,  t_13042;
/* u0_4615 Output nets */
wire t_13043,  t_13044;
/* u0_4616 Output nets */
wire t_13045,  t_13046;
/* u0_4617 Output nets */
wire t_13047,  t_13048;
/* u0_4618 Output nets */
wire t_13049,  t_13050;
/* u0_4619 Output nets */
wire t_13051,  t_13052;
/* u0_4620 Output nets */
wire t_13053,  t_13054;
/* u0_4621 Output nets */
wire t_13055,  t_13056;
/* u0_4622 Output nets */
wire t_13057,  t_13058;
/* u0_4623 Output nets */
wire t_13059,  t_13060;
/* u0_4624 Output nets */
wire t_13061,  t_13062;
/* u0_4625 Output nets */
wire t_13063,  t_13064;
/* u0_4626 Output nets */
wire t_13065,  t_13066;
/* u0_4627 Output nets */
wire t_13067,  t_13068;
/* u0_4628 Output nets */
wire t_13069,  t_13070;
/* u1_4629 Output nets */
wire t_13071,  t_13072;
/* u0_4630 Output nets */
wire t_13073,  t_13074;
/* u1_4631 Output nets */
wire t_13075,  t_13076;
/* u1_4632 Output nets */
wire t_13077,  t_13078;
/* u1_4633 Output nets */
wire t_13079,  t_13080;
/* u1_4634 Output nets */
wire t_13081,  t_13082;
/* u1_4635 Output nets */
wire t_13083,  t_13084;
/* u1_4636 Output nets */
wire t_13085,  t_13086;
/* u1_4637 Output nets */
wire t_13087,  t_13088;
/* u1_4638 Output nets */
wire t_13089,  t_13090;
/* u1_4639 Output nets */
wire t_13091,  t_13092;
/* u1_4640 Output nets */
wire t_13093,  t_13094;
/* u1_4641 Output nets */
wire t_13095,  t_13096;
/* u1_4642 Output nets */
wire t_13097,  t_13098;
/* u1_4643 Output nets */
wire t_13099,  t_13100;
/* u1_4644 Output nets */
wire t_13101,  t_13102;
/* u1_4645 Output nets */
wire t_13103,  t_13104;
/* u1_4646 Output nets */
wire t_13105,  t_13106;
/* u1_4647 Output nets */
wire t_13107,  t_13108;
/* u1_4648 Output nets */
wire t_13109,  t_13110;
/* u1_4649 Output nets */
wire t_13111,  t_13112;
/* u1_4650 Output nets */
wire t_13113,  t_13114;
/* u1_4651 Output nets */
wire t_13115,  t_13116;
/* u1_4652 Output nets */
wire t_13117,  t_13118;
/* u1_4653 Output nets */
wire t_13119,  t_13120;
/* u1_4654 Output nets */
wire t_13121,  t_13122;
/* u1_4655 Output nets */
wire t_13123,  t_13124;
/* u1_4656 Output nets */
wire t_13125,  t_13126;
/* u1_4657 Output nets */
wire t_13127,  t_13128;
/* u1_4658 Output nets */
wire t_13129,  t_13130;
/* u1_4659 Output nets */
wire t_13131,  t_13132;
/* u0_4660 Output nets */
wire t_13133,  t_13134;
/* u0_4661 Output nets */
wire t_13135,  t_13136;
/* u1_4662 Output nets */
wire t_13137,  t_13138;
/* u1_4663 Output nets */
wire t_13139,  t_13140;
/* u1_4664 Output nets */
wire t_13141,  t_13142;
/* u1_4665 Output nets */
wire t_13143,  t_13144;
/* u1_4666 Output nets */
wire t_13145,  t_13146;
/* u1_4667 Output nets */
wire t_13147,  t_13148;
/* u1_4668 Output nets */
wire t_13149,  t_13150;
/* u1_4669 Output nets */
wire t_13151,  t_13152;
/* u1_4670 Output nets */
wire t_13153,  t_13154;
/* u1_4671 Output nets */
wire t_13155,  t_13156;
/* u1_4672 Output nets */
wire t_13157,  t_13158;
/* u1_4673 Output nets */
wire t_13159,  t_13160;
/* u1_4674 Output nets */
wire t_13161,  t_13162;
/* u0_4675 Output nets */
wire t_13163,  t_13164;
/* u0_4676 Output nets */
wire t_13165,  t_13166;
/* u1_4677 Output nets */
wire t_13167,  t_13168;
/* u1_4678 Output nets */
wire t_13169,  t_13170;
/* u1_4679 Output nets */
wire t_13171,  t_13172;
/* u1_4680 Output nets */
wire t_13173,  t_13174;
/* u1_4681 Output nets */
wire t_13175,  t_13176;
/* u0_4682 Output nets */
wire t_13177,  t_13178;
/* u0_4683 Output nets */
wire t_13179,  t_13180;
/* u1_4684 Output nets */
wire t_13181,  t_13182;
/* u0_4685 Output nets */
wire t_13183,  t_13184;
/* u0_4686 Output nets */
wire t_13185,  t_13186;
/* u0_4687 Output nets */
wire t_13187,  t_13188;
/* u0_4688 Output nets */
wire t_13189,  t_13190;
/* u1_4689 Output nets */
wire t_13191,  t_13192;
/* u1_4690 Output nets */
wire t_13193,  t_13194;
/* u0_4691 Output nets */
wire t_13195,  t_13196;
/* u0_4692 Output nets */
wire t_13197,  t_13198;
/* u1_4693 Output nets */
wire t_13199,  t_13200;
/* u0_4694 Output nets */
wire t_13201,  t_13202;
/* u0_4695 Output nets */
wire t_13203,  t_13204;
/* u0_4696 Output nets */
wire t_13205,  t_13206;
/* u0_4697 Output nets */
wire t_13207,  t_13208;
/* u1_4698 Output nets */
wire t_13209,  t_13210;
/* u0_4699 Output nets */
wire t_13211,  t_13212;
/* u0_4700 Output nets */
wire t_13213,  t_13214;
/* u0_4701 Output nets */
wire t_13215,  t_13216;
/* u0_4702 Output nets */
wire t_13217,  t_13218;
/* u0_4703 Output nets */
wire t_13219,  t_13220;
/* u0_4704 Output nets */
wire t_13221,  t_13222;
/* u0_4705 Output nets */
wire t_13223,  t_13224;
/* u0_4706 Output nets */
wire t_13225,  t_13226;
/* u0_4707 Output nets */
wire t_13227,  t_13228;
/* u0_4708 Output nets */
wire t_13229,  t_13230;
/* u0_4709 Output nets */
wire t_13231,  t_13232;
/* u0_4710 Output nets */
wire t_13233,  t_13234;
/* u0_4711 Output nets */
wire t_13235,  t_13236;
/* u0_4712 Output nets */
wire t_13237,  t_13238;
/* u0_4713 Output nets */
wire t_13239,  t_13240;
/* u0_4714 Output nets */
wire t_13241,  t_13242;
/* u0_4715 Output nets */
wire t_13243,  t_13244;
/* u0_4716 Output nets */
wire t_13245,  t_13246;
/* u0_4717 Output nets */
wire t_13247,  t_13248;
/* u0_4718 Output nets */
wire t_13249,  t_13250;
/* u0_4719 Output nets */
wire t_13251,  t_13252;
/* u0_4720 Output nets */
wire t_13253,  t_13254;
/* u0_4721 Output nets */
wire t_13255,  t_13256;
/* u0_4722 Output nets */
wire t_13257,  t_13258;
/* u1_4723 Output nets */
wire t_13259,  t_13260;
/* u0_4724 Output nets */
wire t_13261,  t_13262;
/* u0_4725 Output nets */
wire t_13263,  t_13264;
/* u0_4726 Output nets */
wire t_13265,  t_13266;
/* u0_4727 Output nets */
wire t_13267,  t_13268;
/* u0_4728 Output nets */
wire t_13269,  t_13270;
/* u0_4729 Output nets */
wire t_13271,  t_13272;
/* u0_4730 Output nets */
wire t_13273,  t_13274;
/* u0_4731 Output nets */
wire t_13275,  t_13276;
/* u0_4732 Output nets */
wire t_13277,  t_13278;
/* u0_4733 Output nets */
wire t_13279,  t_13280;
/* u0_4734 Output nets */
wire t_13281,  t_13282;
/* u0_4735 Output nets */
wire t_13283,  t_13284;
/* u0_4736 Output nets */
wire t_13285,  t_13286;
/* u0_4737 Output nets */
wire t_13287,  t_13288;
/* u0_4738 Output nets */
wire t_13289,  t_13290;
/* u0_4739 Output nets */
wire t_13291,  t_13292;
/* u0_4740 Output nets */
wire t_13293,  t_13294;
/* u0_4741 Output nets */
wire t_13295,  t_13296;
/* u0_4742 Output nets */
wire t_13297,  t_13298;
/* u0_4743 Output nets */
wire t_13299,  t_13300;
/* u0_4744 Output nets */
wire t_13301,  t_13302;
/* u0_4745 Output nets */
wire t_13303,  t_13304;
/* u0_4746 Output nets */
wire t_13305,  t_13306;
/* u0_4747 Output nets */
wire t_13307,  t_13308;
/* u0_4748 Output nets */
wire t_13309,  t_13310;
/* u0_4749 Output nets */
wire t_13311,  t_13312;
/* u0_4750 Output nets */
wire t_13313,  t_13314;
/* u0_4751 Output nets */
wire t_13315,  t_13316;
/* u0_4752 Output nets */
wire t_13317,  t_13318;
/* u0_4753 Output nets */
wire t_13319,  t_13320;
/* u0_4754 Output nets */
wire t_13321,  t_13322;
/* u0_4755 Output nets */
wire t_13323,  t_13324;
/* u0_4756 Output nets */
wire t_13325,  t_13326;
/* u0_4757 Output nets */
wire t_13327,  t_13328;
/* u0_4758 Output nets */
wire t_13329,  t_13330;
/* u0_4759 Output nets */
wire t_13331,  t_13332;
/* u0_4760 Output nets */
wire t_13333,  t_13334;
/* u0_4761 Output nets */
wire t_13335,  t_13336;
/* u0_4762 Output nets */
wire t_13337,  t_13338;
/* u0_4763 Output nets */
wire t_13339,  t_13340;
/* u0_4764 Output nets */
wire t_13341,  t_13342;
/* u0_4765 Output nets */
wire t_13343,  t_13344;
/* u0_4766 Output nets */
wire t_13345,  t_13346;
/* u0_4767 Output nets */
wire t_13347,  t_13348;
/* u0_4768 Output nets */
wire t_13349,  t_13350;
/* u0_4769 Output nets */
wire t_13351,  t_13352;
/* u0_4770 Output nets */
wire t_13353,  t_13354;
/* u0_4771 Output nets */
wire t_13355,  t_13356;
/* u0_4772 Output nets */
wire t_13357,  t_13358;
/* u0_4773 Output nets */
wire t_13359,  t_13360;
/* u0_4774 Output nets */
wire t_13361,  t_13362;
/* u0_4775 Output nets */
wire t_13363,  t_13364;
/* u0_4776 Output nets */
wire t_13365,  t_13366;
/* u0_4777 Output nets */
wire t_13367,  t_13368;
/* u0_4778 Output nets */
wire t_13369,  t_13370;
/* u0_4779 Output nets */
wire t_13371,  t_13372;
/* u0_4780 Output nets */
wire t_13373,  t_13374;
/* u0_4781 Output nets */
wire t_13375,  t_13376;
/* u0_4782 Output nets */
wire t_13377,  t_13378;
/* u0_4783 Output nets */
wire t_13379,  t_13380;
/* u0_4784 Output nets */
wire t_13381,  t_13382;
/* u0_4785 Output nets */
wire t_13383,  t_13384;
/* u0_4786 Output nets */
wire t_13385,  t_13386;
/* u0_4787 Output nets */
wire t_13387,  t_13388;
/* u0_4788 Output nets */
wire t_13389,  t_13390;
/* u0_4789 Output nets */
wire t_13391,  t_13392;
/* u0_4790 Output nets */
wire t_13393,  t_13394;
/* u0_4791 Output nets */
wire t_13395,  t_13396;
/* u0_4792 Output nets */
wire t_13397,  t_13398;
/* u0_4793 Output nets */
wire t_13399,  t_13400;
/* u0_4794 Output nets */
wire t_13401,  t_13402;
/* u0_4795 Output nets */
wire t_13403,  t_13404;
/* u0_4796 Output nets */
wire t_13405,  t_13406;
/* u0_4797 Output nets */
wire t_13407,  t_13408;
/* u0_4798 Output nets */
wire t_13409,  t_13410;
/* u0_4799 Output nets */
wire t_13411,  t_13412;
/* u0_4800 Output nets */
wire t_13413,  t_13414;
/* u0_4801 Output nets */
wire t_13415,  t_13416;
/* u0_4802 Output nets */
wire t_13417,  t_13418;
/* u0_4803 Output nets */
wire t_13419,  t_13420;
/* u0_4804 Output nets */
wire t_13421,  t_13422;
/* u0_4805 Output nets */
wire t_13423,  t_13424;
/* u0_4806 Output nets */
wire t_13425,  t_13426;
/* u0_4807 Output nets */
wire t_13427,  t_13428;
/* u0_4808 Output nets */
wire t_13429,  t_13430;
/* u0_4809 Output nets */
wire t_13431,  t_13432;
/* u0_4810 Output nets */
wire t_13433,  t_13434;
/* u0_4811 Output nets */
wire t_13435,  t_13436;
/* u0_4812 Output nets */
wire t_13437,  t_13438;
/* u0_4813 Output nets */
wire t_13439,  t_13440;
/* u0_4814 Output nets */
wire t_13441,  t_13442;
/* u0_4815 Output nets */
wire t_13443,  t_13444;
/* u0_4816 Output nets */
wire t_13445;

/* compress stage 6 */
half_adder u0_4567(.a(t_12351), .b(t_11373), .o(t_12947), .cout(t_12948));
half_adder u0_4568(.a(t_12354), .b(t_12353), .o(t_12949), .cout(t_12950));
half_adder u0_4569(.a(t_12356), .b(t_12355), .o(t_12951), .cout(t_12952));
half_adder u0_4570(.a(t_12358), .b(t_12357), .o(t_12953), .cout(t_12954));
half_adder u0_4571(.a(t_12360), .b(t_12359), .o(t_12955), .cout(t_12956));
half_adder u0_4572(.a(t_12362), .b(t_12361), .o(t_12957), .cout(t_12958));
half_adder u0_4573(.a(t_12364), .b(t_12363), .o(t_12959), .cout(t_12960));
half_adder u0_4574(.a(t_12366), .b(t_12365), .o(t_12961), .cout(t_12962));
half_adder u0_4575(.a(t_12368), .b(t_12367), .o(t_12963), .cout(t_12964));
half_adder u0_4576(.a(t_12370), .b(t_12369), .o(t_12965), .cout(t_12966));
half_adder u0_4577(.a(t_12372), .b(t_12371), .o(t_12967), .cout(t_12968));
half_adder u0_4578(.a(t_12374), .b(t_12373), .o(t_12969), .cout(t_12970));
half_adder u0_4579(.a(t_12376), .b(t_12375), .o(t_12971), .cout(t_12972));
half_adder u0_4580(.a(t_12378), .b(t_12377), .o(t_12973), .cout(t_12974));
half_adder u0_4581(.a(t_12380), .b(t_12379), .o(t_12975), .cout(t_12976));
half_adder u0_4582(.a(t_12382), .b(t_12381), .o(t_12977), .cout(t_12978));
half_adder u0_4583(.a(t_12384), .b(t_12383), .o(t_12979), .cout(t_12980));
half_adder u0_4584(.a(t_12386), .b(t_12385), .o(t_12981), .cout(t_12982));
half_adder u0_4585(.a(t_12388), .b(t_12387), .o(t_12983), .cout(t_12984));
half_adder u0_4586(.a(t_12390), .b(t_12389), .o(t_12985), .cout(t_12986));
half_adder u0_4587(.a(t_12392), .b(t_12391), .o(t_12987), .cout(t_12988));
half_adder u0_4588(.a(t_12394), .b(t_12393), .o(t_12989), .cout(t_12990));
half_adder u0_4589(.a(t_12396), .b(t_12395), .o(t_12991), .cout(t_12992));
half_adder u0_4590(.a(t_12398), .b(t_12397), .o(t_12993), .cout(t_12994));
half_adder u0_4591(.a(t_12400), .b(t_12399), .o(t_12995), .cout(t_12996));
half_adder u0_4592(.a(t_12402), .b(t_12401), .o(t_12997), .cout(t_12998));
half_adder u0_4593(.a(t_12404), .b(t_12403), .o(t_12999), .cout(t_13000));
half_adder u0_4594(.a(t_12406), .b(t_12405), .o(t_13001), .cout(t_13002));
half_adder u0_4595(.a(t_12408), .b(t_12407), .o(t_13003), .cout(t_13004));
half_adder u0_4596(.a(t_12410), .b(t_12409), .o(t_13005), .cout(t_13006));
half_adder u0_4597(.a(t_12412), .b(t_12411), .o(t_13007), .cout(t_13008));
half_adder u0_4598(.a(t_12414), .b(t_12413), .o(t_13009), .cout(t_13010));
half_adder u0_4599(.a(t_12416), .b(t_12415), .o(t_13011), .cout(t_13012));
half_adder u0_4600(.a(t_12418), .b(t_12417), .o(t_13013), .cout(t_13014));
half_adder u0_4601(.a(t_12420), .b(t_12419), .o(t_13015), .cout(t_13016));
half_adder u0_4602(.a(t_12422), .b(t_12421), .o(t_13017), .cout(t_13018));
half_adder u0_4603(.a(t_12424), .b(t_12423), .o(t_13019), .cout(t_13020));
half_adder u0_4604(.a(t_12426), .b(t_12425), .o(t_13021), .cout(t_13022));
half_adder u0_4605(.a(t_12428), .b(t_12427), .o(t_13023), .cout(t_13024));
half_adder u0_4606(.a(t_12430), .b(t_12429), .o(t_13025), .cout(t_13026));
half_adder u0_4607(.a(t_12432), .b(t_12431), .o(t_13027), .cout(t_13028));
half_adder u0_4608(.a(t_12434), .b(t_12433), .o(t_13029), .cout(t_13030));
half_adder u0_4609(.a(t_12436), .b(t_12435), .o(t_13031), .cout(t_13032));
half_adder u0_4610(.a(t_12438), .b(t_12437), .o(t_13033), .cout(t_13034));
half_adder u0_4611(.a(t_12440), .b(t_12439), .o(t_13035), .cout(t_13036));
half_adder u0_4612(.a(t_12442), .b(t_12441), .o(t_13037), .cout(t_13038));
half_adder u0_4613(.a(t_12444), .b(t_12443), .o(t_13039), .cout(t_13040));
half_adder u0_4614(.a(t_12446), .b(t_12445), .o(t_13041), .cout(t_13042));
half_adder u0_4615(.a(t_12448), .b(t_12447), .o(t_13043), .cout(t_13044));
half_adder u0_4616(.a(t_12450), .b(t_12449), .o(t_13045), .cout(t_13046));
half_adder u0_4617(.a(t_12452), .b(t_12451), .o(t_13047), .cout(t_13048));
half_adder u0_4618(.a(t_12454), .b(t_12453), .o(t_13049), .cout(t_13050));
half_adder u0_4619(.a(t_12456), .b(t_12455), .o(t_13051), .cout(t_13052));
half_adder u0_4620(.a(t_12458), .b(t_12457), .o(t_13053), .cout(t_13054));
half_adder u0_4621(.a(t_12460), .b(t_12459), .o(t_13055), .cout(t_13056));
half_adder u0_4622(.a(t_12462), .b(t_12461), .o(t_13057), .cout(t_13058));
half_adder u0_4623(.a(t_12464), .b(t_12463), .o(t_13059), .cout(t_13060));
half_adder u0_4624(.a(t_12466), .b(t_12465), .o(t_13061), .cout(t_13062));
half_adder u0_4625(.a(t_12468), .b(t_12467), .o(t_13063), .cout(t_13064));
half_adder u0_4626(.a(t_12470), .b(t_12469), .o(t_13065), .cout(t_13066));
half_adder u0_4627(.a(t_12472), .b(t_12471), .o(t_13067), .cout(t_13068));
half_adder u0_4628(.a(t_12474), .b(t_12473), .o(t_13069), .cout(t_13070));
compressor_3_2 u1_4629(.a(t_12476), .b(t_12475), .cin(t_11519), .o(t_13071), .cout(t_13072));
half_adder u0_4630(.a(t_12478), .b(t_12477), .o(t_13073), .cout(t_13074));
compressor_3_2 u1_4631(.a(t_12480), .b(t_12479), .cin(t_11530), .o(t_13075), .cout(t_13076));
compressor_3_2 u1_4632(.a(t_12482), .b(t_12481), .cin(t_11535), .o(t_13077), .cout(t_13078));
compressor_3_2 u1_4633(.a(t_12484), .b(t_12483), .cin(t_11540), .o(t_13079), .cout(t_13080));
compressor_3_2 u1_4634(.a(t_12486), .b(t_12485), .cin(t_11545), .o(t_13081), .cout(t_13082));
compressor_3_2 u1_4635(.a(t_12488), .b(t_12487), .cin(t_11550), .o(t_13083), .cout(t_13084));
compressor_3_2 u1_4636(.a(t_12490), .b(t_12489), .cin(t_11555), .o(t_13085), .cout(t_13086));
compressor_3_2 u1_4637(.a(t_12492), .b(t_12491), .cin(t_11560), .o(t_13087), .cout(t_13088));
compressor_3_2 u1_4638(.a(t_12494), .b(t_12493), .cin(t_11565), .o(t_13089), .cout(t_13090));
compressor_3_2 u1_4639(.a(t_12496), .b(t_12495), .cin(t_11570), .o(t_13091), .cout(t_13092));
compressor_3_2 u1_4640(.a(t_12498), .b(t_12497), .cin(t_11575), .o(t_13093), .cout(t_13094));
compressor_3_2 u1_4641(.a(t_12500), .b(t_12499), .cin(t_11580), .o(t_13095), .cout(t_13096));
compressor_3_2 u1_4642(.a(t_12502), .b(t_12501), .cin(t_11585), .o(t_13097), .cout(t_13098));
compressor_3_2 u1_4643(.a(t_12504), .b(t_12503), .cin(t_11590), .o(t_13099), .cout(t_13100));
compressor_3_2 u1_4644(.a(t_12506), .b(t_12505), .cin(t_11595), .o(t_13101), .cout(t_13102));
compressor_3_2 u1_4645(.a(t_12508), .b(t_12507), .cin(t_11600), .o(t_13103), .cout(t_13104));
compressor_3_2 u1_4646(.a(t_12510), .b(t_12509), .cin(t_11605), .o(t_13105), .cout(t_13106));
compressor_3_2 u1_4647(.a(t_12512), .b(t_12511), .cin(t_11610), .o(t_13107), .cout(t_13108));
compressor_3_2 u1_4648(.a(t_12514), .b(t_12513), .cin(t_11615), .o(t_13109), .cout(t_13110));
compressor_3_2 u1_4649(.a(t_12516), .b(t_12515), .cin(t_11620), .o(t_13111), .cout(t_13112));
compressor_3_2 u1_4650(.a(t_12518), .b(t_12517), .cin(t_11625), .o(t_13113), .cout(t_13114));
compressor_3_2 u1_4651(.a(t_12520), .b(t_12519), .cin(t_11630), .o(t_13115), .cout(t_13116));
compressor_3_2 u1_4652(.a(t_12522), .b(t_12521), .cin(t_11635), .o(t_13117), .cout(t_13118));
compressor_3_2 u1_4653(.a(t_12524), .b(t_12523), .cin(t_11640), .o(t_13119), .cout(t_13120));
compressor_3_2 u1_4654(.a(t_12526), .b(t_12525), .cin(t_11645), .o(t_13121), .cout(t_13122));
compressor_3_2 u1_4655(.a(t_12528), .b(t_12527), .cin(t_11650), .o(t_13123), .cout(t_13124));
compressor_3_2 u1_4656(.a(t_12530), .b(t_12529), .cin(t_11655), .o(t_13125), .cout(t_13126));
compressor_3_2 u1_4657(.a(t_12532), .b(t_12531), .cin(t_11660), .o(t_13127), .cout(t_13128));
compressor_3_2 u1_4658(.a(t_12534), .b(t_12533), .cin(t_11665), .o(t_13129), .cout(t_13130));
compressor_3_2 u1_4659(.a(t_12536), .b(t_12535), .cin(t_11670), .o(t_13131), .cout(t_13132));
half_adder u0_4660(.a(t_12538), .b(t_12537), .o(t_13133), .cout(t_13134));
half_adder u0_4661(.a(t_12541), .b(t_12539), .o(t_13135), .cout(t_13136));
compressor_3_2 u1_4662(.a(t_12544), .b(t_12542), .cin(t_11685), .o(t_13137), .cout(t_13138));
compressor_3_2 u1_4663(.a(t_12547), .b(t_12545), .cin(t_11690), .o(t_13139), .cout(t_13140));
compressor_3_2 u1_4664(.a(t_12550), .b(t_12548), .cin(t_11695), .o(t_13141), .cout(t_13142));
compressor_3_2 u1_4665(.a(t_12553), .b(t_12551), .cin(t_11700), .o(t_13143), .cout(t_13144));
compressor_3_2 u1_4666(.a(t_12556), .b(t_12554), .cin(t_11705), .o(t_13145), .cout(t_13146));
compressor_3_2 u1_4667(.a(t_12559), .b(t_12557), .cin(t_11710), .o(t_13147), .cout(t_13148));
compressor_3_2 u1_4668(.a(t_12562), .b(t_12560), .cin(t_11715), .o(t_13149), .cout(t_13150));
compressor_3_2 u1_4669(.a(t_12565), .b(t_12563), .cin(t_11720), .o(t_13151), .cout(t_13152));
compressor_3_2 u1_4670(.a(t_12568), .b(t_12566), .cin(t_11725), .o(t_13153), .cout(t_13154));
compressor_3_2 u1_4671(.a(t_12571), .b(t_12569), .cin(t_11730), .o(t_13155), .cout(t_13156));
compressor_3_2 u1_4672(.a(t_12574), .b(t_12572), .cin(t_11735), .o(t_13157), .cout(t_13158));
compressor_3_2 u1_4673(.a(t_12577), .b(t_12575), .cin(t_11740), .o(t_13159), .cout(t_13160));
compressor_3_2 u1_4674(.a(t_12580), .b(t_12578), .cin(t_11745), .o(t_13161), .cout(t_13162));
half_adder u0_4675(.a(t_12583), .b(t_12581), .o(t_13163), .cout(t_13164));
half_adder u0_4676(.a(t_12586), .b(t_12584), .o(t_13165), .cout(t_13166));
compressor_3_2 u1_4677(.a(t_12589), .b(t_12587), .cin(t_11762), .o(t_13167), .cout(t_13168));
compressor_3_2 u1_4678(.a(t_12592), .b(t_12590), .cin(t_11768), .o(t_13169), .cout(t_13170));
compressor_3_2 u1_4679(.a(t_12595), .b(t_12593), .cin(t_11774), .o(t_13171), .cout(t_13172));
compressor_3_2 u1_4680(.a(t_12598), .b(t_12596), .cin(t_11780), .o(t_13173), .cout(t_13174));
compressor_3_2 u1_4681(.a(t_12601), .b(t_12599), .cin(t_11786), .o(t_13175), .cout(t_13176));
half_adder u0_4682(.a(t_12604), .b(t_12602), .o(t_13177), .cout(t_13178));
half_adder u0_4683(.a(t_12607), .b(t_12605), .o(t_13179), .cout(t_13180));
compressor_3_2 u1_4684(.a(t_12610), .b(t_12608), .cin(t_11804), .o(t_13181), .cout(t_13182));
half_adder u0_4685(.a(t_12613), .b(t_12611), .o(t_13183), .cout(t_13184));
half_adder u0_4686(.a(t_12616), .b(t_12614), .o(t_13185), .cout(t_13186));
half_adder u0_4687(.a(t_12619), .b(t_12617), .o(t_13187), .cout(t_13188));
half_adder u0_4688(.a(t_12622), .b(t_12620), .o(t_13189), .cout(t_13190));
compressor_3_2 u1_4689(.a(t_12625), .b(t_12623), .cin(t_11834), .o(t_13191), .cout(t_13192));
compressor_3_2 u1_4690(.a(t_12628), .b(t_12626), .cin(t_11840), .o(t_13193), .cout(t_13194));
half_adder u0_4691(.a(t_12631), .b(t_12629), .o(t_13195), .cout(t_13196));
half_adder u0_4692(.a(t_12634), .b(t_12632), .o(t_13197), .cout(t_13198));
compressor_3_2 u1_4693(.a(t_12637), .b(t_12635), .cin(t_11858), .o(t_13199), .cout(t_13200));
half_adder u0_4694(.a(t_12640), .b(t_12638), .o(t_13201), .cout(t_13202));
half_adder u0_4695(.a(t_12643), .b(t_12641), .o(t_13203), .cout(t_13204));
half_adder u0_4696(.a(t_12646), .b(t_12644), .o(t_13205), .cout(t_13206));
half_adder u0_4697(.a(t_12649), .b(t_12647), .o(t_13207), .cout(t_13208));
compressor_3_2 u1_4698(.a(t_12652), .b(t_12650), .cin(t_11888), .o(t_13209), .cout(t_13210));
half_adder u0_4699(.a(t_12655), .b(t_12653), .o(t_13211), .cout(t_13212));
half_adder u0_4700(.a(t_12658), .b(t_12656), .o(t_13213), .cout(t_13214));
half_adder u0_4701(.a(t_12661), .b(t_12659), .o(t_13215), .cout(t_13216));
half_adder u0_4702(.a(t_12664), .b(t_12662), .o(t_13217), .cout(t_13218));
half_adder u0_4703(.a(t_12667), .b(t_12665), .o(t_13219), .cout(t_13220));
half_adder u0_4704(.a(t_12670), .b(t_12668), .o(t_13221), .cout(t_13222));
half_adder u0_4705(.a(t_12673), .b(t_12671), .o(t_13223), .cout(t_13224));
half_adder u0_4706(.a(t_12676), .b(t_12674), .o(t_13225), .cout(t_13226));
half_adder u0_4707(.a(t_12679), .b(t_12677), .o(t_13227), .cout(t_13228));
half_adder u0_4708(.a(t_12682), .b(t_12680), .o(t_13229), .cout(t_13230));
half_adder u0_4709(.a(t_12685), .b(t_12683), .o(t_13231), .cout(t_13232));
half_adder u0_4710(.a(t_12688), .b(t_12686), .o(t_13233), .cout(t_13234));
half_adder u0_4711(.a(t_12691), .b(t_12689), .o(t_13235), .cout(t_13236));
half_adder u0_4712(.a(t_12694), .b(t_12692), .o(t_13237), .cout(t_13238));
half_adder u0_4713(.a(t_12697), .b(t_12695), .o(t_13239), .cout(t_13240));
half_adder u0_4714(.a(t_12700), .b(t_12698), .o(t_13241), .cout(t_13242));
half_adder u0_4715(.a(t_12703), .b(t_12701), .o(t_13243), .cout(t_13244));
half_adder u0_4716(.a(t_12706), .b(t_12704), .o(t_13245), .cout(t_13246));
half_adder u0_4717(.a(t_12709), .b(t_12707), .o(t_13247), .cout(t_13248));
half_adder u0_4718(.a(t_12712), .b(t_12710), .o(t_13249), .cout(t_13250));
half_adder u0_4719(.a(t_12715), .b(t_12713), .o(t_13251), .cout(t_13252));
half_adder u0_4720(.a(t_12718), .b(t_12716), .o(t_13253), .cout(t_13254));
half_adder u0_4721(.a(t_12721), .b(t_12719), .o(t_13255), .cout(t_13256));
half_adder u0_4722(.a(t_12724), .b(t_12722), .o(t_13257), .cout(t_13258));
compressor_3_2 u1_4723(.a(t_12727), .b(t_12725), .cin(t_12038), .o(t_13259), .cout(t_13260));
half_adder u0_4724(.a(t_12730), .b(t_12728), .o(t_13261), .cout(t_13262));
half_adder u0_4725(.a(t_12733), .b(t_12731), .o(t_13263), .cout(t_13264));
half_adder u0_4726(.a(t_12736), .b(t_12734), .o(t_13265), .cout(t_13266));
half_adder u0_4727(.a(t_12739), .b(t_12737), .o(t_13267), .cout(t_13268));
half_adder u0_4728(.a(t_12742), .b(t_12740), .o(t_13269), .cout(t_13270));
half_adder u0_4729(.a(t_12745), .b(t_12743), .o(t_13271), .cout(t_13272));
half_adder u0_4730(.a(t_12748), .b(t_12746), .o(t_13273), .cout(t_13274));
half_adder u0_4731(.a(t_12751), .b(t_12749), .o(t_13275), .cout(t_13276));
half_adder u0_4732(.a(t_12754), .b(t_12752), .o(t_13277), .cout(t_13278));
half_adder u0_4733(.a(t_12757), .b(t_12755), .o(t_13279), .cout(t_13280));
half_adder u0_4734(.a(t_12760), .b(t_12758), .o(t_13281), .cout(t_13282));
half_adder u0_4735(.a(t_12763), .b(t_12761), .o(t_13283), .cout(t_13284));
half_adder u0_4736(.a(t_12766), .b(t_12764), .o(t_13285), .cout(t_13286));
half_adder u0_4737(.a(t_12769), .b(t_12767), .o(t_13287), .cout(t_13288));
half_adder u0_4738(.a(t_12772), .b(t_12770), .o(t_13289), .cout(t_13290));
half_adder u0_4739(.a(t_12775), .b(t_12773), .o(t_13291), .cout(t_13292));
half_adder u0_4740(.a(t_12778), .b(t_12776), .o(t_13293), .cout(t_13294));
half_adder u0_4741(.a(t_12781), .b(t_12779), .o(t_13295), .cout(t_13296));
half_adder u0_4742(.a(t_12784), .b(t_12782), .o(t_13297), .cout(t_13298));
half_adder u0_4743(.a(t_12787), .b(t_12785), .o(t_13299), .cout(t_13300));
half_adder u0_4744(.a(t_12790), .b(t_12788), .o(t_13301), .cout(t_13302));
half_adder u0_4745(.a(t_12793), .b(t_12791), .o(t_13303), .cout(t_13304));
half_adder u0_4746(.a(t_12796), .b(t_12794), .o(t_13305), .cout(t_13306));
half_adder u0_4747(.a(t_12799), .b(t_12797), .o(t_13307), .cout(t_13308));
half_adder u0_4748(.a(t_12802), .b(t_12800), .o(t_13309), .cout(t_13310));
half_adder u0_4749(.a(t_12805), .b(t_12803), .o(t_13311), .cout(t_13312));
half_adder u0_4750(.a(t_12808), .b(t_12806), .o(t_13313), .cout(t_13314));
half_adder u0_4751(.a(t_12811), .b(t_12809), .o(t_13315), .cout(t_13316));
half_adder u0_4752(.a(t_12814), .b(t_12812), .o(t_13317), .cout(t_13318));
half_adder u0_4753(.a(t_12817), .b(t_12815), .o(t_13319), .cout(t_13320));
half_adder u0_4754(.a(t_12820), .b(t_12818), .o(t_13321), .cout(t_13322));
half_adder u0_4755(.a(t_12823), .b(t_12821), .o(t_13323), .cout(t_13324));
half_adder u0_4756(.a(t_12826), .b(t_12824), .o(t_13325), .cout(t_13326));
half_adder u0_4757(.a(t_12828), .b(t_12827), .o(t_13327), .cout(t_13328));
half_adder u0_4758(.a(t_12830), .b(t_12829), .o(t_13329), .cout(t_13330));
half_adder u0_4759(.a(t_12832), .b(t_12831), .o(t_13331), .cout(t_13332));
half_adder u0_4760(.a(t_12834), .b(t_12833), .o(t_13333), .cout(t_13334));
half_adder u0_4761(.a(t_12836), .b(t_12835), .o(t_13335), .cout(t_13336));
half_adder u0_4762(.a(t_12838), .b(t_12837), .o(t_13337), .cout(t_13338));
half_adder u0_4763(.a(t_12840), .b(t_12839), .o(t_13339), .cout(t_13340));
half_adder u0_4764(.a(t_12842), .b(t_12841), .o(t_13341), .cout(t_13342));
half_adder u0_4765(.a(t_12844), .b(t_12843), .o(t_13343), .cout(t_13344));
half_adder u0_4766(.a(t_12846), .b(t_12845), .o(t_13345), .cout(t_13346));
half_adder u0_4767(.a(t_12848), .b(t_12847), .o(t_13347), .cout(t_13348));
half_adder u0_4768(.a(t_12850), .b(t_12849), .o(t_13349), .cout(t_13350));
half_adder u0_4769(.a(t_12852), .b(t_12851), .o(t_13351), .cout(t_13352));
half_adder u0_4770(.a(t_12854), .b(t_12853), .o(t_13353), .cout(t_13354));
half_adder u0_4771(.a(t_12856), .b(t_12855), .o(t_13355), .cout(t_13356));
half_adder u0_4772(.a(t_12858), .b(t_12857), .o(t_13357), .cout(t_13358));
half_adder u0_4773(.a(t_12860), .b(t_12859), .o(t_13359), .cout(t_13360));
half_adder u0_4774(.a(t_12862), .b(t_12861), .o(t_13361), .cout(t_13362));
half_adder u0_4775(.a(t_12864), .b(t_12863), .o(t_13363), .cout(t_13364));
half_adder u0_4776(.a(t_12866), .b(t_12865), .o(t_13365), .cout(t_13366));
half_adder u0_4777(.a(t_12868), .b(t_12867), .o(t_13367), .cout(t_13368));
half_adder u0_4778(.a(t_12870), .b(t_12869), .o(t_13369), .cout(t_13370));
half_adder u0_4779(.a(t_12872), .b(t_12871), .o(t_13371), .cout(t_13372));
half_adder u0_4780(.a(t_12874), .b(t_12873), .o(t_13373), .cout(t_13374));
half_adder u0_4781(.a(t_12876), .b(t_12875), .o(t_13375), .cout(t_13376));
half_adder u0_4782(.a(t_12878), .b(t_12877), .o(t_13377), .cout(t_13378));
half_adder u0_4783(.a(t_12880), .b(t_12879), .o(t_13379), .cout(t_13380));
half_adder u0_4784(.a(t_12882), .b(t_12881), .o(t_13381), .cout(t_13382));
half_adder u0_4785(.a(t_12884), .b(t_12883), .o(t_13383), .cout(t_13384));
half_adder u0_4786(.a(t_12886), .b(t_12885), .o(t_13385), .cout(t_13386));
half_adder u0_4787(.a(t_12888), .b(t_12887), .o(t_13387), .cout(t_13388));
half_adder u0_4788(.a(t_12890), .b(t_12889), .o(t_13389), .cout(t_13390));
half_adder u0_4789(.a(t_12892), .b(t_12891), .o(t_13391), .cout(t_13392));
half_adder u0_4790(.a(t_12894), .b(t_12893), .o(t_13393), .cout(t_13394));
half_adder u0_4791(.a(t_12896), .b(t_12895), .o(t_13395), .cout(t_13396));
half_adder u0_4792(.a(t_12898), .b(t_12897), .o(t_13397), .cout(t_13398));
half_adder u0_4793(.a(t_12900), .b(t_12899), .o(t_13399), .cout(t_13400));
half_adder u0_4794(.a(t_12902), .b(t_12901), .o(t_13401), .cout(t_13402));
half_adder u0_4795(.a(t_12904), .b(t_12903), .o(t_13403), .cout(t_13404));
half_adder u0_4796(.a(t_12906), .b(t_12905), .o(t_13405), .cout(t_13406));
half_adder u0_4797(.a(t_12908), .b(t_12907), .o(t_13407), .cout(t_13408));
half_adder u0_4798(.a(t_12910), .b(t_12909), .o(t_13409), .cout(t_13410));
half_adder u0_4799(.a(t_12912), .b(t_12911), .o(t_13411), .cout(t_13412));
half_adder u0_4800(.a(t_12914), .b(t_12913), .o(t_13413), .cout(t_13414));
half_adder u0_4801(.a(t_12916), .b(t_12915), .o(t_13415), .cout(t_13416));
half_adder u0_4802(.a(t_12918), .b(t_12917), .o(t_13417), .cout(t_13418));
half_adder u0_4803(.a(t_12920), .b(t_12919), .o(t_13419), .cout(t_13420));
half_adder u0_4804(.a(t_12922), .b(t_12921), .o(t_13421), .cout(t_13422));
half_adder u0_4805(.a(t_12924), .b(t_12923), .o(t_13423), .cout(t_13424));
half_adder u0_4806(.a(t_12926), .b(t_12925), .o(t_13425), .cout(t_13426));
half_adder u0_4807(.a(t_12928), .b(t_12927), .o(t_13427), .cout(t_13428));
half_adder u0_4808(.a(t_12930), .b(t_12929), .o(t_13429), .cout(t_13430));
half_adder u0_4809(.a(t_12932), .b(t_12931), .o(t_13431), .cout(t_13432));
half_adder u0_4810(.a(t_12934), .b(t_12933), .o(t_13433), .cout(t_13434));
half_adder u0_4811(.a(t_12936), .b(t_12935), .o(t_13435), .cout(t_13436));
half_adder u0_4812(.a(t_12938), .b(t_12937), .o(t_13437), .cout(t_13438));
half_adder u0_4813(.a(t_12940), .b(t_12939), .o(t_13439), .cout(t_13440));
half_adder u0_4814(.a(t_12942), .b(t_12941), .o(t_13441), .cout(t_13442));
half_adder u0_4815(.a(t_12944), .b(t_12943), .o(t_13443), .cout(t_13444));
half_adder u0_4816(.a(t_12946), .b(t_12945), .o(t_13445), .cout());

/* Output nets Compression result */
assign compress_a = {
 t_13444, t_13442, t_13440, t_13438,
 t_13436, t_13434, t_13432, t_13430,
 t_13428, t_13426, t_13424, t_13422,
 t_13420, t_13418, t_13416, t_13414,
 t_13412, t_13410, t_13408, t_13406,
 t_13404, t_13402, t_13400, t_13398,
 t_13396, t_13394, t_13392, t_13390,
 t_13388, t_13386, t_13384, t_13382,
 t_13380, t_13378, t_13376, t_13374,
 t_13372, t_13370, t_13368, t_13366,
 t_13364, t_13362, t_13360, t_13358,
 t_13356, t_13354, t_13352, t_13350,
 t_13348, t_13346, t_13344, t_13342,
 t_13340, t_13338, t_13336, t_13334,
 t_13332, t_13330, t_13328, t_13326,
 t_13324, t_13322, t_13320, t_13318,
 t_13316, t_13314, t_13312, t_13310,
 t_13308, t_13306, t_13304, t_13302,
 t_13300, t_13298, t_13296, t_13294,
 t_13292, t_13290, t_13288, t_13286,
 t_13284, t_13282, t_13280, t_13278,
 t_13276, t_13274, t_13272, t_13270,
 t_13268, t_13266, t_13264, t_13262,
 t_13260, t_13258, t_13256, t_13254,
 t_13252, t_13250, t_13248, t_13246,
 t_13244, t_13242, t_13240, t_13238,
 t_13236, t_13234, t_13232, t_13230,
 t_13228, t_13226, t_13224, t_13222,
 t_13220, t_13218, t_13216, t_13214,
 t_13212, t_13210, t_13208, t_13206,
 t_13204, t_13202, t_13200, t_13198,
 t_13196, t_13194, t_13192, t_13190,
 t_13188, t_13186, t_13184, t_13182,
 t_13180, t_13178, t_13176, t_13174,
 t_13172, t_13170, t_13168, t_13166,
 t_13164, t_13162, t_13160, t_13158,
 t_13156, t_13154, t_13152, t_13150,
 t_13148, t_13146, t_13144, t_13142,
 t_13140, t_13138, t_13136, t_13134,
 t_13132, t_13130, t_13128, t_13126,
 t_13124, t_13122, t_13120, t_13118,
 t_13116, t_13114, t_13112, t_13110,
 t_13108, t_13106, t_13104, t_13102,
 t_13100, t_13098, t_13096, t_13094,
 t_13092, t_13090, t_13088, t_13086,
 t_13084, t_13082, t_13080, t_13078,
 t_13076, t_13074, t_13072, t_13070,
 t_13068, t_13066, t_13064, t_13062,
 t_13060, t_13058, t_13056, t_13054,
 t_13052, t_13050, t_13048, t_13046,
 t_13044, t_13042, t_13040, t_13038,
 t_13036, t_13034, t_13032, t_13030,
 t_13028, t_13026, t_13024, t_13022,
 t_13020, t_13018, t_13016, t_13014,
 t_13012, t_13010, t_13008, t_13006,
 t_13004, t_13002, t_13000, t_12998,
 t_12996, t_12994, t_12992, t_12990,
 t_12988, t_12986, t_12984, t_12982,
 t_12980, t_12978, t_12976, t_12974,
 t_12972, t_12970, t_12968, t_12966,
 t_12964, t_12962, t_12960, t_12958,
 t_12956, t_12954, t_12952, t_12950,
 t_12949, t_12352, t_12947, t_12350,
 t_11371,  t_9620,  t_6335,     t_0
};
assign compress_b = {
 t_13445, t_13443, t_13441, t_13439,
 t_13437, t_13435, t_13433, t_13431,
 t_13429, t_13427, t_13425, t_13423,
 t_13421, t_13419, t_13417, t_13415,
 t_13413, t_13411, t_13409, t_13407,
 t_13405, t_13403, t_13401, t_13399,
 t_13397, t_13395, t_13393, t_13391,
 t_13389, t_13387, t_13385, t_13383,
 t_13381, t_13379, t_13377, t_13375,
 t_13373, t_13371, t_13369, t_13367,
 t_13365, t_13363, t_13361, t_13359,
 t_13357, t_13355, t_13353, t_13351,
 t_13349, t_13347, t_13345, t_13343,
 t_13341, t_13339, t_13337, t_13335,
 t_13333, t_13331, t_13329, t_13327,
 t_13325, t_13323, t_13321, t_13319,
 t_13317, t_13315, t_13313, t_13311,
 t_13309, t_13307, t_13305, t_13303,
 t_13301, t_13299, t_13297, t_13295,
 t_13293, t_13291, t_13289, t_13287,
 t_13285, t_13283, t_13281, t_13279,
 t_13277, t_13275, t_13273, t_13271,
 t_13269, t_13267, t_13265, t_13263,
 t_13261, t_13259, t_13257, t_13255,
 t_13253, t_13251, t_13249, t_13247,
 t_13245, t_13243, t_13241, t_13239,
 t_13237, t_13235, t_13233, t_13231,
 t_13229, t_13227, t_13225, t_13223,
 t_13221, t_13219, t_13217, t_13215,
 t_13213, t_13211, t_13209, t_13207,
 t_13205, t_13203, t_13201, t_13199,
 t_13197, t_13195, t_13193, t_13191,
 t_13189, t_13187, t_13185, t_13183,
 t_13181, t_13179, t_13177, t_13175,
 t_13173, t_13171, t_13169, t_13167,
 t_13165, t_13163, t_13161, t_13159,
 t_13157, t_13155, t_13153, t_13151,
 t_13149, t_13147, t_13145, t_13143,
 t_13141, t_13139, t_13137, t_13135,
 t_13133, t_13131, t_13129, t_13127,
 t_13125, t_13123, t_13121, t_13119,
 t_13117, t_13115, t_13113, t_13111,
 t_13109, t_13107, t_13105, t_13103,
 t_13101, t_13099, t_13097, t_13095,
 t_13093, t_13091, t_13089, t_13087,
 t_13085, t_13083, t_13081, t_13079,
 t_13077, t_13075, t_13073, t_13071,
 t_13069, t_13067, t_13065, t_13063,
 t_13061, t_13059, t_13057, t_13055,
 t_13053, t_13051, t_13049, t_13047,
 t_13045, t_13043, t_13041, t_13039,
 t_13037, t_13035, t_13033, t_13031,
 t_13029, t_13027, t_13025, t_13023,
 t_13021, t_13019, t_13017, t_13015,
 t_13013, t_13011, t_13009, t_13007,
 t_13005, t_13003, t_13001, t_12999,
 t_12997, t_12995, t_12993, t_12991,
 t_12989, t_12987, t_12985, t_12983,
 t_12981, t_12979, t_12977, t_12975,
 t_12973, t_12971, t_12969, t_12967,
 t_12965, t_12963, t_12961, t_12959,
 t_12957, t_12955, t_12953, t_12951,
    1'b0, t_12948,    1'b0,    1'b0,
    1'b0,    1'b0,    1'b0,    1'b0
};

endmodule

/********************************************************************************/

module booth_coder(
//inputs
	sign,
	a,
	b,
//outputs
	partial_products,
	carry
);

parameter width = 8;

input wire sign;
input wire [width-1:0] a;
input wire [width-1:0] b;
output wire [(width+2)*(width/2+1)-1:0] partial_products;
output reg [width/2-1:0] carry;

reg [(width+2)*(width/2)-1:0] codingdata;
wire [width:0] b_ = {sign&b[width-1], b};
wire [width:0] a_temp = {a, 1'b0};

generate
	genvar i;
	for (i=0; i<width; i=i+2)
	begin: encoder
		always @ (*)
		begin
			case (a_temp[i+2:i])
			3'b0, 3'd7: begin
				codingdata[`INDEX] = {1'b1, {(width+1){1'b0}}};
				carry[i/2] = 1'b0;
			end
			3'd1, 3'd2: begin
				codingdata[`INDEX] = {~b_[width], b_};
				carry[i/2] = 1'b0;
			end
			3'd3: begin
				codingdata[`INDEX] = {~b_[width], b, 1'b0};
				carry[i/2] = 1'b0;
			end
			3'd4: begin
				codingdata[`INDEX] = {b_[width], ~b, 1'b1};
				carry[i/2] = 1'b1;
			end
			3'd5, 3'd6: begin
				codingdata[`INDEX] = {b_[width], ~b_};
				carry[i/2] = 1'b1;
			end
			default: begin
				codingdata[`INDEX] = {(width+2){1'b0}};
				carry[i/2] = 1'b0;
			end
			endcase
		end
	end
endgenerate

function [255:0] sign_sum(input integer n);
integer i;
begin
	for (sign_sum=0, i=0; i<n; i=i+2)
		sign_sum = sign_sum + ({256{1'b1}} << (n-i-2));
	sign_sum = sign_sum << 3;
end
endfunction

wire [width+1:0] signsum = sign_sum(width);
wire [width-1:0] unsign_correct = {width{ a[width-1]&(~sign) }} & b;
wire [width+1:0] extra_product = {signsum[width+1:2]+unsign_correct, signsum[1:0]};

assign partial_products = {extra_product, codingdata};

endmodule

/********************************************************************************/

module multer(
//inputs
    sign,
    A,
    B,
//outputs
    P
);

parameter width = 8;

input wire sign;
input wire [width-1:0] A;
input wire [width-1:0] B;
output wire [2*width-1:0] P;

wire [(width+2)*(width/2+1)-1:0] partial_products;
wire [width/2-1:0] carry;
wire [2*width-1:0] compress_a;
wire [2*width-1:0] compress_b;

booth_coder encoder(.sign(sign), .a(A), .b(B), .partial_products(partial_products), .carry(carry));
defparam
    encoder.width=width;

generate
	case (width)
		32 : _32_wallace_tree compressor(.partial_products(partial_products), .carry(carry), .compress_a(compress_a), .compress_b(compress_b));
		64 : _64_wallace_tree compressor(.partial_products(partial_products), .carry(carry), .compress_a(compress_a), .compress_b(compress_b));
		128: _128_wallace_tree compressor(.partial_products(partial_products), .carry(carry), .compress_a(compress_a), .compress_b(compress_b));
		default: _32_wallace_tree compressor(.partial_products(partial_products), .carry(carry), .compress_a(compress_a), .compress_b(compress_b));
	endcase
endgenerate

assign P = compress_a + compress_b;

endmodule

`undef INDEX
